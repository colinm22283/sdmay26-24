magic
tech sky130A
magscale 1 2
timestamp 1763051408
<< obsli1 >>
rect 1104 2159 58880 57681
<< obsm1 >>
rect 934 2128 59786 57712
<< metal2 >>
rect 14922 0 14978 800
rect 44914 0 44970 800
<< obsm2 >>
rect 938 856 59780 57701
rect 938 800 14866 856
rect 15034 800 44858 856
rect 45026 800 59780 856
<< metal3 >>
rect 59200 55496 60000 55616
rect 0 55224 800 55344
rect 59200 54680 60000 54800
rect 59200 53864 60000 53984
rect 0 53592 800 53712
rect 59200 53048 60000 53168
rect 59200 52232 60000 52352
rect 0 51960 800 52080
rect 59200 51416 60000 51536
rect 59200 50600 60000 50720
rect 0 50328 800 50448
rect 59200 49784 60000 49904
rect 59200 48968 60000 49088
rect 0 48696 800 48816
rect 59200 48152 60000 48272
rect 59200 47336 60000 47456
rect 0 47064 800 47184
rect 59200 46520 60000 46640
rect 59200 45704 60000 45824
rect 0 45432 800 45552
rect 59200 44888 60000 45008
rect 59200 44072 60000 44192
rect 0 43800 800 43920
rect 59200 43256 60000 43376
rect 59200 42440 60000 42560
rect 0 42168 800 42288
rect 59200 41624 60000 41744
rect 59200 40808 60000 40928
rect 0 40536 800 40656
rect 59200 39992 60000 40112
rect 59200 39176 60000 39296
rect 0 38904 800 39024
rect 59200 38360 60000 38480
rect 59200 37544 60000 37664
rect 0 37272 800 37392
rect 59200 36728 60000 36848
rect 59200 35912 60000 36032
rect 0 35640 800 35760
rect 59200 35096 60000 35216
rect 59200 34280 60000 34400
rect 0 34008 800 34128
rect 59200 33464 60000 33584
rect 59200 32648 60000 32768
rect 0 32376 800 32496
rect 59200 31832 60000 31952
rect 59200 31016 60000 31136
rect 0 30744 800 30864
rect 59200 30200 60000 30320
rect 59200 29384 60000 29504
rect 0 29112 800 29232
rect 59200 28568 60000 28688
rect 59200 27752 60000 27872
rect 0 27480 800 27600
rect 59200 26936 60000 27056
rect 59200 26120 60000 26240
rect 0 25848 800 25968
rect 59200 25304 60000 25424
rect 59200 24488 60000 24608
rect 0 24216 800 24336
rect 59200 23672 60000 23792
rect 59200 22856 60000 22976
rect 0 22584 800 22704
rect 59200 22040 60000 22160
rect 59200 21224 60000 21344
rect 0 20952 800 21072
rect 59200 20408 60000 20528
rect 59200 19592 60000 19712
rect 0 19320 800 19440
rect 59200 18776 60000 18896
rect 59200 17960 60000 18080
rect 0 17688 800 17808
rect 59200 17144 60000 17264
rect 59200 16328 60000 16448
rect 0 16056 800 16176
rect 59200 15512 60000 15632
rect 59200 14696 60000 14816
rect 0 14424 800 14544
rect 59200 13880 60000 14000
rect 59200 13064 60000 13184
rect 0 12792 800 12912
rect 59200 12248 60000 12368
rect 59200 11432 60000 11552
rect 0 11160 800 11280
rect 59200 10616 60000 10736
rect 59200 9800 60000 9920
rect 0 9528 800 9648
rect 59200 8984 60000 9104
rect 59200 8168 60000 8288
rect 0 7896 800 8016
rect 59200 7352 60000 7472
rect 59200 6536 60000 6656
rect 0 6264 800 6384
rect 59200 5720 60000 5840
rect 59200 4904 60000 5024
rect 0 4632 800 4752
rect 59200 4088 60000 4208
<< obsm3 >>
rect 798 55696 59200 57697
rect 798 55424 59120 55696
rect 880 55416 59120 55424
rect 880 55144 59200 55416
rect 798 54880 59200 55144
rect 798 54600 59120 54880
rect 798 54064 59200 54600
rect 798 53792 59120 54064
rect 880 53784 59120 53792
rect 880 53512 59200 53784
rect 798 53248 59200 53512
rect 798 52968 59120 53248
rect 798 52432 59200 52968
rect 798 52160 59120 52432
rect 880 52152 59120 52160
rect 880 51880 59200 52152
rect 798 51616 59200 51880
rect 798 51336 59120 51616
rect 798 50800 59200 51336
rect 798 50528 59120 50800
rect 880 50520 59120 50528
rect 880 50248 59200 50520
rect 798 49984 59200 50248
rect 798 49704 59120 49984
rect 798 49168 59200 49704
rect 798 48896 59120 49168
rect 880 48888 59120 48896
rect 880 48616 59200 48888
rect 798 48352 59200 48616
rect 798 48072 59120 48352
rect 798 47536 59200 48072
rect 798 47264 59120 47536
rect 880 47256 59120 47264
rect 880 46984 59200 47256
rect 798 46720 59200 46984
rect 798 46440 59120 46720
rect 798 45904 59200 46440
rect 798 45632 59120 45904
rect 880 45624 59120 45632
rect 880 45352 59200 45624
rect 798 45088 59200 45352
rect 798 44808 59120 45088
rect 798 44272 59200 44808
rect 798 44000 59120 44272
rect 880 43992 59120 44000
rect 880 43720 59200 43992
rect 798 43456 59200 43720
rect 798 43176 59120 43456
rect 798 42640 59200 43176
rect 798 42368 59120 42640
rect 880 42360 59120 42368
rect 880 42088 59200 42360
rect 798 41824 59200 42088
rect 798 41544 59120 41824
rect 798 41008 59200 41544
rect 798 40736 59120 41008
rect 880 40728 59120 40736
rect 880 40456 59200 40728
rect 798 40192 59200 40456
rect 798 39912 59120 40192
rect 798 39376 59200 39912
rect 798 39104 59120 39376
rect 880 39096 59120 39104
rect 880 38824 59200 39096
rect 798 38560 59200 38824
rect 798 38280 59120 38560
rect 798 37744 59200 38280
rect 798 37472 59120 37744
rect 880 37464 59120 37472
rect 880 37192 59200 37464
rect 798 36928 59200 37192
rect 798 36648 59120 36928
rect 798 36112 59200 36648
rect 798 35840 59120 36112
rect 880 35832 59120 35840
rect 880 35560 59200 35832
rect 798 35296 59200 35560
rect 798 35016 59120 35296
rect 798 34480 59200 35016
rect 798 34208 59120 34480
rect 880 34200 59120 34208
rect 880 33928 59200 34200
rect 798 33664 59200 33928
rect 798 33384 59120 33664
rect 798 32848 59200 33384
rect 798 32576 59120 32848
rect 880 32568 59120 32576
rect 880 32296 59200 32568
rect 798 32032 59200 32296
rect 798 31752 59120 32032
rect 798 31216 59200 31752
rect 798 30944 59120 31216
rect 880 30936 59120 30944
rect 880 30664 59200 30936
rect 798 30400 59200 30664
rect 798 30120 59120 30400
rect 798 29584 59200 30120
rect 798 29312 59120 29584
rect 880 29304 59120 29312
rect 880 29032 59200 29304
rect 798 28768 59200 29032
rect 798 28488 59120 28768
rect 798 27952 59200 28488
rect 798 27680 59120 27952
rect 880 27672 59120 27680
rect 880 27400 59200 27672
rect 798 27136 59200 27400
rect 798 26856 59120 27136
rect 798 26320 59200 26856
rect 798 26048 59120 26320
rect 880 26040 59120 26048
rect 880 25768 59200 26040
rect 798 25504 59200 25768
rect 798 25224 59120 25504
rect 798 24688 59200 25224
rect 798 24416 59120 24688
rect 880 24408 59120 24416
rect 880 24136 59200 24408
rect 798 23872 59200 24136
rect 798 23592 59120 23872
rect 798 23056 59200 23592
rect 798 22784 59120 23056
rect 880 22776 59120 22784
rect 880 22504 59200 22776
rect 798 22240 59200 22504
rect 798 21960 59120 22240
rect 798 21424 59200 21960
rect 798 21152 59120 21424
rect 880 21144 59120 21152
rect 880 20872 59200 21144
rect 798 20608 59200 20872
rect 798 20328 59120 20608
rect 798 19792 59200 20328
rect 798 19520 59120 19792
rect 880 19512 59120 19520
rect 880 19240 59200 19512
rect 798 18976 59200 19240
rect 798 18696 59120 18976
rect 798 18160 59200 18696
rect 798 17888 59120 18160
rect 880 17880 59120 17888
rect 880 17608 59200 17880
rect 798 17344 59200 17608
rect 798 17064 59120 17344
rect 798 16528 59200 17064
rect 798 16256 59120 16528
rect 880 16248 59120 16256
rect 880 15976 59200 16248
rect 798 15712 59200 15976
rect 798 15432 59120 15712
rect 798 14896 59200 15432
rect 798 14624 59120 14896
rect 880 14616 59120 14624
rect 880 14344 59200 14616
rect 798 14080 59200 14344
rect 798 13800 59120 14080
rect 798 13264 59200 13800
rect 798 12992 59120 13264
rect 880 12984 59120 12992
rect 880 12712 59200 12984
rect 798 12448 59200 12712
rect 798 12168 59120 12448
rect 798 11632 59200 12168
rect 798 11360 59120 11632
rect 880 11352 59120 11360
rect 880 11080 59200 11352
rect 798 10816 59200 11080
rect 798 10536 59120 10816
rect 798 10000 59200 10536
rect 798 9728 59120 10000
rect 880 9720 59120 9728
rect 880 9448 59200 9720
rect 798 9184 59200 9448
rect 798 8904 59120 9184
rect 798 8368 59200 8904
rect 798 8096 59120 8368
rect 880 8088 59120 8096
rect 880 7816 59200 8088
rect 798 7552 59200 7816
rect 798 7272 59120 7552
rect 798 6736 59200 7272
rect 798 6464 59120 6736
rect 880 6456 59120 6464
rect 880 6184 59200 6456
rect 798 5920 59200 6184
rect 798 5640 59120 5920
rect 798 5104 59200 5640
rect 798 4832 59120 5104
rect 880 4824 59120 4832
rect 880 4552 59200 4824
rect 798 4288 59200 4552
rect 798 4008 59120 4288
rect 798 2143 59200 4008
<< metal4 >>
rect 4208 2128 4528 57712
rect 19568 2128 19888 57712
rect 34928 2128 35248 57712
rect 50288 2128 50608 57712
<< obsm4 >>
rect 6131 6427 19488 48109
rect 19968 6427 34848 48109
rect 35328 6427 50208 48109
rect 50688 6427 57901 48109
<< labels >>
rlabel metal3 s 59200 4088 60000 4208 6 a_i[0]
port 1 nsew signal input
rlabel metal3 s 59200 12248 60000 12368 6 a_i[10]
port 2 nsew signal input
rlabel metal3 s 59200 13064 60000 13184 6 a_i[11]
port 3 nsew signal input
rlabel metal3 s 59200 13880 60000 14000 6 a_i[12]
port 4 nsew signal input
rlabel metal3 s 59200 14696 60000 14816 6 a_i[13]
port 5 nsew signal input
rlabel metal3 s 59200 15512 60000 15632 6 a_i[14]
port 6 nsew signal input
rlabel metal3 s 59200 16328 60000 16448 6 a_i[15]
port 7 nsew signal input
rlabel metal3 s 59200 17144 60000 17264 6 a_i[16]
port 8 nsew signal input
rlabel metal3 s 59200 17960 60000 18080 6 a_i[17]
port 9 nsew signal input
rlabel metal3 s 59200 18776 60000 18896 6 a_i[18]
port 10 nsew signal input
rlabel metal3 s 59200 19592 60000 19712 6 a_i[19]
port 11 nsew signal input
rlabel metal3 s 59200 4904 60000 5024 6 a_i[1]
port 12 nsew signal input
rlabel metal3 s 59200 20408 60000 20528 6 a_i[20]
port 13 nsew signal input
rlabel metal3 s 59200 21224 60000 21344 6 a_i[21]
port 14 nsew signal input
rlabel metal3 s 59200 22040 60000 22160 6 a_i[22]
port 15 nsew signal input
rlabel metal3 s 59200 22856 60000 22976 6 a_i[23]
port 16 nsew signal input
rlabel metal3 s 59200 23672 60000 23792 6 a_i[24]
port 17 nsew signal input
rlabel metal3 s 59200 24488 60000 24608 6 a_i[25]
port 18 nsew signal input
rlabel metal3 s 59200 25304 60000 25424 6 a_i[26]
port 19 nsew signal input
rlabel metal3 s 59200 26120 60000 26240 6 a_i[27]
port 20 nsew signal input
rlabel metal3 s 59200 26936 60000 27056 6 a_i[28]
port 21 nsew signal input
rlabel metal3 s 59200 27752 60000 27872 6 a_i[29]
port 22 nsew signal input
rlabel metal3 s 59200 5720 60000 5840 6 a_i[2]
port 23 nsew signal input
rlabel metal3 s 59200 28568 60000 28688 6 a_i[30]
port 24 nsew signal input
rlabel metal3 s 59200 29384 60000 29504 6 a_i[31]
port 25 nsew signal input
rlabel metal3 s 59200 6536 60000 6656 6 a_i[3]
port 26 nsew signal input
rlabel metal3 s 59200 7352 60000 7472 6 a_i[4]
port 27 nsew signal input
rlabel metal3 s 59200 8168 60000 8288 6 a_i[5]
port 28 nsew signal input
rlabel metal3 s 59200 8984 60000 9104 6 a_i[6]
port 29 nsew signal input
rlabel metal3 s 59200 9800 60000 9920 6 a_i[7]
port 30 nsew signal input
rlabel metal3 s 59200 10616 60000 10736 6 a_i[8]
port 31 nsew signal input
rlabel metal3 s 59200 11432 60000 11552 6 a_i[9]
port 32 nsew signal input
rlabel metal3 s 59200 30200 60000 30320 6 b_i[0]
port 33 nsew signal input
rlabel metal3 s 59200 38360 60000 38480 6 b_i[10]
port 34 nsew signal input
rlabel metal3 s 59200 39176 60000 39296 6 b_i[11]
port 35 nsew signal input
rlabel metal3 s 59200 39992 60000 40112 6 b_i[12]
port 36 nsew signal input
rlabel metal3 s 59200 40808 60000 40928 6 b_i[13]
port 37 nsew signal input
rlabel metal3 s 59200 41624 60000 41744 6 b_i[14]
port 38 nsew signal input
rlabel metal3 s 59200 42440 60000 42560 6 b_i[15]
port 39 nsew signal input
rlabel metal3 s 59200 43256 60000 43376 6 b_i[16]
port 40 nsew signal input
rlabel metal3 s 59200 44072 60000 44192 6 b_i[17]
port 41 nsew signal input
rlabel metal3 s 59200 44888 60000 45008 6 b_i[18]
port 42 nsew signal input
rlabel metal3 s 59200 45704 60000 45824 6 b_i[19]
port 43 nsew signal input
rlabel metal3 s 59200 31016 60000 31136 6 b_i[1]
port 44 nsew signal input
rlabel metal3 s 59200 46520 60000 46640 6 b_i[20]
port 45 nsew signal input
rlabel metal3 s 59200 47336 60000 47456 6 b_i[21]
port 46 nsew signal input
rlabel metal3 s 59200 48152 60000 48272 6 b_i[22]
port 47 nsew signal input
rlabel metal3 s 59200 48968 60000 49088 6 b_i[23]
port 48 nsew signal input
rlabel metal3 s 59200 49784 60000 49904 6 b_i[24]
port 49 nsew signal input
rlabel metal3 s 59200 50600 60000 50720 6 b_i[25]
port 50 nsew signal input
rlabel metal3 s 59200 51416 60000 51536 6 b_i[26]
port 51 nsew signal input
rlabel metal3 s 59200 52232 60000 52352 6 b_i[27]
port 52 nsew signal input
rlabel metal3 s 59200 53048 60000 53168 6 b_i[28]
port 53 nsew signal input
rlabel metal3 s 59200 53864 60000 53984 6 b_i[29]
port 54 nsew signal input
rlabel metal3 s 59200 31832 60000 31952 6 b_i[2]
port 55 nsew signal input
rlabel metal3 s 59200 54680 60000 54800 6 b_i[30]
port 56 nsew signal input
rlabel metal3 s 59200 55496 60000 55616 6 b_i[31]
port 57 nsew signal input
rlabel metal3 s 59200 32648 60000 32768 6 b_i[3]
port 58 nsew signal input
rlabel metal3 s 59200 33464 60000 33584 6 b_i[4]
port 59 nsew signal input
rlabel metal3 s 59200 34280 60000 34400 6 b_i[5]
port 60 nsew signal input
rlabel metal3 s 59200 35096 60000 35216 6 b_i[6]
port 61 nsew signal input
rlabel metal3 s 59200 35912 60000 36032 6 b_i[7]
port 62 nsew signal input
rlabel metal3 s 59200 36728 60000 36848 6 b_i[8]
port 63 nsew signal input
rlabel metal3 s 59200 37544 60000 37664 6 b_i[9]
port 64 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 clk
port 65 nsew signal input
rlabel metal2 s 44914 0 44970 800 6 nrst
port 66 nsew signal input
rlabel metal4 s 4208 2128 4528 57712 6 vccd1
port 67 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 57712 6 vccd1
port 67 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 57712 6 vssd1
port 68 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 57712 6 vssd1
port 68 nsew ground bidirectional
rlabel metal3 s 0 4632 800 4752 6 y_o[0]
port 69 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 y_o[10]
port 70 nsew signal output
rlabel metal3 s 0 22584 800 22704 6 y_o[11]
port 71 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 y_o[12]
port 72 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 y_o[13]
port 73 nsew signal output
rlabel metal3 s 0 27480 800 27600 6 y_o[14]
port 74 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 y_o[15]
port 75 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 y_o[16]
port 76 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 y_o[17]
port 77 nsew signal output
rlabel metal3 s 0 34008 800 34128 6 y_o[18]
port 78 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 y_o[19]
port 79 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 y_o[1]
port 80 nsew signal output
rlabel metal3 s 0 37272 800 37392 6 y_o[20]
port 81 nsew signal output
rlabel metal3 s 0 38904 800 39024 6 y_o[21]
port 82 nsew signal output
rlabel metal3 s 0 40536 800 40656 6 y_o[22]
port 83 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 y_o[23]
port 84 nsew signal output
rlabel metal3 s 0 43800 800 43920 6 y_o[24]
port 85 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 y_o[25]
port 86 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 y_o[26]
port 87 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 y_o[27]
port 88 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 y_o[28]
port 89 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 y_o[29]
port 90 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 y_o[2]
port 91 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 y_o[30]
port 92 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 y_o[31]
port 93 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 y_o[3]
port 94 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 y_o[4]
port 95 nsew signal output
rlabel metal3 s 0 12792 800 12912 6 y_o[5]
port 96 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 y_o[6]
port 97 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 y_o[7]
port 98 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 y_o[8]
port 99 nsew signal output
rlabel metal3 s 0 19320 800 19440 6 y_o[9]
port 100 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11355254
string GDS_FILE /home/sforde22/Caravel/sdmay26-24/openlane/mac_pipe/runs/25_11_13_10_25/results/signoff/mac_piped.magic.gds
string GDS_START 458822
<< end >>

