magic
tech sky130A
magscale 1 2
timestamp 1760900936
<< obsli1 >>
rect 1104 2159 118864 87601
<< obsm1 >>
rect 198 8 119126 87712
<< metal2 >>
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8206 0 8262 800
rect 8574 0 8630 800
rect 8942 0 8998 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10782 0 10838 800
rect 11150 0 11206 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13358 0 13414 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15934 0 15990 800
rect 16302 0 16358 800
rect 16670 0 16726 800
rect 17038 0 17094 800
rect 17406 0 17462 800
rect 17774 0 17830 800
rect 18142 0 18198 800
rect 18510 0 18566 800
rect 18878 0 18934 800
rect 19246 0 19302 800
rect 19614 0 19670 800
rect 19982 0 20038 800
rect 20350 0 20406 800
rect 20718 0 20774 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21822 0 21878 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22926 0 22982 800
rect 23294 0 23350 800
rect 23662 0 23718 800
rect 24030 0 24086 800
rect 24398 0 24454 800
rect 24766 0 24822 800
rect 25134 0 25190 800
rect 25502 0 25558 800
rect 25870 0 25926 800
rect 26238 0 26294 800
rect 26606 0 26662 800
rect 26974 0 27030 800
rect 27342 0 27398 800
rect 27710 0 27766 800
rect 28078 0 28134 800
rect 28446 0 28502 800
rect 28814 0 28870 800
rect 29182 0 29238 800
rect 29550 0 29606 800
rect 29918 0 29974 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31390 0 31446 800
rect 31758 0 31814 800
rect 32126 0 32182 800
rect 32494 0 32550 800
rect 32862 0 32918 800
rect 33230 0 33286 800
rect 33598 0 33654 800
rect 33966 0 34022 800
rect 34334 0 34390 800
rect 34702 0 34758 800
rect 35070 0 35126 800
rect 35438 0 35494 800
rect 35806 0 35862 800
rect 36174 0 36230 800
rect 36542 0 36598 800
rect 36910 0 36966 800
rect 37278 0 37334 800
rect 37646 0 37702 800
rect 38014 0 38070 800
rect 38382 0 38438 800
rect 38750 0 38806 800
rect 39118 0 39174 800
rect 39486 0 39542 800
rect 39854 0 39910 800
rect 40222 0 40278 800
rect 40590 0 40646 800
rect 40958 0 41014 800
rect 41326 0 41382 800
rect 41694 0 41750 800
rect 42062 0 42118 800
rect 42430 0 42486 800
rect 42798 0 42854 800
rect 43166 0 43222 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44270 0 44326 800
rect 44638 0 44694 800
rect 45006 0 45062 800
rect 45374 0 45430 800
rect 45742 0 45798 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46846 0 46902 800
rect 47214 0 47270 800
rect 47582 0 47638 800
rect 47950 0 48006 800
rect 48318 0 48374 800
rect 48686 0 48742 800
rect 49054 0 49110 800
rect 49422 0 49478 800
rect 49790 0 49846 800
rect 50158 0 50214 800
rect 50526 0 50582 800
rect 50894 0 50950 800
rect 51262 0 51318 800
rect 51630 0 51686 800
rect 51998 0 52054 800
rect 52366 0 52422 800
rect 52734 0 52790 800
rect 53102 0 53158 800
rect 53470 0 53526 800
rect 53838 0 53894 800
rect 54206 0 54262 800
rect 54574 0 54630 800
rect 54942 0 54998 800
rect 55310 0 55366 800
rect 55678 0 55734 800
rect 56046 0 56102 800
rect 56414 0 56470 800
rect 56782 0 56838 800
rect 57150 0 57206 800
rect 57518 0 57574 800
rect 57886 0 57942 800
rect 58254 0 58310 800
rect 58622 0 58678 800
rect 58990 0 59046 800
rect 59358 0 59414 800
rect 59726 0 59782 800
rect 60094 0 60150 800
rect 60462 0 60518 800
rect 60830 0 60886 800
rect 61198 0 61254 800
rect 61566 0 61622 800
rect 61934 0 61990 800
rect 62302 0 62358 800
rect 62670 0 62726 800
rect 63038 0 63094 800
rect 63406 0 63462 800
rect 63774 0 63830 800
rect 64142 0 64198 800
rect 64510 0 64566 800
rect 64878 0 64934 800
rect 65246 0 65302 800
rect 65614 0 65670 800
rect 65982 0 66038 800
rect 66350 0 66406 800
rect 66718 0 66774 800
rect 67086 0 67142 800
rect 67454 0 67510 800
rect 67822 0 67878 800
rect 68190 0 68246 800
rect 68558 0 68614 800
rect 68926 0 68982 800
rect 69294 0 69350 800
rect 69662 0 69718 800
rect 70030 0 70086 800
rect 70398 0 70454 800
rect 70766 0 70822 800
rect 71134 0 71190 800
rect 71502 0 71558 800
rect 71870 0 71926 800
rect 72238 0 72294 800
rect 72606 0 72662 800
rect 72974 0 73030 800
rect 73342 0 73398 800
rect 73710 0 73766 800
rect 74078 0 74134 800
rect 74446 0 74502 800
rect 74814 0 74870 800
rect 75182 0 75238 800
rect 75550 0 75606 800
rect 75918 0 75974 800
rect 76286 0 76342 800
rect 76654 0 76710 800
rect 77022 0 77078 800
rect 77390 0 77446 800
rect 77758 0 77814 800
rect 78126 0 78182 800
rect 78494 0 78550 800
rect 78862 0 78918 800
rect 79230 0 79286 800
rect 79598 0 79654 800
rect 79966 0 80022 800
rect 80334 0 80390 800
rect 80702 0 80758 800
rect 81070 0 81126 800
rect 81438 0 81494 800
rect 81806 0 81862 800
rect 82174 0 82230 800
rect 82542 0 82598 800
rect 82910 0 82966 800
rect 83278 0 83334 800
rect 83646 0 83702 800
rect 84014 0 84070 800
rect 84382 0 84438 800
rect 84750 0 84806 800
rect 85118 0 85174 800
rect 85486 0 85542 800
rect 85854 0 85910 800
rect 86222 0 86278 800
rect 86590 0 86646 800
rect 86958 0 87014 800
rect 87326 0 87382 800
rect 87694 0 87750 800
rect 88062 0 88118 800
rect 88430 0 88486 800
rect 88798 0 88854 800
rect 89166 0 89222 800
rect 89534 0 89590 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90638 0 90694 800
rect 91006 0 91062 800
rect 91374 0 91430 800
rect 91742 0 91798 800
rect 92110 0 92166 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93214 0 93270 800
rect 93582 0 93638 800
rect 93950 0 94006 800
rect 94318 0 94374 800
rect 94686 0 94742 800
rect 95054 0 95110 800
rect 95422 0 95478 800
rect 95790 0 95846 800
rect 96158 0 96214 800
rect 96526 0 96582 800
rect 96894 0 96950 800
rect 97262 0 97318 800
rect 97630 0 97686 800
rect 97998 0 98054 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99102 0 99158 800
rect 99470 0 99526 800
rect 99838 0 99894 800
rect 100206 0 100262 800
rect 100574 0 100630 800
rect 100942 0 100998 800
rect 101310 0 101366 800
rect 101678 0 101734 800
rect 102046 0 102102 800
rect 102414 0 102470 800
rect 102782 0 102838 800
rect 103150 0 103206 800
rect 103518 0 103574 800
rect 103886 0 103942 800
rect 104254 0 104310 800
rect 104622 0 104678 800
rect 104990 0 105046 800
rect 105358 0 105414 800
rect 105726 0 105782 800
rect 106094 0 106150 800
rect 106462 0 106518 800
rect 106830 0 106886 800
rect 107198 0 107254 800
rect 107566 0 107622 800
rect 107934 0 107990 800
rect 108302 0 108358 800
rect 108670 0 108726 800
rect 109038 0 109094 800
rect 109406 0 109462 800
rect 109774 0 109830 800
rect 110142 0 110198 800
rect 110510 0 110566 800
rect 110878 0 110934 800
rect 111246 0 111302 800
rect 111614 0 111670 800
rect 111982 0 112038 800
rect 112350 0 112406 800
rect 112718 0 112774 800
rect 113086 0 113142 800
<< obsm2 >>
rect 110 856 119122 87718
rect 110 2 6678 856
rect 6846 2 7046 856
rect 7214 2 7414 856
rect 7582 2 7782 856
rect 7950 2 8150 856
rect 8318 2 8518 856
rect 8686 2 8886 856
rect 9054 2 9254 856
rect 9422 2 9622 856
rect 9790 2 9990 856
rect 10158 2 10358 856
rect 10526 2 10726 856
rect 10894 2 11094 856
rect 11262 2 11462 856
rect 11630 2 11830 856
rect 11998 2 12198 856
rect 12366 2 12566 856
rect 12734 2 12934 856
rect 13102 2 13302 856
rect 13470 2 13670 856
rect 13838 2 14038 856
rect 14206 2 14406 856
rect 14574 2 14774 856
rect 14942 2 15142 856
rect 15310 2 15510 856
rect 15678 2 15878 856
rect 16046 2 16246 856
rect 16414 2 16614 856
rect 16782 2 16982 856
rect 17150 2 17350 856
rect 17518 2 17718 856
rect 17886 2 18086 856
rect 18254 2 18454 856
rect 18622 2 18822 856
rect 18990 2 19190 856
rect 19358 2 19558 856
rect 19726 2 19926 856
rect 20094 2 20294 856
rect 20462 2 20662 856
rect 20830 2 21030 856
rect 21198 2 21398 856
rect 21566 2 21766 856
rect 21934 2 22134 856
rect 22302 2 22502 856
rect 22670 2 22870 856
rect 23038 2 23238 856
rect 23406 2 23606 856
rect 23774 2 23974 856
rect 24142 2 24342 856
rect 24510 2 24710 856
rect 24878 2 25078 856
rect 25246 2 25446 856
rect 25614 2 25814 856
rect 25982 2 26182 856
rect 26350 2 26550 856
rect 26718 2 26918 856
rect 27086 2 27286 856
rect 27454 2 27654 856
rect 27822 2 28022 856
rect 28190 2 28390 856
rect 28558 2 28758 856
rect 28926 2 29126 856
rect 29294 2 29494 856
rect 29662 2 29862 856
rect 30030 2 30230 856
rect 30398 2 30598 856
rect 30766 2 30966 856
rect 31134 2 31334 856
rect 31502 2 31702 856
rect 31870 2 32070 856
rect 32238 2 32438 856
rect 32606 2 32806 856
rect 32974 2 33174 856
rect 33342 2 33542 856
rect 33710 2 33910 856
rect 34078 2 34278 856
rect 34446 2 34646 856
rect 34814 2 35014 856
rect 35182 2 35382 856
rect 35550 2 35750 856
rect 35918 2 36118 856
rect 36286 2 36486 856
rect 36654 2 36854 856
rect 37022 2 37222 856
rect 37390 2 37590 856
rect 37758 2 37958 856
rect 38126 2 38326 856
rect 38494 2 38694 856
rect 38862 2 39062 856
rect 39230 2 39430 856
rect 39598 2 39798 856
rect 39966 2 40166 856
rect 40334 2 40534 856
rect 40702 2 40902 856
rect 41070 2 41270 856
rect 41438 2 41638 856
rect 41806 2 42006 856
rect 42174 2 42374 856
rect 42542 2 42742 856
rect 42910 2 43110 856
rect 43278 2 43478 856
rect 43646 2 43846 856
rect 44014 2 44214 856
rect 44382 2 44582 856
rect 44750 2 44950 856
rect 45118 2 45318 856
rect 45486 2 45686 856
rect 45854 2 46054 856
rect 46222 2 46422 856
rect 46590 2 46790 856
rect 46958 2 47158 856
rect 47326 2 47526 856
rect 47694 2 47894 856
rect 48062 2 48262 856
rect 48430 2 48630 856
rect 48798 2 48998 856
rect 49166 2 49366 856
rect 49534 2 49734 856
rect 49902 2 50102 856
rect 50270 2 50470 856
rect 50638 2 50838 856
rect 51006 2 51206 856
rect 51374 2 51574 856
rect 51742 2 51942 856
rect 52110 2 52310 856
rect 52478 2 52678 856
rect 52846 2 53046 856
rect 53214 2 53414 856
rect 53582 2 53782 856
rect 53950 2 54150 856
rect 54318 2 54518 856
rect 54686 2 54886 856
rect 55054 2 55254 856
rect 55422 2 55622 856
rect 55790 2 55990 856
rect 56158 2 56358 856
rect 56526 2 56726 856
rect 56894 2 57094 856
rect 57262 2 57462 856
rect 57630 2 57830 856
rect 57998 2 58198 856
rect 58366 2 58566 856
rect 58734 2 58934 856
rect 59102 2 59302 856
rect 59470 2 59670 856
rect 59838 2 60038 856
rect 60206 2 60406 856
rect 60574 2 60774 856
rect 60942 2 61142 856
rect 61310 2 61510 856
rect 61678 2 61878 856
rect 62046 2 62246 856
rect 62414 2 62614 856
rect 62782 2 62982 856
rect 63150 2 63350 856
rect 63518 2 63718 856
rect 63886 2 64086 856
rect 64254 2 64454 856
rect 64622 2 64822 856
rect 64990 2 65190 856
rect 65358 2 65558 856
rect 65726 2 65926 856
rect 66094 2 66294 856
rect 66462 2 66662 856
rect 66830 2 67030 856
rect 67198 2 67398 856
rect 67566 2 67766 856
rect 67934 2 68134 856
rect 68302 2 68502 856
rect 68670 2 68870 856
rect 69038 2 69238 856
rect 69406 2 69606 856
rect 69774 2 69974 856
rect 70142 2 70342 856
rect 70510 2 70710 856
rect 70878 2 71078 856
rect 71246 2 71446 856
rect 71614 2 71814 856
rect 71982 2 72182 856
rect 72350 2 72550 856
rect 72718 2 72918 856
rect 73086 2 73286 856
rect 73454 2 73654 856
rect 73822 2 74022 856
rect 74190 2 74390 856
rect 74558 2 74758 856
rect 74926 2 75126 856
rect 75294 2 75494 856
rect 75662 2 75862 856
rect 76030 2 76230 856
rect 76398 2 76598 856
rect 76766 2 76966 856
rect 77134 2 77334 856
rect 77502 2 77702 856
rect 77870 2 78070 856
rect 78238 2 78438 856
rect 78606 2 78806 856
rect 78974 2 79174 856
rect 79342 2 79542 856
rect 79710 2 79910 856
rect 80078 2 80278 856
rect 80446 2 80646 856
rect 80814 2 81014 856
rect 81182 2 81382 856
rect 81550 2 81750 856
rect 81918 2 82118 856
rect 82286 2 82486 856
rect 82654 2 82854 856
rect 83022 2 83222 856
rect 83390 2 83590 856
rect 83758 2 83958 856
rect 84126 2 84326 856
rect 84494 2 84694 856
rect 84862 2 85062 856
rect 85230 2 85430 856
rect 85598 2 85798 856
rect 85966 2 86166 856
rect 86334 2 86534 856
rect 86702 2 86902 856
rect 87070 2 87270 856
rect 87438 2 87638 856
rect 87806 2 88006 856
rect 88174 2 88374 856
rect 88542 2 88742 856
rect 88910 2 89110 856
rect 89278 2 89478 856
rect 89646 2 89846 856
rect 90014 2 90214 856
rect 90382 2 90582 856
rect 90750 2 90950 856
rect 91118 2 91318 856
rect 91486 2 91686 856
rect 91854 2 92054 856
rect 92222 2 92422 856
rect 92590 2 92790 856
rect 92958 2 93158 856
rect 93326 2 93526 856
rect 93694 2 93894 856
rect 94062 2 94262 856
rect 94430 2 94630 856
rect 94798 2 94998 856
rect 95166 2 95366 856
rect 95534 2 95734 856
rect 95902 2 96102 856
rect 96270 2 96470 856
rect 96638 2 96838 856
rect 97006 2 97206 856
rect 97374 2 97574 856
rect 97742 2 97942 856
rect 98110 2 98310 856
rect 98478 2 98678 856
rect 98846 2 99046 856
rect 99214 2 99414 856
rect 99582 2 99782 856
rect 99950 2 100150 856
rect 100318 2 100518 856
rect 100686 2 100886 856
rect 101054 2 101254 856
rect 101422 2 101622 856
rect 101790 2 101990 856
rect 102158 2 102358 856
rect 102526 2 102726 856
rect 102894 2 103094 856
rect 103262 2 103462 856
rect 103630 2 103830 856
rect 103998 2 104198 856
rect 104366 2 104566 856
rect 104734 2 104934 856
rect 105102 2 105302 856
rect 105470 2 105670 856
rect 105838 2 106038 856
rect 106206 2 106406 856
rect 106574 2 106774 856
rect 106942 2 107142 856
rect 107310 2 107510 856
rect 107678 2 107878 856
rect 108046 2 108246 856
rect 108414 2 108614 856
rect 108782 2 108982 856
rect 109150 2 109350 856
rect 109518 2 109718 856
rect 109886 2 110086 856
rect 110254 2 110454 856
rect 110622 2 110822 856
rect 110990 2 111190 856
rect 111358 2 111558 856
rect 111726 2 111926 856
rect 112094 2 112294 856
rect 112462 2 112662 856
rect 112830 2 113030 856
rect 113198 2 119122 856
<< metal3 >>
rect 0 76440 800 76560
rect 119200 76440 120000 76560
rect 0 75896 800 76016
rect 119200 75896 120000 76016
rect 0 75352 800 75472
rect 119200 75352 120000 75472
rect 0 74808 800 74928
rect 119200 74808 120000 74928
rect 0 74264 800 74384
rect 119200 74264 120000 74384
rect 0 73720 800 73840
rect 119200 73720 120000 73840
rect 0 73176 800 73296
rect 119200 73176 120000 73296
rect 0 72632 800 72752
rect 119200 72632 120000 72752
rect 0 72088 800 72208
rect 119200 72088 120000 72208
rect 0 71544 800 71664
rect 119200 71544 120000 71664
rect 0 71000 800 71120
rect 119200 71000 120000 71120
rect 0 70456 800 70576
rect 119200 70456 120000 70576
rect 0 69912 800 70032
rect 119200 69912 120000 70032
rect 0 69368 800 69488
rect 119200 69368 120000 69488
rect 0 68824 800 68944
rect 119200 68824 120000 68944
rect 0 68280 800 68400
rect 119200 68280 120000 68400
rect 0 67736 800 67856
rect 119200 67736 120000 67856
rect 0 67192 800 67312
rect 119200 67192 120000 67312
rect 0 66648 800 66768
rect 119200 66648 120000 66768
rect 0 66104 800 66224
rect 119200 66104 120000 66224
rect 0 65560 800 65680
rect 119200 65560 120000 65680
rect 0 65016 800 65136
rect 119200 65016 120000 65136
rect 0 64472 800 64592
rect 119200 64472 120000 64592
rect 0 63928 800 64048
rect 119200 63928 120000 64048
rect 0 63384 800 63504
rect 119200 63384 120000 63504
rect 0 62840 800 62960
rect 119200 62840 120000 62960
rect 0 62296 800 62416
rect 119200 62296 120000 62416
rect 0 61752 800 61872
rect 119200 61752 120000 61872
rect 0 61208 800 61328
rect 119200 61208 120000 61328
rect 0 60664 800 60784
rect 119200 60664 120000 60784
rect 0 60120 800 60240
rect 119200 60120 120000 60240
rect 0 59576 800 59696
rect 119200 59576 120000 59696
rect 0 59032 800 59152
rect 119200 59032 120000 59152
rect 0 58488 800 58608
rect 119200 58488 120000 58608
rect 0 57944 800 58064
rect 119200 57944 120000 58064
rect 0 57400 800 57520
rect 119200 57400 120000 57520
rect 0 56856 800 56976
rect 119200 56856 120000 56976
rect 0 56312 800 56432
rect 119200 56312 120000 56432
rect 0 55768 800 55888
rect 119200 55768 120000 55888
rect 0 55224 800 55344
rect 119200 55224 120000 55344
rect 0 54680 800 54800
rect 119200 54680 120000 54800
rect 0 54136 800 54256
rect 119200 54136 120000 54256
rect 0 53592 800 53712
rect 119200 53592 120000 53712
rect 0 53048 800 53168
rect 119200 53048 120000 53168
rect 0 52504 800 52624
rect 119200 52504 120000 52624
rect 0 51960 800 52080
rect 119200 51960 120000 52080
rect 0 51416 800 51536
rect 119200 51416 120000 51536
rect 0 50872 800 50992
rect 119200 50872 120000 50992
rect 0 50328 800 50448
rect 119200 50328 120000 50448
rect 0 49784 800 49904
rect 119200 49784 120000 49904
rect 0 49240 800 49360
rect 119200 49240 120000 49360
rect 0 48696 800 48816
rect 119200 48696 120000 48816
rect 0 48152 800 48272
rect 119200 48152 120000 48272
rect 0 47608 800 47728
rect 119200 47608 120000 47728
rect 0 47064 800 47184
rect 119200 47064 120000 47184
rect 0 46520 800 46640
rect 119200 46520 120000 46640
rect 0 45976 800 46096
rect 119200 45976 120000 46096
rect 0 45432 800 45552
rect 119200 45432 120000 45552
rect 0 44888 800 45008
rect 119200 44888 120000 45008
rect 0 44344 800 44464
rect 119200 44344 120000 44464
rect 0 43800 800 43920
rect 119200 43800 120000 43920
rect 0 43256 800 43376
rect 119200 43256 120000 43376
rect 0 42712 800 42832
rect 119200 42712 120000 42832
rect 0 42168 800 42288
rect 119200 42168 120000 42288
rect 0 41624 800 41744
rect 119200 41624 120000 41744
rect 0 41080 800 41200
rect 119200 41080 120000 41200
rect 0 40536 800 40656
rect 119200 40536 120000 40656
rect 0 39992 800 40112
rect 119200 39992 120000 40112
rect 0 39448 800 39568
rect 119200 39448 120000 39568
rect 0 38904 800 39024
rect 119200 38904 120000 39024
rect 0 38360 800 38480
rect 119200 38360 120000 38480
rect 0 37816 800 37936
rect 119200 37816 120000 37936
rect 0 37272 800 37392
rect 119200 37272 120000 37392
rect 0 36728 800 36848
rect 119200 36728 120000 36848
rect 0 36184 800 36304
rect 119200 36184 120000 36304
rect 0 35640 800 35760
rect 119200 35640 120000 35760
rect 0 35096 800 35216
rect 119200 35096 120000 35216
rect 0 34552 800 34672
rect 119200 34552 120000 34672
rect 0 34008 800 34128
rect 119200 34008 120000 34128
rect 0 33464 800 33584
rect 119200 33464 120000 33584
rect 0 32920 800 33040
rect 119200 32920 120000 33040
rect 0 32376 800 32496
rect 119200 32376 120000 32496
rect 0 31832 800 31952
rect 119200 31832 120000 31952
rect 0 31288 800 31408
rect 119200 31288 120000 31408
rect 0 30744 800 30864
rect 119200 30744 120000 30864
rect 0 30200 800 30320
rect 119200 30200 120000 30320
rect 0 29656 800 29776
rect 119200 29656 120000 29776
rect 0 29112 800 29232
rect 119200 29112 120000 29232
rect 0 28568 800 28688
rect 119200 28568 120000 28688
rect 0 28024 800 28144
rect 119200 28024 120000 28144
rect 0 27480 800 27600
rect 119200 27480 120000 27600
rect 0 26936 800 27056
rect 119200 26936 120000 27056
rect 0 26392 800 26512
rect 119200 26392 120000 26512
rect 0 25848 800 25968
rect 119200 25848 120000 25968
rect 0 25304 800 25424
rect 119200 25304 120000 25424
rect 0 24760 800 24880
rect 119200 24760 120000 24880
rect 0 24216 800 24336
rect 119200 24216 120000 24336
rect 0 23672 800 23792
rect 119200 23672 120000 23792
rect 0 23128 800 23248
rect 119200 23128 120000 23248
rect 0 22584 800 22704
rect 119200 22584 120000 22704
rect 0 22040 800 22160
rect 119200 22040 120000 22160
rect 0 21496 800 21616
rect 119200 21496 120000 21616
rect 0 20952 800 21072
rect 119200 20952 120000 21072
rect 0 20408 800 20528
rect 119200 20408 120000 20528
rect 0 19864 800 19984
rect 119200 19864 120000 19984
rect 0 19320 800 19440
rect 119200 19320 120000 19440
rect 0 18776 800 18896
rect 119200 18776 120000 18896
rect 0 18232 800 18352
rect 119200 18232 120000 18352
rect 0 17688 800 17808
rect 119200 17688 120000 17808
rect 0 17144 800 17264
rect 119200 17144 120000 17264
rect 0 16600 800 16720
rect 119200 16600 120000 16720
rect 0 16056 800 16176
rect 119200 16056 120000 16176
rect 0 15512 800 15632
rect 119200 15512 120000 15632
rect 0 14968 800 15088
rect 119200 14968 120000 15088
rect 0 14424 800 14544
rect 119200 14424 120000 14544
rect 0 13880 800 14000
rect 119200 13880 120000 14000
rect 0 13336 800 13456
rect 119200 13336 120000 13456
<< obsm3 >>
rect 105 76640 119200 87617
rect 880 76360 119120 76640
rect 105 76096 119200 76360
rect 880 75816 119120 76096
rect 105 75552 119200 75816
rect 880 75272 119120 75552
rect 105 75008 119200 75272
rect 880 74728 119120 75008
rect 105 74464 119200 74728
rect 880 74184 119120 74464
rect 105 73920 119200 74184
rect 880 73640 119120 73920
rect 105 73376 119200 73640
rect 880 73096 119120 73376
rect 105 72832 119200 73096
rect 880 72552 119120 72832
rect 105 72288 119200 72552
rect 880 72008 119120 72288
rect 105 71744 119200 72008
rect 880 71464 119120 71744
rect 105 71200 119200 71464
rect 880 70920 119120 71200
rect 105 70656 119200 70920
rect 880 70376 119120 70656
rect 105 70112 119200 70376
rect 880 69832 119120 70112
rect 105 69568 119200 69832
rect 880 69288 119120 69568
rect 105 69024 119200 69288
rect 880 68744 119120 69024
rect 105 68480 119200 68744
rect 880 68200 119120 68480
rect 105 67936 119200 68200
rect 880 67656 119120 67936
rect 105 67392 119200 67656
rect 880 67112 119120 67392
rect 105 66848 119200 67112
rect 880 66568 119120 66848
rect 105 66304 119200 66568
rect 880 66024 119120 66304
rect 105 65760 119200 66024
rect 880 65480 119120 65760
rect 105 65216 119200 65480
rect 880 64936 119120 65216
rect 105 64672 119200 64936
rect 880 64392 119120 64672
rect 105 64128 119200 64392
rect 880 63848 119120 64128
rect 105 63584 119200 63848
rect 880 63304 119120 63584
rect 105 63040 119200 63304
rect 880 62760 119120 63040
rect 105 62496 119200 62760
rect 880 62216 119120 62496
rect 105 61952 119200 62216
rect 880 61672 119120 61952
rect 105 61408 119200 61672
rect 880 61128 119120 61408
rect 105 60864 119200 61128
rect 880 60584 119120 60864
rect 105 60320 119200 60584
rect 880 60040 119120 60320
rect 105 59776 119200 60040
rect 880 59496 119120 59776
rect 105 59232 119200 59496
rect 880 58952 119120 59232
rect 105 58688 119200 58952
rect 880 58408 119120 58688
rect 105 58144 119200 58408
rect 880 57864 119120 58144
rect 105 57600 119200 57864
rect 880 57320 119120 57600
rect 105 57056 119200 57320
rect 880 56776 119120 57056
rect 105 56512 119200 56776
rect 880 56232 119120 56512
rect 105 55968 119200 56232
rect 880 55688 119120 55968
rect 105 55424 119200 55688
rect 880 55144 119120 55424
rect 105 54880 119200 55144
rect 880 54600 119120 54880
rect 105 54336 119200 54600
rect 880 54056 119120 54336
rect 105 53792 119200 54056
rect 880 53512 119120 53792
rect 105 53248 119200 53512
rect 880 52968 119120 53248
rect 105 52704 119200 52968
rect 880 52424 119120 52704
rect 105 52160 119200 52424
rect 880 51880 119120 52160
rect 105 51616 119200 51880
rect 880 51336 119120 51616
rect 105 51072 119200 51336
rect 880 50792 119120 51072
rect 105 50528 119200 50792
rect 880 50248 119120 50528
rect 105 49984 119200 50248
rect 880 49704 119120 49984
rect 105 49440 119200 49704
rect 880 49160 119120 49440
rect 105 48896 119200 49160
rect 880 48616 119120 48896
rect 105 48352 119200 48616
rect 880 48072 119120 48352
rect 105 47808 119200 48072
rect 880 47528 119120 47808
rect 105 47264 119200 47528
rect 880 46984 119120 47264
rect 105 46720 119200 46984
rect 880 46440 119120 46720
rect 105 46176 119200 46440
rect 880 45896 119120 46176
rect 105 45632 119200 45896
rect 880 45352 119120 45632
rect 105 45088 119200 45352
rect 880 44808 119120 45088
rect 105 44544 119200 44808
rect 880 44264 119120 44544
rect 105 44000 119200 44264
rect 880 43720 119120 44000
rect 105 43456 119200 43720
rect 880 43176 119120 43456
rect 105 42912 119200 43176
rect 880 42632 119120 42912
rect 105 42368 119200 42632
rect 880 42088 119120 42368
rect 105 41824 119200 42088
rect 880 41544 119120 41824
rect 105 41280 119200 41544
rect 880 41000 119120 41280
rect 105 40736 119200 41000
rect 880 40456 119120 40736
rect 105 40192 119200 40456
rect 880 39912 119120 40192
rect 105 39648 119200 39912
rect 880 39368 119120 39648
rect 105 39104 119200 39368
rect 880 38824 119120 39104
rect 105 38560 119200 38824
rect 880 38280 119120 38560
rect 105 38016 119200 38280
rect 880 37736 119120 38016
rect 105 37472 119200 37736
rect 880 37192 119120 37472
rect 105 36928 119200 37192
rect 880 36648 119120 36928
rect 105 36384 119200 36648
rect 880 36104 119120 36384
rect 105 35840 119200 36104
rect 880 35560 119120 35840
rect 105 35296 119200 35560
rect 880 35016 119120 35296
rect 105 34752 119200 35016
rect 880 34472 119120 34752
rect 105 34208 119200 34472
rect 880 33928 119120 34208
rect 105 33664 119200 33928
rect 880 33384 119120 33664
rect 105 33120 119200 33384
rect 880 32840 119120 33120
rect 105 32576 119200 32840
rect 880 32296 119120 32576
rect 105 32032 119200 32296
rect 880 31752 119120 32032
rect 105 31488 119200 31752
rect 880 31208 119120 31488
rect 105 30944 119200 31208
rect 880 30664 119120 30944
rect 105 30400 119200 30664
rect 880 30120 119120 30400
rect 105 29856 119200 30120
rect 880 29576 119120 29856
rect 105 29312 119200 29576
rect 880 29032 119120 29312
rect 105 28768 119200 29032
rect 880 28488 119120 28768
rect 105 28224 119200 28488
rect 880 27944 119120 28224
rect 105 27680 119200 27944
rect 880 27400 119120 27680
rect 105 27136 119200 27400
rect 880 26856 119120 27136
rect 105 26592 119200 26856
rect 880 26312 119120 26592
rect 105 26048 119200 26312
rect 880 25768 119120 26048
rect 105 25504 119200 25768
rect 880 25224 119120 25504
rect 105 24960 119200 25224
rect 880 24680 119120 24960
rect 105 24416 119200 24680
rect 880 24136 119120 24416
rect 105 23872 119200 24136
rect 880 23592 119120 23872
rect 105 23328 119200 23592
rect 880 23048 119120 23328
rect 105 22784 119200 23048
rect 880 22504 119120 22784
rect 105 22240 119200 22504
rect 880 21960 119120 22240
rect 105 21696 119200 21960
rect 880 21416 119120 21696
rect 105 21152 119200 21416
rect 880 20872 119120 21152
rect 105 20608 119200 20872
rect 880 20328 119120 20608
rect 105 20064 119200 20328
rect 880 19784 119120 20064
rect 105 19520 119200 19784
rect 880 19240 119120 19520
rect 105 18976 119200 19240
rect 880 18696 119120 18976
rect 105 18432 119200 18696
rect 880 18152 119120 18432
rect 105 17888 119200 18152
rect 880 17608 119120 17888
rect 105 17344 119200 17608
rect 880 17064 119120 17344
rect 105 16800 119200 17064
rect 880 16520 119120 16800
rect 105 16256 119200 16520
rect 880 15976 119120 16256
rect 105 15712 119200 15976
rect 880 15432 119120 15712
rect 105 15168 119200 15432
rect 880 14888 119120 15168
rect 105 14624 119200 14888
rect 880 14344 119120 14624
rect 105 14080 119200 14344
rect 880 13800 119120 14080
rect 105 13536 119200 13800
rect 880 13256 119120 13536
rect 105 35 119200 13256
<< metal4 >>
rect 4208 2128 4528 87632
rect 19568 2128 19888 87632
rect 34928 2128 35248 87632
rect 50288 2128 50608 87632
rect 65648 2128 65968 87632
rect 81008 2128 81328 87632
rect 96368 2128 96688 87632
rect 111728 2128 112048 87632
<< obsm4 >>
rect 611 2048 4128 80613
rect 4608 2048 19488 80613
rect 19968 2048 34848 80613
rect 35328 2048 50208 80613
rect 50688 2048 65568 80613
rect 66048 2048 80928 80613
rect 81408 2048 96288 80613
rect 96768 2048 111648 80613
rect 112128 2048 114941 80613
rect 611 171 114941 2048
<< labels >>
rlabel metal2 s 6734 0 6790 800 6 clk_i
port 1 nsew signal input
rlabel metal3 s 119200 13336 120000 13456 6 mstream_i
port 2 nsew signal input
rlabel metal3 s 119200 13880 120000 14000 6 mstream_o[0]
port 3 nsew signal output
rlabel metal3 s 119200 68280 120000 68400 6 mstream_o[100]
port 4 nsew signal output
rlabel metal3 s 119200 68824 120000 68944 6 mstream_o[101]
port 5 nsew signal output
rlabel metal3 s 119200 69368 120000 69488 6 mstream_o[102]
port 6 nsew signal output
rlabel metal3 s 119200 69912 120000 70032 6 mstream_o[103]
port 7 nsew signal output
rlabel metal3 s 119200 70456 120000 70576 6 mstream_o[104]
port 8 nsew signal output
rlabel metal3 s 119200 71000 120000 71120 6 mstream_o[105]
port 9 nsew signal output
rlabel metal3 s 119200 71544 120000 71664 6 mstream_o[106]
port 10 nsew signal output
rlabel metal3 s 119200 72088 120000 72208 6 mstream_o[107]
port 11 nsew signal output
rlabel metal3 s 119200 72632 120000 72752 6 mstream_o[108]
port 12 nsew signal output
rlabel metal3 s 119200 73176 120000 73296 6 mstream_o[109]
port 13 nsew signal output
rlabel metal3 s 119200 19320 120000 19440 6 mstream_o[10]
port 14 nsew signal output
rlabel metal3 s 119200 73720 120000 73840 6 mstream_o[110]
port 15 nsew signal output
rlabel metal3 s 119200 74264 120000 74384 6 mstream_o[111]
port 16 nsew signal output
rlabel metal3 s 119200 74808 120000 74928 6 mstream_o[112]
port 17 nsew signal output
rlabel metal3 s 119200 75352 120000 75472 6 mstream_o[113]
port 18 nsew signal output
rlabel metal3 s 119200 75896 120000 76016 6 mstream_o[114]
port 19 nsew signal output
rlabel metal3 s 119200 76440 120000 76560 6 mstream_o[115]
port 20 nsew signal output
rlabel metal3 s 119200 19864 120000 19984 6 mstream_o[11]
port 21 nsew signal output
rlabel metal3 s 119200 20408 120000 20528 6 mstream_o[12]
port 22 nsew signal output
rlabel metal3 s 119200 20952 120000 21072 6 mstream_o[13]
port 23 nsew signal output
rlabel metal3 s 119200 21496 120000 21616 6 mstream_o[14]
port 24 nsew signal output
rlabel metal3 s 119200 22040 120000 22160 6 mstream_o[15]
port 25 nsew signal output
rlabel metal3 s 119200 22584 120000 22704 6 mstream_o[16]
port 26 nsew signal output
rlabel metal3 s 119200 23128 120000 23248 6 mstream_o[17]
port 27 nsew signal output
rlabel metal3 s 119200 23672 120000 23792 6 mstream_o[18]
port 28 nsew signal output
rlabel metal3 s 119200 24216 120000 24336 6 mstream_o[19]
port 29 nsew signal output
rlabel metal3 s 119200 14424 120000 14544 6 mstream_o[1]
port 30 nsew signal output
rlabel metal3 s 119200 24760 120000 24880 6 mstream_o[20]
port 31 nsew signal output
rlabel metal3 s 119200 25304 120000 25424 6 mstream_o[21]
port 32 nsew signal output
rlabel metal3 s 119200 25848 120000 25968 6 mstream_o[22]
port 33 nsew signal output
rlabel metal3 s 119200 26392 120000 26512 6 mstream_o[23]
port 34 nsew signal output
rlabel metal3 s 119200 26936 120000 27056 6 mstream_o[24]
port 35 nsew signal output
rlabel metal3 s 119200 27480 120000 27600 6 mstream_o[25]
port 36 nsew signal output
rlabel metal3 s 119200 28024 120000 28144 6 mstream_o[26]
port 37 nsew signal output
rlabel metal3 s 119200 28568 120000 28688 6 mstream_o[27]
port 38 nsew signal output
rlabel metal3 s 119200 29112 120000 29232 6 mstream_o[28]
port 39 nsew signal output
rlabel metal3 s 119200 29656 120000 29776 6 mstream_o[29]
port 40 nsew signal output
rlabel metal3 s 119200 14968 120000 15088 6 mstream_o[2]
port 41 nsew signal output
rlabel metal3 s 119200 30200 120000 30320 6 mstream_o[30]
port 42 nsew signal output
rlabel metal3 s 119200 30744 120000 30864 6 mstream_o[31]
port 43 nsew signal output
rlabel metal3 s 119200 31288 120000 31408 6 mstream_o[32]
port 44 nsew signal output
rlabel metal3 s 119200 31832 120000 31952 6 mstream_o[33]
port 45 nsew signal output
rlabel metal3 s 119200 32376 120000 32496 6 mstream_o[34]
port 46 nsew signal output
rlabel metal3 s 119200 32920 120000 33040 6 mstream_o[35]
port 47 nsew signal output
rlabel metal3 s 119200 33464 120000 33584 6 mstream_o[36]
port 48 nsew signal output
rlabel metal3 s 119200 34008 120000 34128 6 mstream_o[37]
port 49 nsew signal output
rlabel metal3 s 119200 34552 120000 34672 6 mstream_o[38]
port 50 nsew signal output
rlabel metal3 s 119200 35096 120000 35216 6 mstream_o[39]
port 51 nsew signal output
rlabel metal3 s 119200 15512 120000 15632 6 mstream_o[3]
port 52 nsew signal output
rlabel metal3 s 119200 35640 120000 35760 6 mstream_o[40]
port 53 nsew signal output
rlabel metal3 s 119200 36184 120000 36304 6 mstream_o[41]
port 54 nsew signal output
rlabel metal3 s 119200 36728 120000 36848 6 mstream_o[42]
port 55 nsew signal output
rlabel metal3 s 119200 37272 120000 37392 6 mstream_o[43]
port 56 nsew signal output
rlabel metal3 s 119200 37816 120000 37936 6 mstream_o[44]
port 57 nsew signal output
rlabel metal3 s 119200 38360 120000 38480 6 mstream_o[45]
port 58 nsew signal output
rlabel metal3 s 119200 38904 120000 39024 6 mstream_o[46]
port 59 nsew signal output
rlabel metal3 s 119200 39448 120000 39568 6 mstream_o[47]
port 60 nsew signal output
rlabel metal3 s 119200 39992 120000 40112 6 mstream_o[48]
port 61 nsew signal output
rlabel metal3 s 119200 40536 120000 40656 6 mstream_o[49]
port 62 nsew signal output
rlabel metal3 s 119200 16056 120000 16176 6 mstream_o[4]
port 63 nsew signal output
rlabel metal3 s 119200 41080 120000 41200 6 mstream_o[50]
port 64 nsew signal output
rlabel metal3 s 119200 41624 120000 41744 6 mstream_o[51]
port 65 nsew signal output
rlabel metal3 s 119200 42168 120000 42288 6 mstream_o[52]
port 66 nsew signal output
rlabel metal3 s 119200 42712 120000 42832 6 mstream_o[53]
port 67 nsew signal output
rlabel metal3 s 119200 43256 120000 43376 6 mstream_o[54]
port 68 nsew signal output
rlabel metal3 s 119200 43800 120000 43920 6 mstream_o[55]
port 69 nsew signal output
rlabel metal3 s 119200 44344 120000 44464 6 mstream_o[56]
port 70 nsew signal output
rlabel metal3 s 119200 44888 120000 45008 6 mstream_o[57]
port 71 nsew signal output
rlabel metal3 s 119200 45432 120000 45552 6 mstream_o[58]
port 72 nsew signal output
rlabel metal3 s 119200 45976 120000 46096 6 mstream_o[59]
port 73 nsew signal output
rlabel metal3 s 119200 16600 120000 16720 6 mstream_o[5]
port 74 nsew signal output
rlabel metal3 s 119200 46520 120000 46640 6 mstream_o[60]
port 75 nsew signal output
rlabel metal3 s 119200 47064 120000 47184 6 mstream_o[61]
port 76 nsew signal output
rlabel metal3 s 119200 47608 120000 47728 6 mstream_o[62]
port 77 nsew signal output
rlabel metal3 s 119200 48152 120000 48272 6 mstream_o[63]
port 78 nsew signal output
rlabel metal3 s 119200 48696 120000 48816 6 mstream_o[64]
port 79 nsew signal output
rlabel metal3 s 119200 49240 120000 49360 6 mstream_o[65]
port 80 nsew signal output
rlabel metal3 s 119200 49784 120000 49904 6 mstream_o[66]
port 81 nsew signal output
rlabel metal3 s 119200 50328 120000 50448 6 mstream_o[67]
port 82 nsew signal output
rlabel metal3 s 119200 50872 120000 50992 6 mstream_o[68]
port 83 nsew signal output
rlabel metal3 s 119200 51416 120000 51536 6 mstream_o[69]
port 84 nsew signal output
rlabel metal3 s 119200 17144 120000 17264 6 mstream_o[6]
port 85 nsew signal output
rlabel metal3 s 119200 51960 120000 52080 6 mstream_o[70]
port 86 nsew signal output
rlabel metal3 s 119200 52504 120000 52624 6 mstream_o[71]
port 87 nsew signal output
rlabel metal3 s 119200 53048 120000 53168 6 mstream_o[72]
port 88 nsew signal output
rlabel metal3 s 119200 53592 120000 53712 6 mstream_o[73]
port 89 nsew signal output
rlabel metal3 s 119200 54136 120000 54256 6 mstream_o[74]
port 90 nsew signal output
rlabel metal3 s 119200 54680 120000 54800 6 mstream_o[75]
port 91 nsew signal output
rlabel metal3 s 119200 55224 120000 55344 6 mstream_o[76]
port 92 nsew signal output
rlabel metal3 s 119200 55768 120000 55888 6 mstream_o[77]
port 93 nsew signal output
rlabel metal3 s 119200 56312 120000 56432 6 mstream_o[78]
port 94 nsew signal output
rlabel metal3 s 119200 56856 120000 56976 6 mstream_o[79]
port 95 nsew signal output
rlabel metal3 s 119200 17688 120000 17808 6 mstream_o[7]
port 96 nsew signal output
rlabel metal3 s 119200 57400 120000 57520 6 mstream_o[80]
port 97 nsew signal output
rlabel metal3 s 119200 57944 120000 58064 6 mstream_o[81]
port 98 nsew signal output
rlabel metal3 s 119200 58488 120000 58608 6 mstream_o[82]
port 99 nsew signal output
rlabel metal3 s 119200 59032 120000 59152 6 mstream_o[83]
port 100 nsew signal output
rlabel metal3 s 119200 59576 120000 59696 6 mstream_o[84]
port 101 nsew signal output
rlabel metal3 s 119200 60120 120000 60240 6 mstream_o[85]
port 102 nsew signal output
rlabel metal3 s 119200 60664 120000 60784 6 mstream_o[86]
port 103 nsew signal output
rlabel metal3 s 119200 61208 120000 61328 6 mstream_o[87]
port 104 nsew signal output
rlabel metal3 s 119200 61752 120000 61872 6 mstream_o[88]
port 105 nsew signal output
rlabel metal3 s 119200 62296 120000 62416 6 mstream_o[89]
port 106 nsew signal output
rlabel metal3 s 119200 18232 120000 18352 6 mstream_o[8]
port 107 nsew signal output
rlabel metal3 s 119200 62840 120000 62960 6 mstream_o[90]
port 108 nsew signal output
rlabel metal3 s 119200 63384 120000 63504 6 mstream_o[91]
port 109 nsew signal output
rlabel metal3 s 119200 63928 120000 64048 6 mstream_o[92]
port 110 nsew signal output
rlabel metal3 s 119200 64472 120000 64592 6 mstream_o[93]
port 111 nsew signal output
rlabel metal3 s 119200 65016 120000 65136 6 mstream_o[94]
port 112 nsew signal output
rlabel metal3 s 119200 65560 120000 65680 6 mstream_o[95]
port 113 nsew signal output
rlabel metal3 s 119200 66104 120000 66224 6 mstream_o[96]
port 114 nsew signal output
rlabel metal3 s 119200 66648 120000 66768 6 mstream_o[97]
port 115 nsew signal output
rlabel metal3 s 119200 67192 120000 67312 6 mstream_o[98]
port 116 nsew signal output
rlabel metal3 s 119200 67736 120000 67856 6 mstream_o[99]
port 117 nsew signal output
rlabel metal3 s 119200 18776 120000 18896 6 mstream_o[9]
port 118 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 nrst_i
port 119 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 sstream_i[0]
port 120 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 sstream_i[100]
port 121 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 sstream_i[101]
port 122 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 sstream_i[102]
port 123 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 sstream_i[103]
port 124 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 sstream_i[104]
port 125 nsew signal input
rlabel metal3 s 0 70456 800 70576 6 sstream_i[105]
port 126 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 sstream_i[106]
port 127 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 sstream_i[107]
port 128 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 sstream_i[108]
port 129 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 sstream_i[109]
port 130 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 sstream_i[10]
port 131 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 sstream_i[110]
port 132 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 sstream_i[111]
port 133 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 sstream_i[112]
port 134 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 sstream_i[113]
port 135 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 sstream_i[114]
port 136 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 sstream_i[115]
port 137 nsew signal input
rlabel metal3 s 0 19320 800 19440 6 sstream_i[11]
port 138 nsew signal input
rlabel metal3 s 0 19864 800 19984 6 sstream_i[12]
port 139 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 sstream_i[13]
port 140 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 sstream_i[14]
port 141 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 sstream_i[15]
port 142 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 sstream_i[16]
port 143 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 sstream_i[17]
port 144 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 sstream_i[18]
port 145 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 sstream_i[19]
port 146 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 sstream_i[1]
port 147 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 sstream_i[20]
port 148 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 sstream_i[21]
port 149 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 sstream_i[22]
port 150 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 sstream_i[23]
port 151 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 sstream_i[24]
port 152 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 sstream_i[25]
port 153 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 sstream_i[26]
port 154 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 sstream_i[27]
port 155 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 sstream_i[28]
port 156 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 sstream_i[29]
port 157 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 sstream_i[2]
port 158 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 sstream_i[30]
port 159 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 sstream_i[31]
port 160 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 sstream_i[32]
port 161 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 sstream_i[33]
port 162 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 sstream_i[34]
port 163 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 sstream_i[35]
port 164 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 sstream_i[36]
port 165 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 sstream_i[37]
port 166 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 sstream_i[38]
port 167 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 sstream_i[39]
port 168 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 sstream_i[3]
port 169 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 sstream_i[40]
port 170 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 sstream_i[41]
port 171 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 sstream_i[42]
port 172 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 sstream_i[43]
port 173 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 sstream_i[44]
port 174 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 sstream_i[45]
port 175 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 sstream_i[46]
port 176 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 sstream_i[47]
port 177 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 sstream_i[48]
port 178 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 sstream_i[49]
port 179 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 sstream_i[4]
port 180 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 sstream_i[50]
port 181 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 sstream_i[51]
port 182 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 sstream_i[52]
port 183 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 sstream_i[53]
port 184 nsew signal input
rlabel metal3 s 0 42712 800 42832 6 sstream_i[54]
port 185 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 sstream_i[55]
port 186 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 sstream_i[56]
port 187 nsew signal input
rlabel metal3 s 0 44344 800 44464 6 sstream_i[57]
port 188 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 sstream_i[58]
port 189 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 sstream_i[59]
port 190 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 sstream_i[5]
port 191 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 sstream_i[60]
port 192 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 sstream_i[61]
port 193 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 sstream_i[62]
port 194 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 sstream_i[63]
port 195 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 sstream_i[64]
port 196 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 sstream_i[65]
port 197 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 sstream_i[66]
port 198 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 sstream_i[67]
port 199 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 sstream_i[68]
port 200 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 sstream_i[69]
port 201 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 sstream_i[6]
port 202 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 sstream_i[70]
port 203 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 sstream_i[71]
port 204 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 sstream_i[72]
port 205 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 sstream_i[73]
port 206 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 sstream_i[74]
port 207 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 sstream_i[75]
port 208 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 sstream_i[76]
port 209 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 sstream_i[77]
port 210 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 sstream_i[78]
port 211 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 sstream_i[79]
port 212 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 sstream_i[7]
port 213 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 sstream_i[80]
port 214 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 sstream_i[81]
port 215 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 sstream_i[82]
port 216 nsew signal input
rlabel metal3 s 0 58488 800 58608 6 sstream_i[83]
port 217 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 sstream_i[84]
port 218 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 sstream_i[85]
port 219 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 sstream_i[86]
port 220 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 sstream_i[87]
port 221 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 sstream_i[88]
port 222 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 sstream_i[89]
port 223 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 sstream_i[8]
port 224 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 sstream_i[90]
port 225 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 sstream_i[91]
port 226 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 sstream_i[92]
port 227 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 sstream_i[93]
port 228 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 sstream_i[94]
port 229 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 sstream_i[95]
port 230 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 sstream_i[96]
port 231 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 sstream_i[97]
port 232 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 sstream_i[98]
port 233 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 sstream_i[99]
port 234 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 sstream_i[9]
port 235 nsew signal input
rlabel metal3 s 0 76440 800 76560 6 sstream_o
port 236 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 t0x[0]
port 237 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 t0x[10]
port 238 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 t0x[11]
port 239 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 t0x[12]
port 240 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 t0x[13]
port 241 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 t0x[14]
port 242 nsew signal input
rlabel metal2 s 75918 0 75974 800 6 t0x[15]
port 243 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 t0x[16]
port 244 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 t0x[17]
port 245 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 t0x[18]
port 246 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 t0x[19]
port 247 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 t0x[1]
port 248 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 t0x[20]
port 249 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 t0x[21]
port 250 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 t0x[22]
port 251 nsew signal input
rlabel metal2 s 93582 0 93638 800 6 t0x[23]
port 252 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 t0x[24]
port 253 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 t0x[25]
port 254 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 t0x[26]
port 255 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 t0x[27]
port 256 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 t0x[28]
port 257 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 t0x[29]
port 258 nsew signal input
rlabel metal2 s 47214 0 47270 800 6 t0x[2]
port 259 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 t0x[30]
port 260 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 t0x[31]
port 261 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 t0x[3]
port 262 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 t0x[4]
port 263 nsew signal input
rlabel metal2 s 53838 0 53894 800 6 t0x[5]
port 264 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 t0x[6]
port 265 nsew signal input
rlabel metal2 s 58254 0 58310 800 6 t0x[7]
port 266 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 t0x[8]
port 267 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 t0x[9]
port 268 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 t0y[0]
port 269 nsew signal input
rlabel metal2 s 65246 0 65302 800 6 t0y[10]
port 270 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 t0y[11]
port 271 nsew signal input
rlabel metal2 s 69662 0 69718 800 6 t0y[12]
port 272 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 t0y[13]
port 273 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 t0y[14]
port 274 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 t0y[15]
port 275 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 t0y[16]
port 276 nsew signal input
rlabel metal2 s 80702 0 80758 800 6 t0y[17]
port 277 nsew signal input
rlabel metal2 s 82910 0 82966 800 6 t0y[18]
port 278 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 t0y[19]
port 279 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 t0y[1]
port 280 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 t0y[20]
port 281 nsew signal input
rlabel metal2 s 89534 0 89590 800 6 t0y[21]
port 282 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 t0y[22]
port 283 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 t0y[23]
port 284 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 t0y[24]
port 285 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 t0y[25]
port 286 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 t0y[26]
port 287 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 t0y[27]
port 288 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 t0y[28]
port 289 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 t0y[29]
port 290 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 t0y[2]
port 291 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 t0y[30]
port 292 nsew signal input
rlabel metal2 s 111614 0 111670 800 6 t0y[31]
port 293 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 t0y[3]
port 294 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 t0y[4]
port 295 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 t0y[5]
port 296 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 t0y[6]
port 297 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 t0y[7]
port 298 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 t0y[8]
port 299 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 t0y[9]
port 300 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 t1x[0]
port 301 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 t1x[10]
port 302 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 t1x[11]
port 303 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 t1x[12]
port 304 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 t1x[13]
port 305 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 t1x[14]
port 306 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 t1x[15]
port 307 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 t1x[16]
port 308 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 t1x[17]
port 309 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 t1x[18]
port 310 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 t1x[19]
port 311 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 t1x[1]
port 312 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 t1x[20]
port 313 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 t1x[21]
port 314 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 t1x[22]
port 315 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 t1x[23]
port 316 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 t1x[24]
port 317 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 t1x[25]
port 318 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 t1x[26]
port 319 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 t1x[27]
port 320 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 t1x[28]
port 321 nsew signal input
rlabel metal2 s 107566 0 107622 800 6 t1x[29]
port 322 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 t1x[2]
port 323 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 t1x[30]
port 324 nsew signal input
rlabel metal2 s 111982 0 112038 800 6 t1x[31]
port 325 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 t1x[3]
port 326 nsew signal input
rlabel metal2 s 52366 0 52422 800 6 t1x[4]
port 327 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 t1x[5]
port 328 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 t1x[6]
port 329 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 t1x[7]
port 330 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 t1x[8]
port 331 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 t1x[9]
port 332 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 t1y[0]
port 333 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 t1y[10]
port 334 nsew signal input
rlabel metal2 s 68190 0 68246 800 6 t1y[11]
port 335 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 t1y[12]
port 336 nsew signal input
rlabel metal2 s 72606 0 72662 800 6 t1y[13]
port 337 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 t1y[14]
port 338 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 t1y[15]
port 339 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 t1y[16]
port 340 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 t1y[17]
port 341 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 t1y[18]
port 342 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 t1y[19]
port 343 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 t1y[1]
port 344 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 t1y[20]
port 345 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 t1y[21]
port 346 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 t1y[22]
port 347 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 t1y[23]
port 348 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 t1y[24]
port 349 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 t1y[25]
port 350 nsew signal input
rlabel metal2 s 101310 0 101366 800 6 t1y[26]
port 351 nsew signal input
rlabel metal2 s 103518 0 103574 800 6 t1y[27]
port 352 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 t1y[28]
port 353 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 t1y[29]
port 354 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 t1y[2]
port 355 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 t1y[30]
port 356 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 t1y[31]
port 357 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 t1y[3]
port 358 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 t1y[4]
port 359 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 t1y[5]
port 360 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 t1y[6]
port 361 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 t1y[7]
port 362 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 t1y[8]
port 363 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 t1y[9]
port 364 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 t2x[0]
port 365 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 t2x[10]
port 366 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 t2x[11]
port 367 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 t2x[12]
port 368 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 t2x[13]
port 369 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 t2x[14]
port 370 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 t2x[15]
port 371 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 t2x[16]
port 372 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 t2x[17]
port 373 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 t2x[18]
port 374 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 t2x[19]
port 375 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 t2x[1]
port 376 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 t2x[20]
port 377 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 t2x[21]
port 378 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 t2x[22]
port 379 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 t2x[23]
port 380 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 t2x[24]
port 381 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 t2x[25]
port 382 nsew signal input
rlabel metal2 s 101678 0 101734 800 6 t2x[26]
port 383 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 t2x[27]
port 384 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 t2x[28]
port 385 nsew signal input
rlabel metal2 s 108302 0 108358 800 6 t2x[29]
port 386 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 t2x[2]
port 387 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 t2x[30]
port 388 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 t2x[31]
port 389 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 t2x[3]
port 390 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 t2x[4]
port 391 nsew signal input
rlabel metal2 s 55310 0 55366 800 6 t2x[5]
port 392 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 t2x[6]
port 393 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 t2x[7]
port 394 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 t2x[8]
port 395 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 t2x[9]
port 396 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 t2y[0]
port 397 nsew signal input
rlabel metal2 s 66718 0 66774 800 6 t2y[10]
port 398 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 t2y[11]
port 399 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 t2y[12]
port 400 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 t2y[13]
port 401 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 t2y[14]
port 402 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 t2y[15]
port 403 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 t2y[16]
port 404 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 t2y[17]
port 405 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 t2y[18]
port 406 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 t2y[19]
port 407 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 t2y[1]
port 408 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 t2y[20]
port 409 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 t2y[21]
port 410 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 t2y[22]
port 411 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 t2y[23]
port 412 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 t2y[24]
port 413 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 t2y[25]
port 414 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 t2y[26]
port 415 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 t2y[27]
port 416 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 t2y[28]
port 417 nsew signal input
rlabel metal2 s 108670 0 108726 800 6 t2y[29]
port 418 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 t2y[2]
port 419 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 t2y[30]
port 420 nsew signal input
rlabel metal2 s 113086 0 113142 800 6 t2y[31]
port 421 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 t2y[3]
port 422 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 t2y[4]
port 423 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 t2y[5]
port 424 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 t2y[6]
port 425 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 t2y[7]
port 426 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 t2y[8]
port 427 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 t2y[9]
port 428 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 v0z[0]
port 429 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 v0z[10]
port 430 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 v0z[11]
port 431 nsew signal input
rlabel metal2 s 20718 0 20774 800 6 v0z[12]
port 432 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 v0z[13]
port 433 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 v0z[14]
port 434 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 v0z[15]
port 435 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 v0z[16]
port 436 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 v0z[17]
port 437 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 v0z[18]
port 438 nsew signal input
rlabel metal2 s 28446 0 28502 800 6 v0z[19]
port 439 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 v0z[1]
port 440 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 v0z[20]
port 441 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 v0z[21]
port 442 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 v0z[22]
port 443 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 v0z[23]
port 444 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 v0z[24]
port 445 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 v0z[25]
port 446 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 v0z[26]
port 447 nsew signal input
rlabel metal2 s 37278 0 37334 800 6 v0z[27]
port 448 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 v0z[28]
port 449 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 v0z[29]
port 450 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 v0z[2]
port 451 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 v0z[30]
port 452 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 v0z[31]
port 453 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 v0z[3]
port 454 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 v0z[4]
port 455 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 v0z[5]
port 456 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 v0z[6]
port 457 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 v0z[7]
port 458 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 v0z[8]
port 459 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 v0z[9]
port 460 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 v1z[0]
port 461 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 v1z[10]
port 462 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 v1z[11]
port 463 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 v1z[12]
port 464 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 v1z[13]
port 465 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 v1z[14]
port 466 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 v1z[15]
port 467 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 v1z[16]
port 468 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 v1z[17]
port 469 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 v1z[18]
port 470 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 v1z[19]
port 471 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 v1z[1]
port 472 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 v1z[20]
port 473 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 v1z[21]
port 474 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 v1z[22]
port 475 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 v1z[23]
port 476 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 v1z[24]
port 477 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 v1z[25]
port 478 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 v1z[26]
port 479 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 v1z[27]
port 480 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 v1z[28]
port 481 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 v1z[29]
port 482 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 v1z[2]
port 483 nsew signal input
rlabel metal2 s 40958 0 41014 800 6 v1z[30]
port 484 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 v1z[31]
port 485 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 v1z[3]
port 486 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 v1z[4]
port 487 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 v1z[5]
port 488 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 v1z[6]
port 489 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 v1z[7]
port 490 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 v1z[8]
port 491 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 v1z[9]
port 492 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 v2z[0]
port 493 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 v2z[10]
port 494 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 v2z[11]
port 495 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 v2z[12]
port 496 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 v2z[13]
port 497 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 v2z[14]
port 498 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 v2z[15]
port 499 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 v2z[16]
port 500 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 v2z[17]
port 501 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 v2z[18]
port 502 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 v2z[19]
port 503 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 v2z[1]
port 504 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 v2z[20]
port 505 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 v2z[21]
port 506 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 v2z[22]
port 507 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 v2z[23]
port 508 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 v2z[24]
port 509 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 v2z[25]
port 510 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 v2z[26]
port 511 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 v2z[27]
port 512 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 v2z[28]
port 513 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 v2z[29]
port 514 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 v2z[2]
port 515 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 v2z[30]
port 516 nsew signal input
rlabel metal2 s 42430 0 42486 800 6 v2z[31]
port 517 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 v2z[3]
port 518 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 v2z[4]
port 519 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 v2z[5]
port 520 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 v2z[6]
port 521 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 v2z[7]
port 522 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 v2z[8]
port 523 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 v2z[9]
port 524 nsew signal input
rlabel metal4 s 4208 2128 4528 87632 6 vccd1
port 525 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 87632 6 vccd1
port 525 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 87632 6 vccd1
port 525 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 87632 6 vccd1
port 525 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 87632 6 vssd1
port 526 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 87632 6 vssd1
port 526 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 87632 6 vssd1
port 526 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 87632 6 vssd1
port 526 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 120000 90000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 40696618
string GDS_FILE /local/colinm22/sdmay26-24/openlane/wavg_pipe/runs/25_10_19_13_59/results/signoff/wavg_pipe_m.magic.gds
string GDS_START 1378202
<< end >>

