* NGSPICE file created from wavg_pipe_m.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_2 abstract view
.subckt sky130_fd_sc_hd__a32oi_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_1 abstract view
.subckt sky130_fd_sc_hd__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

.subckt wavg_pipe_m clk_i mstream_i mstream_o[0] mstream_o[100] mstream_o[101] mstream_o[102]
+ mstream_o[103] mstream_o[104] mstream_o[105] mstream_o[106] mstream_o[107] mstream_o[108]
+ mstream_o[109] mstream_o[10] mstream_o[110] mstream_o[111] mstream_o[112] mstream_o[113]
+ mstream_o[114] mstream_o[115] mstream_o[11] mstream_o[12] mstream_o[13] mstream_o[14]
+ mstream_o[15] mstream_o[16] mstream_o[17] mstream_o[18] mstream_o[19] mstream_o[1]
+ mstream_o[20] mstream_o[21] mstream_o[22] mstream_o[23] mstream_o[24] mstream_o[25]
+ mstream_o[26] mstream_o[27] mstream_o[28] mstream_o[29] mstream_o[2] mstream_o[30]
+ mstream_o[31] mstream_o[32] mstream_o[33] mstream_o[34] mstream_o[35] mstream_o[36]
+ mstream_o[37] mstream_o[38] mstream_o[39] mstream_o[3] mstream_o[40] mstream_o[41]
+ mstream_o[42] mstream_o[43] mstream_o[44] mstream_o[45] mstream_o[46] mstream_o[47]
+ mstream_o[48] mstream_o[49] mstream_o[4] mstream_o[50] mstream_o[51] mstream_o[52]
+ mstream_o[53] mstream_o[54] mstream_o[55] mstream_o[56] mstream_o[57] mstream_o[58]
+ mstream_o[59] mstream_o[5] mstream_o[60] mstream_o[61] mstream_o[62] mstream_o[63]
+ mstream_o[64] mstream_o[65] mstream_o[66] mstream_o[67] mstream_o[68] mstream_o[69]
+ mstream_o[6] mstream_o[70] mstream_o[71] mstream_o[72] mstream_o[73] mstream_o[74]
+ mstream_o[75] mstream_o[76] mstream_o[77] mstream_o[78] mstream_o[79] mstream_o[7]
+ mstream_o[80] mstream_o[81] mstream_o[82] mstream_o[83] mstream_o[84] mstream_o[85]
+ mstream_o[86] mstream_o[87] mstream_o[88] mstream_o[89] mstream_o[8] mstream_o[90]
+ mstream_o[91] mstream_o[92] mstream_o[93] mstream_o[94] mstream_o[95] mstream_o[96]
+ mstream_o[97] mstream_o[98] mstream_o[99] mstream_o[9] nrst_i sstream_i[0] sstream_i[100]
+ sstream_i[101] sstream_i[102] sstream_i[103] sstream_i[104] sstream_i[105] sstream_i[106]
+ sstream_i[107] sstream_i[108] sstream_i[109] sstream_i[10] sstream_i[110] sstream_i[111]
+ sstream_i[112] sstream_i[113] sstream_i[114] sstream_i[115] sstream_i[11] sstream_i[12]
+ sstream_i[13] sstream_i[14] sstream_i[15] sstream_i[16] sstream_i[17] sstream_i[18]
+ sstream_i[19] sstream_i[1] sstream_i[20] sstream_i[21] sstream_i[22] sstream_i[23]
+ sstream_i[24] sstream_i[25] sstream_i[26] sstream_i[27] sstream_i[28] sstream_i[29]
+ sstream_i[2] sstream_i[30] sstream_i[31] sstream_i[32] sstream_i[33] sstream_i[34]
+ sstream_i[35] sstream_i[36] sstream_i[37] sstream_i[38] sstream_i[39] sstream_i[3]
+ sstream_i[40] sstream_i[41] sstream_i[42] sstream_i[43] sstream_i[44] sstream_i[45]
+ sstream_i[46] sstream_i[47] sstream_i[48] sstream_i[49] sstream_i[4] sstream_i[50]
+ sstream_i[51] sstream_i[52] sstream_i[53] sstream_i[54] sstream_i[55] sstream_i[56]
+ sstream_i[57] sstream_i[58] sstream_i[59] sstream_i[5] sstream_i[60] sstream_i[61]
+ sstream_i[62] sstream_i[63] sstream_i[64] sstream_i[65] sstream_i[66] sstream_i[67]
+ sstream_i[68] sstream_i[69] sstream_i[6] sstream_i[70] sstream_i[71] sstream_i[72]
+ sstream_i[73] sstream_i[74] sstream_i[75] sstream_i[76] sstream_i[77] sstream_i[78]
+ sstream_i[79] sstream_i[7] sstream_i[80] sstream_i[81] sstream_i[82] sstream_i[83]
+ sstream_i[84] sstream_i[85] sstream_i[86] sstream_i[87] sstream_i[88] sstream_i[89]
+ sstream_i[8] sstream_i[90] sstream_i[91] sstream_i[92] sstream_i[93] sstream_i[94]
+ sstream_i[95] sstream_i[96] sstream_i[97] sstream_i[98] sstream_i[99] sstream_i[9]
+ sstream_o t0x[0] t0x[10] t0x[11] t0x[12] t0x[13] t0x[14] t0x[15] t0x[16] t0x[17]
+ t0x[18] t0x[19] t0x[1] t0x[20] t0x[21] t0x[22] t0x[23] t0x[24] t0x[25] t0x[26] t0x[27]
+ t0x[28] t0x[29] t0x[2] t0x[30] t0x[31] t0x[3] t0x[4] t0x[5] t0x[6] t0x[7] t0x[8]
+ t0x[9] t0y[0] t0y[10] t0y[11] t0y[12] t0y[13] t0y[14] t0y[15] t0y[16] t0y[17] t0y[18]
+ t0y[19] t0y[1] t0y[20] t0y[21] t0y[22] t0y[23] t0y[24] t0y[25] t0y[26] t0y[27] t0y[28]
+ t0y[29] t0y[2] t0y[30] t0y[31] t0y[3] t0y[4] t0y[5] t0y[6] t0y[7] t0y[8] t0y[9]
+ t1x[0] t1x[10] t1x[11] t1x[12] t1x[13] t1x[14] t1x[15] t1x[16] t1x[17] t1x[18] t1x[19]
+ t1x[1] t1x[20] t1x[21] t1x[22] t1x[23] t1x[24] t1x[25] t1x[26] t1x[27] t1x[28] t1x[29]
+ t1x[2] t1x[30] t1x[31] t1x[3] t1x[4] t1x[5] t1x[6] t1x[7] t1x[8] t1x[9] t1y[0] t1y[10]
+ t1y[11] t1y[12] t1y[13] t1y[14] t1y[15] t1y[16] t1y[17] t1y[18] t1y[19] t1y[1] t1y[20]
+ t1y[21] t1y[22] t1y[23] t1y[24] t1y[25] t1y[26] t1y[27] t1y[28] t1y[29] t1y[2] t1y[30]
+ t1y[31] t1y[3] t1y[4] t1y[5] t1y[6] t1y[7] t1y[8] t1y[9] t2x[0] t2x[10] t2x[11]
+ t2x[12] t2x[13] t2x[14] t2x[15] t2x[16] t2x[17] t2x[18] t2x[19] t2x[1] t2x[20] t2x[21]
+ t2x[22] t2x[23] t2x[24] t2x[25] t2x[26] t2x[27] t2x[28] t2x[29] t2x[2] t2x[30] t2x[31]
+ t2x[3] t2x[4] t2x[5] t2x[6] t2x[7] t2x[8] t2x[9] t2y[0] t2y[10] t2y[11] t2y[12]
+ t2y[13] t2y[14] t2y[15] t2y[16] t2y[17] t2y[18] t2y[19] t2y[1] t2y[20] t2y[21] t2y[22]
+ t2y[23] t2y[24] t2y[25] t2y[26] t2y[27] t2y[28] t2y[29] t2y[2] t2y[30] t2y[31] t2y[3]
+ t2y[4] t2y[5] t2y[6] t2y[7] t2y[8] t2y[9] v0z[0] v0z[10] v0z[11] v0z[12] v0z[13]
+ v0z[14] v0z[15] v0z[16] v0z[17] v0z[18] v0z[19] v0z[1] v0z[20] v0z[21] v0z[22] v0z[23]
+ v0z[24] v0z[25] v0z[26] v0z[27] v0z[28] v0z[29] v0z[2] v0z[30] v0z[31] v0z[3] v0z[4]
+ v0z[5] v0z[6] v0z[7] v0z[8] v0z[9] v1z[0] v1z[10] v1z[11] v1z[12] v1z[13] v1z[14]
+ v1z[15] v1z[16] v1z[17] v1z[18] v1z[19] v1z[1] v1z[20] v1z[21] v1z[22] v1z[23] v1z[24]
+ v1z[25] v1z[26] v1z[27] v1z[28] v1z[29] v1z[2] v1z[30] v1z[31] v1z[3] v1z[4] v1z[5]
+ v1z[6] v1z[7] v1z[8] v1z[9] v2z[0] v2z[10] v2z[11] v2z[12] v2z[13] v2z[14] v2z[15]
+ v2z[16] v2z[17] v2z[18] v2z[19] v2z[1] v2z[20] v2z[21] v2z[22] v2z[23] v2z[24] v2z[25]
+ v2z[26] v2z[27] v2z[28] v2z[29] v2z[2] v2z[30] v2z[31] v2z[3] v2z[4] v2z[5] v2z[6]
+ v2z[7] v2z[8] v2z[9] vccd1 vssd1
XFILLER_0_118_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18869_ _18733_/A _18735_/B _18733_/B vssd1 vssd1 vccd1 vccd1 _18874_/A sky130_fd_sc_hd__o21bai_1
XANTENNA__17597__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20900_ _20900_/A _20900_/B vssd1 vssd1 vccd1 vccd1 _20902_/B sky130_fd_sc_hd__nand2_1
X_21880_ _21945_/CLK _21880_/D vssd1 vssd1 vccd1 vccd1 hold208/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20831_ _20830_/B _20830_/C _20830_/A vssd1 vssd1 vccd1 vccd1 _20831_/X sky130_fd_sc_hd__o21a_1
XANTENNA_fanout162_A _17324_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18546__A1 _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20762_ _20759_/Y _20760_/X _20630_/Y _20632_/Y vssd1 vssd1 vccd1 vccd1 _20762_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20693_ _20694_/A _20694_/B vssd1 vssd1 vccd1 vccd1 _20823_/A sky130_fd_sc_hd__or2_1
XFILLER_0_18_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout427_A _21763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_780 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20105__A1 _21832_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20105__B2 _21831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17757__A _18008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17521__A2 _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21314_ hold294/A _21168_/A _21171_/D _21056_/B _21171_/A vssd1 vssd1 vccd1 vccd1
+ _21316_/A sky130_fd_sc_hd__o2111a_1
XFILLER_0_130_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16380__B _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11149__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21245_ _21244_/A _21244_/B _21244_/C vssd1 vssd1 vccd1 vccd1 _21246_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_41_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19972__A _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14181__A _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20333__D _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21176_ _21176_/A _21176_/B vssd1 vssd1 vccd1 vccd1 _21178_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_99_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20127_ _20863_/C _21278_/A _20265_/D _21199_/A vssd1 vssd1 vccd1 vccd1 _20130_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout75_A _21848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20058_ _20203_/B _20056_/Y _19830_/X _19832_/Y vssd1 vssd1 vccd1 vccd1 _20059_/C
+ sky130_fd_sc_hd__a211oi_1
XTAP_3202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15048__B1 _15046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13525__A _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18785__B2 _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11900_ _11900_/A _11900_/B vssd1 vssd1 vccd1 vccd1 _11901_/C sky130_fd_sc_hd__nor2_1
XTAP_3235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ _12880_/A _12880_/B vssd1 vssd1 vccd1 vccd1 _12889_/A sky130_fd_sc_hd__xor2_1
XANTENNA__16796__B1 _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20592__B2 _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_202 hold268/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_213 hold275/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _11801_/A _11801_/B _11801_/C vssd1 vssd1 vccd1 vccd1 _11831_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA_224 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_235 hold299/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_246 _11347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_257 hold262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_268 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14550_ _14690_/B _14548_/C _14548_/A vssd1 vssd1 vccd1 vccd1 _14551_/C sky130_fd_sc_hd__a21o_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11762_ _11761_/A _11761_/C _11761_/B vssd1 vssd1 vccd1 vccd1 _11764_/B sky130_fd_sc_hd__a21o_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_279 hold283/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16555__B _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13501_ _13523_/B _13501_/B _13500_/C _13500_/D vssd1 vssd1 vccd1 vccd1 _13501_/X
+ sky130_fd_sc_hd__or4bb_2
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14481_ _14480_/B _14632_/B _14480_/A vssd1 vssd1 vccd1 vccd1 _14482_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_67_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14356__A _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13898__C _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11693_ _12750_/A _12020_/A _12326_/D _12528_/B vssd1 vssd1 vccd1 vccd1 _11694_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16220_ _16221_/B _16221_/A vssd1 vssd1 vccd1 vccd1 _16337_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__13260__A _13554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13432_ _13280_/A _13280_/Y _13430_/X _13431_/Y vssd1 vssd1 vccd1 vccd1 _13496_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19866__B _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14075__B _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11388__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16151_ _16151_/A _16151_/B vssd1 vssd1 vccd1 vccd1 _16152_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20647__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13363_ _13363_/A _13363_/B vssd1 vssd1 vccd1 vccd1 _13518_/C sky130_fd_sc_hd__nand2_4
XFILLER_0_23_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15102_ _15226_/A _15101_/C _15101_/A vssd1 vssd1 vccd1 vccd1 _15103_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_122_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12314_ _12315_/A _12315_/B vssd1 vssd1 vccd1 vccd1 _12314_/X sky130_fd_sc_hd__and2b_1
X_16082_ _16079_/X _16080_/Y _15909_/B _15948_/Y vssd1 vssd1 vccd1 vccd1 _16128_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13294_ _14365_/A _14367_/A _15514_/A _15514_/B vssd1 vssd1 vccd1 vccd1 _13445_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_146_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15033_ _15933_/C _16409_/A _15034_/C _15127_/A vssd1 vssd1 vccd1 vccd1 _15035_/B
+ sky130_fd_sc_hd__a22o_1
X_19910_ _19909_/B _20001_/B _19909_/A vssd1 vssd1 vccd1 vccd1 _19911_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_32_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12245_ _12269_/A _12245_/B _12246_/C _12246_/D vssd1 vssd1 vccd1 vccd1 _12245_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_82_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17276__B2 _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ _12168_/A _12168_/C _12168_/B vssd1 vssd1 vccd1 vccd1 _12176_/Y sky130_fd_sc_hd__o21ai_1
X_19841_ _19841_/A _19841_/B vssd1 vssd1 vccd1 vccd1 _19843_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1087 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11127_ hold225/X _11126_/A _11126_/B hold200/X vssd1 vssd1 vccd1 vccd1 _11127_/X
+ sky130_fd_sc_hd__a22o_1
X_16984_ _16984_/A _16984_/B vssd1 vssd1 vccd1 vccd1 _16986_/B sky130_fd_sc_hd__xnor2_1
X_19772_ _19772_/A _19772_/B vssd1 vssd1 vccd1 vccd1 _19773_/B sky130_fd_sc_hd__xor2_2
XANTENNA__20813__A1_N _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15935_ _15936_/B _15936_/A vssd1 vssd1 vccd1 vccd1 _16069_/A sky130_fd_sc_hd__nand2b_1
X_11058_ _11057_/Y hold42/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21658_/D sky130_fd_sc_hd__mux2_1
X_18723_ _18563_/Y _18566_/X _18721_/Y _18722_/X vssd1 vssd1 vccd1 vccd1 _18847_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18010__B _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17552__D _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18654_ _18653_/B _18653_/C _18653_/A vssd1 vssd1 vccd1 vccd1 _18656_/B sky130_fd_sc_hd__a21o_1
X_15866_ _15863_/Y _15864_/X _15726_/X _15728_/X vssd1 vssd1 vccd1 vccd1 _15867_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_14_clk_i_A _21806_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14817_ _16374_/A _16196_/A _14817_/C _14817_/D vssd1 vssd1 vccd1 vccd1 _14820_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_99_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17605_ _17605_/A vssd1 vssd1 vccd1 vccd1 _17607_/A sky130_fd_sc_hd__inv_2
X_18585_ _19644_/A _19382_/B _18583_/Y _18584_/X vssd1 vssd1 vccd1 vccd1 _18587_/A
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15797_ _15798_/A _15798_/B vssd1 vssd1 vccd1 vccd1 _15986_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_118_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17536_ _17536_/A _17536_/B _17536_/C vssd1 vssd1 vccd1 vccd1 _17536_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__21532__A0 hold262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14748_ _14588_/A _14588_/B _14586_/Y vssd1 vssd1 vccd1 vccd1 _14750_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_47_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12993__B _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17467_ _17466_/A _17466_/B _17466_/C _17466_/D vssd1 vssd1 vccd1 vccd1 _17467_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_156_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10794__A _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14679_ _14679_/A _14679_/B _14679_/C vssd1 vssd1 vccd1 vccd1 _14682_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15211__B1 _10926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18961__A _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16418_ _16418_/A _16418_/B vssd1 vssd1 vccd1 vccd1 _16420_/A sky130_fd_sc_hd__nand2_1
X_19206_ _19195_/Y _19206_/B _19206_/C vssd1 vssd1 vccd1 vccd1 _19363_/A sky130_fd_sc_hd__and3b_1
X_17398_ _17398_/A _17398_/B vssd1 vssd1 vccd1 vccd1 _17400_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11379__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19137_ _18975_/B _18975_/Y _19135_/X _19136_/Y vssd1 vssd1 vccd1 vccd1 _19139_/B
+ sky130_fd_sc_hd__a211o_2
X_16349_ _16349_/A _16349_/B _16349_/C vssd1 vssd1 vccd1 vccd1 _16368_/B sky130_fd_sc_hd__or3_1
XFILLER_0_15_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13320__D _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17503__A2 _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18700__A1 _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18700__B2 _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21099__A _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19068_ _19692_/A _19535_/B _19068_/C _19238_/C vssd1 vssd1 vccd1 vccd1 _19235_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_113_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14713__B _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18019_ _18018_/A _18018_/B _18018_/C vssd1 vssd1 vccd1 vccd1 _18020_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_112_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19256__A2 _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21030_ hold100/X _21029_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _21914_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_2_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout105 _19691_/D vssd1 vssd1 vccd1 vccd1 _20416_/B sky130_fd_sc_hd__buf_4
XFILLER_0_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout116 _21839_/Q vssd1 vssd1 vccd1 vccd1 _20148_/C sky130_fd_sc_hd__buf_6
Xfanout127 _20910_/A vssd1 vssd1 vccd1 vccd1 _17636_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__20810__A2 _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout138 _18929_/B vssd1 vssd1 vccd1 vccd1 _18767_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout149 _21832_/Q vssd1 vssd1 vccd1 vccd1 _19092_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__18201__A _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16490__A2 _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout377_A _14828_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21932_ _21932_/CLK _21932_/D vssd1 vssd1 vccd1 vccd1 hold191/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21863_ _21932_/CLK _21863_/D vssd1 vssd1 vccd1 vccd1 hold315/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout544_A _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19032__A _19650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21523__A0 hold290/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20814_ _20938_/A _21278_/B _21171_/A _20814_/D vssd1 vssd1 vccd1 vccd1 _20938_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_38_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21794_ _22016_/CLK _21794_/D vssd1 vssd1 vccd1 vccd1 _21794_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_92_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19967__A _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20745_ _20615_/X _20617_/X _20743_/Y _20744_/X vssd1 vssd1 vccd1 vccd1 _20747_/B
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__14176__A _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17742__A2 _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20676_ _21256_/A _21040_/A _20677_/C _20677_/D vssd1 vssd1 vccd1 vccd1 _20678_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__19686__B _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14326__D _14635_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16391__A _16391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15719__B _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16541__D _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17724__A2_N _19053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12030_ _12286_/B _12030_/B vssd1 vssd1 vccd1 vccd1 _12036_/C sky130_fd_sc_hd__or2_1
X_21228_ _21228_/A _21228_/B _21228_/C vssd1 vssd1 vccd1 vccd1 _21229_/B sky130_fd_sc_hd__nor3_1
Xhold170 hold170/A vssd1 vssd1 vccd1 vccd1 hold170/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 hold181/A vssd1 vssd1 vccd1 vccd1 hold181/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12143__B _12242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold192 hold192/A vssd1 vssd1 vccd1 vccd1 hold192/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19852__D _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21159_ _21159_/A _21159_/B vssd1 vssd1 vccd1 vccd1 _21159_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__18749__C _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15454__B _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16481__A2 _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13981_ _13981_/A _13981_/B vssd1 vssd1 vccd1 vccd1 _13989_/A sky130_fd_sc_hd__xnor2_1
X_15720_ _15720_/A _15848_/B vssd1 vssd1 vccd1 vccd1 _15722_/B sky130_fd_sc_hd__or2_1
XTAP_3010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12932_ _12803_/C _12802_/Y _12929_/X _12930_/Y vssd1 vssd1 vccd1 vccd1 _12934_/C
+ sky130_fd_sc_hd__o211ai_4
XTAP_3021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15651_ _15561_/A _15561_/C _15561_/B vssd1 vssd1 vccd1 vccd1 _15687_/A sky130_fd_sc_hd__a21boi_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ _12989_/B _12862_/C _12862_/A vssd1 vssd1 vccd1 vccd1 _12864_/B sky130_fd_sc_hd__a21o_1
XTAP_3076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15441__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14602_ _14603_/B _14603_/C _14911_/A vssd1 vssd1 vccd1 vccd1 _14608_/B sky130_fd_sc_hd__o21a_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18370_ _18220_/C _18219_/Y _18368_/X _18369_/Y vssd1 vssd1 vccd1 vccd1 _18373_/C
+ sky130_fd_sc_hd__o211a_2
XANTENNA__18484__C _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11814_ _11813_/A _11813_/C _11813_/B vssd1 vssd1 vccd1 vccd1 _11816_/B sky130_fd_sc_hd__a21o_1
X_15582_ _15582_/A _15582_/B vssd1 vssd1 vccd1 vccd1 _15585_/A sky130_fd_sc_hd__xnor2_2
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20088__A _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12794_ _12681_/A _12681_/C _12681_/B vssd1 vssd1 vccd1 vccd1 _12795_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_150_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17321_ _17223_/A _20088_/A _17226_/B _17224_/X vssd1 vssd1 vccd1 vccd1 _17331_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14533_ _14412_/A _14411_/B _14409_/X vssd1 vssd1 vccd1 vccd1 _14548_/A sky130_fd_sc_hd__a21o_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ _11744_/A _11744_/C _11744_/B vssd1 vssd1 vccd1 vccd1 _11748_/B sky130_fd_sc_hd__a21o_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18930__A1 _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17252_ _17251_/B _17251_/C _17251_/A vssd1 vssd1 vccd1 vccd1 _17252_/Y sky130_fd_sc_hd__a21oi_2
X_14464_ _14466_/A vssd1 vssd1 vccd1 vccd1 _14629_/A sky130_fd_sc_hd__inv_2
XFILLER_0_138_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11676_ _11673_/X _11676_/B vssd1 vssd1 vccd1 vccd1 _11763_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16203_ _15695_/A _16406_/B _16314_/D _16203_/D vssd1 vssd1 vccd1 vccd1 _16321_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_126_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13415_ _13415_/A _13415_/B vssd1 vssd1 vccd1 vccd1 _13415_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17183_ _17277_/A _17741_/B _17183_/C _17183_/D vssd1 vssd1 vccd1 vccd1 _17186_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_4_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14395_ _14395_/A _14532_/A _14395_/C vssd1 vssd1 vccd1 vccd1 _14532_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_10_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19486__A2 _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12037__C _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16134_ _16134_/A _16134_/B _16134_/C vssd1 vssd1 vccd1 vccd1 _16134_/X sky130_fd_sc_hd__and3_1
XFILLER_0_141_539 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11230__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_271 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13346_ _13343_/X _13344_/Y _13204_/B _13203_/Y vssd1 vssd1 vccd1 vccd1 _13348_/C
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__11230__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18694__B1 _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16065_ _16064_/B _16064_/C _16064_/A vssd1 vssd1 vccd1 vccd1 _16066_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_122_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16451__D _16743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13277_ _13136_/A _13136_/C _13136_/B vssd1 vssd1 vccd1 vccd1 _13278_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_110_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15016_ _16087_/A _16092_/D _15653_/C _15112_/D vssd1 vssd1 vccd1 vccd1 _15017_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__21045__A2 _21816_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12228_ _12228_/A _12228_/B _12228_/C vssd1 vssd1 vccd1 vccd1 _12234_/A sky130_fd_sc_hd__and3_1
XANTENNA__15645__A _15645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19824_ _20462_/D _20193_/D _19825_/C _20043_/A vssd1 vssd1 vccd1 vccd1 _19826_/B
+ sky130_fd_sc_hd__a22o_1
X_12159_ _12160_/A _12160_/B _12160_/C vssd1 vssd1 vccd1 vccd1 _12159_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_75_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20270__B _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19755_ _19752_/X _19753_/Y _19572_/Y _19574_/X vssd1 vssd1 vccd1 vccd1 _19756_/C
+ sky130_fd_sc_hd__a211o_1
X_16967_ _16920_/A _16920_/C _16920_/B vssd1 vssd1 vccd1 vccd1 _16973_/B sky130_fd_sc_hd__a21o_1
XANTENNA__17860__A _19337_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11297__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18706_ _18707_/A _18707_/B vssd1 vssd1 vccd1 vccd1 _18708_/A sky130_fd_sc_hd__and2_1
X_15918_ _16369_/A _16396_/A _15919_/C _15919_/D vssd1 vssd1 vccd1 vccd1 _15920_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__12494__B1 _11048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16898_ _16898_/A _16898_/B vssd1 vssd1 vccd1 vccd1 _16951_/A sky130_fd_sc_hd__nor2_1
X_19686_ _19686_/A _19686_/B _20265_/D vssd1 vssd1 vccd1 vccd1 _19686_/X sky130_fd_sc_hd__and3_1
XFILLER_0_91_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17421__A1 _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15849_ _15849_/A _15849_/B vssd1 vssd1 vccd1 vccd1 _15857_/A sky130_fd_sc_hd__nand2_1
X_18637_ _18787_/B _19092_/C _19262_/C _18787_/A vssd1 vssd1 vccd1 vccd1 _18640_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14235__A1 _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17972__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20308__A1 _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14786__A2 _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20308__B2 _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18568_ _18413_/Y _18416_/X _18565_/Y _18567_/X vssd1 vssd1 vccd1 vccd1 _18572_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_75_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1076 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20859__A2 _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17519_ _17602_/A _17517_/Y _17405_/B _17405_/Y vssd1 vssd1 vccd1 vccd1 _17580_/B
+ sky130_fd_sc_hd__a211o_1
X_18499_ _19123_/B _19872_/C _19972_/C _19123_/A vssd1 vssd1 vccd1 vccd1 _18500_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20530_ _20913_/A _20531_/B vssd1 vssd1 vccd1 vccd1 _20530_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__20148__D _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20461_ _20461_/A _20461_/B vssd1 vssd1 vccd1 vccd1 _20465_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout125_A _20689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20392_ _20249_/A _20249_/B _20250_/A _20248_/B vssd1 vssd1 vccd1 vccd1 _20398_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13761__A3 _14218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22062_ _22063_/CLK _22062_/D vssd1 vssd1 vccd1 vccd1 hold277/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__21036__A2 _21283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout494_A _21745_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21013_ _21012_/B _21012_/C _21012_/A vssd1 vssd1 vccd1 vccd1 _21014_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_10_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17660__A1 _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15274__B _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15671__B1 _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17412__A1 _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21915_ _21949_/CLK hold147/X vssd1 vssd1 vccd1 vccd1 hold146/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__17412__B2 _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15423__B1 _15243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21846_ _21853_/CLK _21846_/D vssd1 vssd1 vccd1 vccd1 _21846_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21777_ _21809_/CLK _21777_/D vssd1 vssd1 vccd1 vccd1 _21777_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_65_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11530_ _11529_/X _19201_/B _11545_/S vssd1 vssd1 vccd1 vccd1 _21848_/D sky130_fd_sc_hd__mux2_1
XANTENNA__11460__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20728_ _20728_/A _20728_/B vssd1 vssd1 vccd1 vccd1 _20747_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout4_A fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11461_ _11460_/X _17666_/A _11470_/S vssd1 vssd1 vccd1 vccd1 _21825_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_34_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20659_ _20913_/A _20660_/B vssd1 vssd1 vccd1 vccd1 _20659_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_80_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13200_ _13199_/B _13199_/C _13199_/A vssd1 vssd1 vccd1 vccd1 _13200_/Y sky130_fd_sc_hd__a21oi_2
X_14180_ _14508_/A _14817_/C _14817_/D _14813_/A vssd1 vssd1 vccd1 vccd1 _14185_/C
+ sky130_fd_sc_hd__a22o_1
X_11392_ _11391_/X _17433_/A _11401_/S vssd1 vssd1 vccd1 vccd1 _21802_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14353__B _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13131_ _13867_/A _13269_/C _13269_/D _13858_/A vssd1 vssd1 vccd1 vccd1 _13132_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13062_ _13062_/A _13062_/B _13062_/C vssd1 vssd1 vccd1 vccd1 _13062_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__12712__A1 _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11993__A _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ _12011_/A _12011_/Y _12012_/Y _11941_/X vssd1 vssd1 vccd1 vccd1 _12029_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12712__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17870_ _17870_/A _17870_/B vssd1 vssd1 vccd1 vccd1 _17878_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16821_ _16822_/A _16822_/B vssd1 vssd1 vccd1 vccd1 _16840_/B sky130_fd_sc_hd__nand2b_1
Xfanout480 _14217_/D vssd1 vssd1 vccd1 vccd1 _16040_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14465__B2 _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12601__B _21340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout491 _21746_/Q vssd1 vssd1 vccd1 vccd1 _14212_/D sky130_fd_sc_hd__buf_4
X_16752_ _16753_/A _16753_/B vssd1 vssd1 vccd1 vccd1 _16773_/B sky130_fd_sc_hd__nand2_1
X_19540_ _19536_/X _19538_/Y _19378_/X _19381_/X vssd1 vssd1 vccd1 vccd1 _19541_/B
+ sky130_fd_sc_hd__a211o_1
X_13964_ _13814_/B _13964_/B vssd1 vssd1 vccd1 vccd1 _14294_/B sky130_fd_sc_hd__and2b_1
X_15703_ _15705_/A vssd1 vssd1 vccd1 vccd1 _15846_/A sky130_fd_sc_hd__inv_2
X_12915_ _12787_/A _12787_/C _12787_/B vssd1 vssd1 vccd1 vccd1 _12916_/C sky130_fd_sc_hd__a21bo_1
X_16683_ _16682_/A _16681_/Y _16657_/X _16658_/Y vssd1 vssd1 vccd1 vccd1 _16686_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__18746__A4 _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19471_ _19472_/A _19472_/B vssd1 vssd1 vccd1 vccd1 _19471_/X sky130_fd_sc_hd__or2_1
X_13895_ _14367_/A _14537_/A vssd1 vssd1 vccd1 vccd1 _13896_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_115_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15634_ _16027_/A _16369_/B _15635_/C _15635_/D vssd1 vssd1 vccd1 vccd1 _15640_/A
+ sky130_fd_sc_hd__a22oi_1
X_18422_ _18307_/X _18310_/Y _18543_/B _18421_/X vssd1 vssd1 vccd1 vccd1 _18542_/A
+ sky130_fd_sc_hd__a211oi_2
X_12846_ _14138_/A _13258_/C _13258_/D _13975_/B vssd1 vssd1 vccd1 vccd1 _12848_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12779__A1 _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12779__B2 _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18353_ _18352_/B _18352_/C _18352_/A vssd1 vssd1 vccd1 vccd1 _18355_/B sky130_fd_sc_hd__a21o_1
X_15565_ _15420_/B _15420_/Y _15563_/Y _15564_/X vssd1 vssd1 vccd1 vccd1 _15567_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12777_ _12775_/X _12777_/B vssd1 vssd1 vccd1 vccd1 _12778_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_127_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17304_ _17621_/C _17636_/B _17301_/Y _17303_/B vssd1 vssd1 vccd1 vccd1 _17305_/B
+ sky130_fd_sc_hd__a22oi_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14516_ _14516_/A _14828_/B _16406_/A _16404_/A vssd1 vssd1 vccd1 vccd1 _14671_/A
+ sky130_fd_sc_hd__nand4_2
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18284_ _19644_/A _19227_/C _19227_/D _19487_/A vssd1 vssd1 vccd1 vccd1 _18286_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11451__A1 _11549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11728_ _11727_/B _11727_/C _11727_/A vssd1 vssd1 vccd1 vccd1 _11734_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_138_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15496_ _15496_/A _15496_/B _15496_/C vssd1 vssd1 vccd1 vccd1 _15497_/B sky130_fd_sc_hd__and3_1
XFILLER_0_86_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16743__B _16743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17235_ _17235_/A _17235_/B vssd1 vssd1 vccd1 vccd1 _17236_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_127_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14447_ _14447_/A _14913_/C vssd1 vssd1 vccd1 vccd1 _14601_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_83_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11659_ _12402_/A _13525_/A _12858_/C _12991_/D vssd1 vssd1 vccd1 vccd1 _11659_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_154_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20265__B _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17166_ _17165_/A _17165_/B _17165_/C vssd1 vssd1 vccd1 vccd1 _17169_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14378_ _14375_/X _14376_/Y _14228_/B _14230_/A vssd1 vssd1 vccd1 vccd1 _14379_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_40_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17277__D _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16117_ _15985_/X _15987_/X _16115_/Y _16116_/X vssd1 vssd1 vccd1 vccd1 _16119_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__20474__B1 _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13329_ _13188_/A _13188_/C _13188_/B vssd1 vssd1 vccd1 vccd1 _13330_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_51_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17097_ _17097_/A _17097_/B vssd1 vssd1 vccd1 vccd1 _17099_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16048_ _16273_/A _16377_/B _16048_/C _16048_/D vssd1 vssd1 vccd1 vccd1 _16165_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_86_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15375__A _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12214__D _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15806__C _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19807_ _19808_/A _19808_/B _19808_/C vssd1 vssd1 vccd1 vccd1 _19807_/X sky130_fd_sc_hd__a21o_1
XANTENNA__20431__D _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14456__A1 _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13259__A2 _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17999_ _17999_/A _17999_/B _17999_/C vssd1 vssd1 vccd1 vccd1 _18002_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12511__B _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14456__B2 _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19738_ _19737_/B _19737_/C _19737_/A vssd1 vssd1 vccd1 vccd1 _19740_/D sky130_fd_sc_hd__a21o_1
XANTENNA__16918__B _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19669_ _19669_/A _19669_/B _19669_/C vssd1 vssd1 vccd1 vccd1 _19671_/B sky130_fd_sc_hd__nand3_2
X_21700_ _22080_/CLK _21700_/D vssd1 vssd1 vccd1 vccd1 hold73/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19013__C _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21631_ _21682_/CLK _21631_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[94] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21562_ mstream_o[25] hold28/X _21562_/S vssd1 vssd1 vccd1 vccd1 _22089_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20513_ _20513_/A _20513_/B vssd1 vssd1 vccd1 vccd1 _20514_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_34_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21493_ hold179/X sstream_i[70] _21494_/S vssd1 vssd1 vccd1 vccd1 _22020_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_15_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout507_A _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20444_ _20444_/A _20444_/B vssd1 vssd1 vccd1 vccd1 _20446_/B sky130_fd_sc_hd__nor2_1
XANTENNA__20606__D _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20375_ _20901_/A _20643_/A vssd1 vssd1 vccd1 vccd1 _20513_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_28_1166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20191__A _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17915__D _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22045_ _22049_/CLK _22045_/D vssd1 vssd1 vccd1 vccd1 hold251/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_103_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18596__A _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10961_ hold36/A hold145/A vssd1 vssd1 vccd1 vccd1 _10961_/X sky130_fd_sc_hd__and2_1
XFILLER_0_134_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13670__A2 _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12700_ _12696_/X _12698_/Y _12585_/Y _12587_/X vssd1 vssd1 vccd1 vccd1 _12701_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_97_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13680_ _14138_/A _13975_/B _14477_/C _14635_/D vssd1 vssd1 vccd1 vccd1 _13835_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_97_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11681__A1 _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ _10892_/A _10892_/B vssd1 vssd1 vccd1 vccd1 _10892_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__20940__A1 _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20940__B2 _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14348__B _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12631_ _12631_/A vssd1 vssd1 vccd1 vccd1 _12631_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_155_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21829_ _21829_/CLK _21829_/D vssd1 vssd1 vccd1 vccd1 _21829_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_155_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15350_ _15350_/A _15350_/B vssd1 vssd1 vccd1 vccd1 _15351_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12562_ _12562_/A _12562_/B vssd1 vssd1 vccd1 vccd1 _12563_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_148_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17659__B _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14301_ _14301_/A _14301_/B vssd1 vssd1 vccd1 vccd1 _14443_/A sky130_fd_sc_hd__or2_1
XFILLER_0_135_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11513_ _21723_/D t1y[21] t0x[21] _11223_/A vssd1 vssd1 vccd1 vccd1 _11513_/X sky130_fd_sc_hd__a22o_1
X_15281_ _15281_/A _15281_/B vssd1 vssd1 vccd1 vccd1 _15284_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12493_ fanout9/X _12493_/B vssd1 vssd1 vccd1 vccd1 _12493_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_124_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17020_ _17144_/A _17019_/C _17124_/C _17129_/B vssd1 vssd1 vccd1 vccd1 _17021_/B
+ sky130_fd_sc_hd__a22o_1
X_14232_ _14713_/B _15098_/B _14083_/X _14084_/X _14557_/D vssd1 vssd1 vccd1 vccd1
+ _14237_/A sky130_fd_sc_hd__a32o_1
XANTENNA__14383__B1 _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11444_ _11447_/A1 hold120/A fanout48/X hold201/A vssd1 vssd1 vccd1 vccd1 _11444_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19874__B _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14163_ _14162_/B _14162_/C _14162_/A vssd1 vssd1 vccd1 vccd1 _14163_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_145_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11375_ _11447_/A1 hold260/X _11126_/B hold182/X vssd1 vssd1 vccd1 vccd1 _11375_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_150_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13114_ _13975_/B _13858_/C _13402_/D _14312_/D vssd1 vssd1 vccd1 vccd1 _13115_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14094_ _14093_/A _14093_/B _14093_/C vssd1 vssd1 vccd1 vccd1 _14095_/C sky130_fd_sc_hd__a21o_1
XANTENNA__17394__B _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18971_ _18807_/A _18807_/C _18807_/B vssd1 vssd1 vccd1 vccd1 _18972_/C sky130_fd_sc_hd__a21bo_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ _14712_/B _14384_/C _14384_/D _14712_/A vssd1 vssd1 vccd1 vccd1 _13046_/B
+ sky130_fd_sc_hd__a22oi_2
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17922_ _17921_/B _17921_/C _17921_/A vssd1 vssd1 vccd1 vccd1 _17923_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__19890__A _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17853_ _18095_/A _17853_/B vssd1 vssd1 vccd1 vccd1 _17958_/A sky130_fd_sc_hd__nor2_1
X_16804_ _16968_/C _16733_/X _16803_/X vssd1 vssd1 vccd1 vccd1 _16805_/B sky130_fd_sc_hd__a21bo_1
X_14996_ _14996_/A _14996_/B vssd1 vssd1 vccd1 vccd1 _15004_/A sky130_fd_sc_hd__xnor2_1
X_17784_ _17782_/X _17784_/B vssd1 vssd1 vccd1 vccd1 _17785_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_92_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19377__B2 _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19523_ _19524_/B _19524_/A vssd1 vssd1 vccd1 vccd1 _19640_/A sky130_fd_sc_hd__and2b_1
XANTENNA__15642__B _15643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13947_ _13948_/A _13948_/B _13948_/C _13948_/D vssd1 vssd1 vccd1 vccd1 _13947_/Y
+ sky130_fd_sc_hd__nor4_2
X_16735_ _16868_/A _16860_/C _16917_/C _16734_/B vssd1 vssd1 vccd1 vccd1 _16736_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11121__A0 _10988_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16666_ _16665_/A _16665_/C _16665_/B vssd1 vssd1 vccd1 vccd1 _16669_/B sky130_fd_sc_hd__a21o_1
X_19454_ _19300_/A _19300_/B _19298_/X vssd1 vssd1 vccd1 vccd1 _19456_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13878_ _13878_/A _13878_/B _14032_/B vssd1 vssd1 vccd1 vccd1 _13878_/X sky130_fd_sc_hd__and3_1
XFILLER_0_5_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15617_ _15614_/Y _15615_/X _15473_/B _15475_/C vssd1 vssd1 vccd1 vccd1 _15617_/X
+ sky130_fd_sc_hd__o211a_1
X_18405_ _19008_/D _19201_/B _18403_/Y _18552_/A vssd1 vssd1 vccd1 vccd1 _18405_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_12829_ _21725_/D hold163/X _11055_/Y fanout6/X _12828_/Y vssd1 vssd1 vccd1 vccd1
+ _12829_/X sky130_fd_sc_hd__a221o_1
X_16597_ _16597_/A _16597_/B vssd1 vssd1 vccd1 vccd1 _16599_/B sky130_fd_sc_hd__xnor2_2
X_19385_ _19383_/X _19385_/B vssd1 vssd1 vccd1 vccd1 _19386_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__12059__A _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15548_ _15548_/A _15548_/B vssd1 vssd1 vccd1 vccd1 _15556_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_29_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18336_ _19732_/A _19732_/B _19546_/D _19906_/C vssd1 vssd1 vccd1 vccd1 _18338_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18267_ _18267_/A _18267_/B vssd1 vssd1 vccd1 vccd1 _18270_/A sky130_fd_sc_hd__xor2_1
X_15479_ _15338_/B _15340_/A _15477_/Y _15478_/X vssd1 vssd1 vccd1 vccd1 _15481_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_126_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17218_ _17219_/A _17297_/A _17219_/C vssd1 vssd1 vccd1 vccd1 _17256_/A sky130_fd_sc_hd__and3_1
X_18198_ _19438_/B _19092_/C _19868_/B _19438_/A vssd1 vssd1 vccd1 vccd1 _18199_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17149_ _17149_/A _17149_/B vssd1 vssd1 vccd1 vccd1 _17149_/X sky130_fd_sc_hd__and2_1
Xfanout7 fanout8/X vssd1 vssd1 vccd1 vccd1 fanout7/X sky130_fd_sc_hd__buf_4
X_20160_ _20161_/A _20161_/B vssd1 vssd1 vccd1 vccd1 _20307_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_126_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20091_ _20091_/A _20091_/B vssd1 vssd1 vccd1 vccd1 _20235_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_23_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19008__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21411__A2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout192_A _21823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11112__A0 _10934_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14449__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20993_ _20994_/B _20994_/A vssd1 vssd1 vccd1 vccd1 _20993_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__17918__A2 _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15929__A1 _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15929__B2 _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout624_A _17557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21614_ _21906_/CLK _21614_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[77] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21720__D _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21545_ mstream_o[8] hold33/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22072_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14184__A _14659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17551__B1 _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14615__C _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19694__B _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21476_ hold131/X sstream_i[53] _21481_/S vssd1 vssd1 vccd1 vccd1 _22003_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20427_ _20427_/A _20427_/B vssd1 vssd1 vccd1 vccd1 _20438_/A sky130_fd_sc_hd__or2_1
XFILLER_0_120_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11160_ hold318/X _11126_/A fanout45/X hold261/A vssd1 vssd1 vccd1 vccd1 _11160_/X
+ sky130_fd_sc_hd__a22o_1
X_20358_ _20355_/Y _20356_/X _20165_/Y _20211_/Y vssd1 vssd1 vccd1 vccd1 _20358_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_12_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11091_ _11045_/X hold9/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21685_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20289_ _20290_/B _20290_/A vssd1 vssd1 vccd1 vccd1 _20440_/A sky130_fd_sc_hd__nand2b_1
X_22028_ _22038_/CLK _22028_/D vssd1 vssd1 vccd1 vccd1 hold304/A sky130_fd_sc_hd__dfxtp_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11351__B1 _11350_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
X_14850_ _14418_/A _14418_/B _14847_/X _14848_/Y vssd1 vssd1 vccd1 vccd1 _14971_/C
+ sky130_fd_sc_hd__o211ai_2
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold74 hold74/A vssd1 vssd1 vccd1 vccd1 hold74/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 hold85/A vssd1 vssd1 vccd1 vccd1 hold85/X sky130_fd_sc_hd__dlygate4sd3_1
X_13801_ _13800_/A _13800_/B _13800_/C _13800_/D vssd1 vssd1 vccd1 vccd1 _13801_/Y
+ sky130_fd_sc_hd__o22ai_4
Xhold96 hold96/A vssd1 vssd1 vccd1 vccd1 hold96/X sky130_fd_sc_hd__dlygate4sd3_1
X_14781_ _14782_/A _14782_/B vssd1 vssd1 vccd1 vccd1 _14783_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11103__A0 _10867_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11993_ _12781_/D _12512_/A vssd1 vssd1 vccd1 vccd1 _11994_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11482__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16520_ _17619_/A _17041_/A _16899_/B _17013_/C vssd1 vssd1 vccd1 vccd1 _16522_/B
+ sky130_fd_sc_hd__a22o_1
X_13732_ _13732_/A _13732_/B _13732_/C vssd1 vssd1 vccd1 vccd1 _13734_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_39_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10944_ _10945_/A _10945_/B _10945_/C vssd1 vssd1 vccd1 vccd1 _10946_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18773__B _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16451_ _17029_/A _17029_/B _16968_/C _16743_/C vssd1 vssd1 vccd1 vccd1 _16451_/X
+ sky130_fd_sc_hd__and4_1
X_13663_ _13664_/A _13964_/B vssd1 vssd1 vccd1 vccd1 _13668_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__16593__A1 _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10875_ mstream_o[46] _10874_/Y _10992_/S vssd1 vssd1 vccd1 vccd1 _21583_/D sky130_fd_sc_hd__mux2_1
XANTENNA__16593__B2 _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15402_ _15402_/A _15402_/B vssd1 vssd1 vccd1 vccd1 _15404_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19170_ hold118/X fanout7/X _14296_/Y _11550_/B vssd1 vssd1 vccd1 vccd1 _19170_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12614_ _12615_/A _12615_/B vssd1 vssd1 vccd1 vccd1 _12614_/X sky130_fd_sc_hd__and2b_1
X_16382_ _16382_/A _16382_/B vssd1 vssd1 vccd1 vccd1 _16384_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13594_ _15514_/A _15514_/B _14365_/D _14212_/C vssd1 vssd1 vccd1 vccd1 _13752_/A
+ sky130_fd_sc_hd__and4_1
X_18121_ _18121_/A _18121_/B vssd1 vssd1 vccd1 vccd1 _18122_/C sky130_fd_sc_hd__or2_1
XFILLER_0_53_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15333_ _15332_/A _15332_/B _15332_/C vssd1 vssd1 vccd1 vccd1 _15334_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13710__B _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16724__D _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12545_ _12432_/X _12434_/X _12543_/X _12544_/Y vssd1 vssd1 vccd1 vccd1 _12583_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12607__A _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18052_ _19692_/A _18789_/A _18049_/Y _18185_/A vssd1 vssd1 vccd1 vccd1 _18054_/C
+ sky130_fd_sc_hd__o2bb2a_1
X_15264_ _16404_/A _16369_/A _15264_/C _15264_/D vssd1 vssd1 vccd1 vccd1 _15400_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_124_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12476_ _12475_/A _12475_/B _12475_/C _12475_/D vssd1 vssd1 vccd1 vccd1 _12476_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_151_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12906__A1 _14712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17003_ _17002_/A _17002_/Y _16956_/Y _16964_/X vssd1 vssd1 vccd1 vccd1 _17005_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12326__B _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20429__B1 _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14215_ _14215_/A _14215_/B vssd1 vssd1 vccd1 vccd1 _14224_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12906__B2 _14712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ hold271/A fanout28/X _11426_/X vssd1 vssd1 vccd1 vccd1 _11427_/X sky130_fd_sc_hd__a21o_1
XANTENNA_5 _11319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15195_ _15195_/A _15195_/B vssd1 vssd1 vccd1 vccd1 _15196_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_21_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14146_ _14146_/A _14146_/B vssd1 vssd1 vccd1 vccd1 _14149_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ hold197/X fanout29/X _11357_/X vssd1 vssd1 vccd1 vccd1 _11358_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_123_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19109__B _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14077_ _14557_/B _14077_/B _14077_/C _14231_/A vssd1 vssd1 vccd1 vccd1 _14231_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11884__C _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18954_ _18952_/X _18954_/B vssd1 vssd1 vccd1 vccd1 _18955_/B sky130_fd_sc_hd__nand2b_1
X_11289_ _11325_/A1 t2y[16] t0y[16] _11507_/A1 vssd1 vssd1 vccd1 vccd1 _11289_/X sky130_fd_sc_hd__a22o_1
XANTENNA__12342__A _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13028_ _13148_/B _13027_/C _13027_/A vssd1 vssd1 vccd1 vccd1 _13029_/C sky130_fd_sc_hd__a21o_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17905_ _17904_/A _17904_/B _17904_/C vssd1 vssd1 vccd1 vccd1 _17906_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13157__B _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18885_ _19159_/A _18885_/B _19006_/A _18885_/D vssd1 vssd1 vccd1 vccd1 _19006_/B
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_83_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17836_ _17833_/Y _17834_/Y _17835_/X fanout2/X hold80/X vssd1 vssd1 vccd1 vccd1
+ _21892_/D sky130_fd_sc_hd__o32a_1
XANTENNA__19125__A _21824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10797__A _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21157__A1 _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17767_ _19664_/B _18624_/A _17643_/X _17642_/X _18319_/B vssd1 vssd1 vccd1 vccd1
+ _17768_/C sky130_fd_sc_hd__a32o_1
X_14979_ _15076_/A _15076_/B _16380_/B _16173_/B vssd1 vssd1 vccd1 vccd1 _15075_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__11392__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19506_ _20462_/D _20733_/C _20606_/D _20026_/B vssd1 vssd1 vccd1 vccd1 _19509_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16718_ _16718_/A _16718_/B _16718_/C vssd1 vssd1 vccd1 vccd1 _16718_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__15091__C _15091_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17698_ _17698_/A _17698_/B _17698_/C vssd1 vssd1 vccd1 vccd1 _17700_/A sky130_fd_sc_hd__or3_1
XFILLER_0_53_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19437_ _19438_/B _20247_/C _20247_/D _19438_/A vssd1 vssd1 vccd1 vccd1 _19441_/A
+ sky130_fd_sc_hd__a22o_1
X_16649_ _16648_/A _16648_/C _16648_/B vssd1 vssd1 vccd1 vccd1 _16653_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_92_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19368_ _19368_/A _19368_/B vssd1 vssd1 vccd1 vccd1 _19370_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__21314__D1 _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14716__B _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20668__B1 _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13620__B _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18319_ _19535_/A _18319_/B _18622_/B _19089_/B vssd1 vssd1 vccd1 vccd1 _18320_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_127_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19299_ _19299_/A _19299_/B vssd1 vssd1 vccd1 vccd1 _19300_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__14347__B1 _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21330_ _21349_/A _11549_/A _11089_/A vssd1 vssd1 vccd1 vccd1 _21390_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_5_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11778__D _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21261_ _21261_/A _21261_/B vssd1 vssd1 vccd1 vccd1 _21263_/A sky130_fd_sc_hd__or2_1
XANTENNA__19286__B1 _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout205_A _19751_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13570__A1 _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20212_ _20212_/A _20212_/B vssd1 vssd1 vccd1 vccd1 _20215_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13570__B2 _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21192_ _21293_/A _21291_/B vssd1 vssd1 vccd1 vccd1 _21193_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20143_ _20143_/A _20143_/B vssd1 vssd1 vccd1 vccd1 _20153_/A sky130_fd_sc_hd__or2_1
XFILLER_0_111_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20074_ _20075_/A _20075_/B vssd1 vssd1 vccd1 vccd1 _20224_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17762__B _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout574_A _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13873__A2 _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16203__A_N _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20976_ _20583_/A _21293_/B _21261_/B _20845_/D vssd1 vssd1 vccd1 vccd1 _20978_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_79_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout20_A _11224_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12427__A _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12330_ _12330_/A _12330_/B vssd1 vssd1 vccd1 vccd1 _12332_/B sky130_fd_sc_hd__and2_1
XFILLER_0_63_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21528_ hold270/X sstream_i[105] _21528_/S vssd1 vssd1 vccd1 vccd1 _22055_/D sky130_fd_sc_hd__mux2_1
XANTENNA__16878__A2 _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11688__D _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12261_ _12261_/A _12269_/B _12268_/B _12269_/C vssd1 vssd1 vccd1 vccd1 _12261_/X
+ sky130_fd_sc_hd__and4_1
X_21459_ hold177/X sstream_i[36] _21494_/S vssd1 vssd1 vccd1 vccd1 _21986_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14000_ _14000_/A _14000_/B _14153_/B vssd1 vssd1 vccd1 vccd1 _14002_/B sky130_fd_sc_hd__nand3_2
X_11212_ hold181/X fanout22/X _11211_/X vssd1 vssd1 vccd1 vccd1 _11212_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16560__C _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12192_ _12185_/A _12185_/B _12185_/C vssd1 vssd1 vccd1 vccd1 _12193_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_43_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13258__A _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19029__B1 _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ hold139/X fanout23/X _11142_/X vssd1 vssd1 vccd1 vccd1 _11143_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15302__A2 _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12162__A _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15951_ _15948_/Y _15949_/X _15784_/B _15823_/X vssd1 vssd1 vccd1 vccd1 _15999_/B
+ sky130_fd_sc_hd__o211a_1
X_11074_ _10892_/Y hold48/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21669_/D sky130_fd_sc_hd__mux2_1
XANTENNA__11324__A0 _14477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13408__D _14663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16569__A _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14902_ _14751_/A _14751_/B _14749_/Y vssd1 vssd1 vccd1 vccd1 _14904_/B sky130_fd_sc_hd__a21boi_2
X_15882_ _15708_/Y _15711_/Y _16011_/A _15881_/X vssd1 vssd1 vccd1 vccd1 _16011_/B
+ sky130_fd_sc_hd__a211oi_2
X_18670_ _18669_/A _18669_/B _18669_/C _18669_/D vssd1 vssd1 vccd1 vccd1 _18670_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_99_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17621_ _17737_/A _17620_/Y _17621_/C _17741_/B vssd1 vssd1 vccd1 vccd1 _17737_/B
+ sky130_fd_sc_hd__and4bb_1
X_14833_ _14833_/A _14833_/B _14833_/C vssd1 vssd1 vccd1 vccd1 _14836_/A sky130_fd_sc_hd__nand3_1
XANTENNA__13705__B _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14089__A _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14764_ _14764_/A _14764_/B vssd1 vssd1 vccd1 vccd1 _14901_/A sky130_fd_sc_hd__or2_1
X_17552_ _17915_/A _19587_/A _19587_/B _17915_/D vssd1 vssd1 vccd1 vccd1 _17552_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_153_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11976_ _11976_/A _11976_/B vssd1 vssd1 vccd1 vccd1 _11979_/B sky130_fd_sc_hd__and2_1
XANTENNA__19752__A1 _21833_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13715_ _13716_/A _13716_/B vssd1 vssd1 vccd1 vccd1 _13846_/A sky130_fd_sc_hd__nand2_1
X_16503_ _16503_/A _17197_/A _16503_/C vssd1 vssd1 vccd1 vccd1 _16553_/A sky130_fd_sc_hd__or3_2
XFILLER_0_156_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17483_ _17483_/A _17483_/B _17483_/C _17483_/D vssd1 vssd1 vccd1 vccd1 _17484_/B
+ sky130_fd_sc_hd__nand4_1
X_10927_ mstream_o[53] _10926_/X _10992_/S vssd1 vssd1 vccd1 vccd1 _21590_/D sky130_fd_sc_hd__mux2_1
XANTENNA__15369__A2 _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14695_ _16027_/A _16328_/A vssd1 vssd1 vccd1 vccd1 _14696_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_50_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14817__A _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19222_ _18732_/C _19221_/X _19220_/X vssd1 vssd1 vccd1 vccd1 _19224_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_156_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16434_ _16434_/A _16434_/B vssd1 vssd1 vccd1 vccd1 _16435_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13646_ _13643_/X _13644_/Y _13491_/C _13490_/Y vssd1 vssd1 vccd1 vccd1 _13648_/D
+ sky130_fd_sc_hd__a211oi_4
X_10858_ _10859_/A _10859_/B _10859_/C vssd1 vssd1 vccd1 vccd1 _10866_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_39_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18008__B _18008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13440__B _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16365_ hold92/X _16364_/X fanout1/X vssd1 vssd1 vccd1 vccd1 hold93/A sky130_fd_sc_hd__mux2_1
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19153_ _19152_/B _19152_/C _19152_/A vssd1 vssd1 vccd1 vccd1 _19154_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13577_ _13578_/A _13578_/B vssd1 vssd1 vccd1 vccd1 _13732_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15316_ _15316_/A _15316_/B vssd1 vssd1 vccd1 vccd1 _15326_/A sky130_fd_sc_hd__or2_1
X_18104_ hold58/X _18103_/X fanout3/X vssd1 vssd1 vccd1 vccd1 _21894_/D sky130_fd_sc_hd__mux2_1
X_12528_ _12750_/A _12528_/B _13152_/C _13152_/D vssd1 vssd1 vccd1 vccd1 _12530_/C
+ sky130_fd_sc_hd__nand4_2
X_16296_ _16297_/A _16297_/B vssd1 vssd1 vccd1 vccd1 _16296_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_125_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19084_ _19084_/A _19084_/B vssd1 vssd1 vccd1 vccd1 _19103_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15648__A _15907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15247_ _15247_/A _15247_/B vssd1 vssd1 vccd1 vccd1 _15249_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_clkbuf_leaf_10_clk_i_A _21806_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18035_ _19892_/A _18624_/A _18175_/A _18035_/D vssd1 vssd1 vccd1 vccd1 _18175_/B
+ sky130_fd_sc_hd__nand4_1
X_12459_ _12357_/C _13034_/D _14386_/B _12458_/A vssd1 vssd1 vccd1 vccd1 _12460_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20273__B _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16470__C _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15178_ _15177_/B _15177_/C _15177_/A vssd1 vssd1 vccd1 vccd1 _15179_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_1_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11563__B1 _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14129_ hold140/X _14128_/X fanout4/X vssd1 vssd1 vccd1 vccd1 hold141/A sky130_fd_sc_hd__mux2_1
Xfanout309 _17490_/A vssd1 vssd1 vccd1 vccd1 _17123_/C sky130_fd_sc_hd__buf_4
X_19986_ _19885_/B _19884_/Y _19983_/Y _20122_/B vssd1 vssd1 vccd1 vccd1 _20164_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18937_ _18775_/A _18775_/C _18775_/B vssd1 vssd1 vccd1 vccd1 _18938_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__11315__B1 _11314_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18868_ _19650_/D _18849_/A _19030_/C _21847_/Q _18713_/X vssd1 vssd1 vccd1 vccd1
+ _18876_/A sky130_fd_sc_hd__a41o_1
XFILLER_0_119_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18794__A2 _19751_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17819_ _17819_/A _17819_/B _17819_/C vssd1 vssd1 vccd1 vccd1 _17821_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_55_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18799_ _19445_/A _19972_/C vssd1 vssd1 vccd1 vccd1 _18802_/A sky130_fd_sc_hd__and2_1
XFILLER_0_55_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20830_ _20830_/A _20830_/B _20830_/C vssd1 vssd1 vccd1 vccd1 _20830_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20761_ _20630_/Y _20632_/Y _20759_/Y _20760_/X vssd1 vssd1 vccd1 vccd1 _20896_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_147_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14727__A _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout155_A _21830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20692_ _20692_/A _20808_/B vssd1 vssd1 vccd1 vccd1 _20694_/B sky130_fd_sc_hd__or2_1
XFILLER_0_92_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout322_A _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20105__A2 _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17757__B _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21313_ _21176_/A _21176_/B _21179_/A vssd1 vssd1 vccd1 vccd1 _21317_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21244_ _21244_/A _21244_/B _21244_/C vssd1 vssd1 vccd1 vccd1 _21246_/A sky130_fd_sc_hd__nor3_1
Xhold330 hold330/A vssd1 vssd1 vccd1 vccd1 hold330/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19972__B _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14181__B _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18482__A1 _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21175_ _21270_/S _21175_/B vssd1 vssd1 vccd1 vccd1 _21176_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_1_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19691__C _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20126_ _20126_/A _20126_/B vssd1 vssd1 vccd1 vccd1 _20159_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_99_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20057_ _19830_/X _19832_/Y _20203_/B _20056_/Y vssd1 vssd1 vccd1 vccd1 _20167_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18785__A2 _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13525__B _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_203 hold268/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11830_ _11833_/B _11830_/B _11830_/C _11830_/D vssd1 vssd1 vccd1 vccd1 _11830_/Y
+ sky130_fd_sc_hd__nand4_2
XTAP_3269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_214 hold275/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_225 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_236 hold299/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_247 _11347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_258 hold262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11761_ _11761_/A _11761_/B _11761_/C vssd1 vssd1 vccd1 vccd1 _11764_/A sky130_fd_sc_hd__nand3_1
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_269 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20959_ _20955_/X _20956_/Y _20822_/Y _20824_/X vssd1 vssd1 vccd1 vccd1 _20960_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_56_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14637__A _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ _13523_/B _13501_/B _13500_/C _13500_/D vssd1 vssd1 vccd1 vccd1 _13500_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17013__A _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14480_ _14480_/A _14480_/B _14632_/B vssd1 vssd1 vccd1 vccd1 _14482_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_82_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11692_ _12750_/A _12528_/B _12020_/A _12326_/D vssd1 vssd1 vccd1 vccd1 _12330_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13898__D _14218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13431_ _13428_/Y _13429_/X _13306_/B _13306_/Y vssd1 vssd1 vccd1 vccd1 _13431_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__13260__B _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19866__C _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16150_ _16150_/A _16150_/B vssd1 vssd1 vccd1 vccd1 _16151_/B sky130_fd_sc_hd__xor2_2
XANTENNA__14075__C _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13362_ _13512_/A _13361_/C _13361_/A vssd1 vssd1 vccd1 vccd1 _13363_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_24_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18170__B1 _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15101_ _15101_/A _15226_/A _15101_/C vssd1 vssd1 vccd1 vccd1 _15226_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_107_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12313_ _12313_/A _12313_/B vssd1 vssd1 vccd1 vccd1 _12315_/B sky130_fd_sc_hd__xnor2_2
X_16081_ _15909_/B _15948_/Y _16079_/X _16080_/Y vssd1 vssd1 vccd1 vccd1 _16128_/A
+ sky130_fd_sc_hd__o211ai_4
X_13293_ _14365_/A _15514_/A _15514_/B _14367_/A vssd1 vssd1 vccd1 vccd1 _13293_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_146_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15032_ _15931_/A _15931_/B _16328_/A _16326_/A vssd1 vssd1 vccd1 vccd1 _15127_/A
+ sky130_fd_sc_hd__nand4_1
X_12244_ _12217_/A _12217_/C _12217_/B vssd1 vssd1 vccd1 vccd1 _12244_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17276__A2 _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19840_ _19840_/A _19840_/B vssd1 vssd1 vccd1 vccd1 _19841_/B sky130_fd_sc_hd__xnor2_1
X_12175_ _12175_/A _12175_/B vssd1 vssd1 vccd1 vccd1 _12175_/Y sky130_fd_sc_hd__xnor2_1
X_11126_ _11126_/A _11126_/B vssd1 vssd1 vccd1 vccd1 _11126_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_43_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19771_ _19772_/A _19772_/B vssd1 vssd1 vccd1 vccd1 _19771_/Y sky130_fd_sc_hd__nor2_1
X_16983_ _16983_/A _16983_/B vssd1 vssd1 vccd1 vccd1 _16986_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_120_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18722_ _18719_/Y _18720_/X _18559_/A _18560_/Y vssd1 vssd1 vccd1 vccd1 _18722_/X
+ sky130_fd_sc_hd__o211a_1
X_15934_ _15934_/A _16056_/B vssd1 vssd1 vccd1 vccd1 _15936_/B sky130_fd_sc_hd__or2_1
X_11057_ _11057_/A _11057_/B vssd1 vssd1 vccd1 vccd1 _11057_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_155_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19973__A1 _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18653_ _18653_/A _18653_/B _18653_/C vssd1 vssd1 vccd1 vccd1 _18656_/A sky130_fd_sc_hd__nand3_1
X_15865_ _15726_/X _15728_/X _15863_/Y _15864_/X vssd1 vssd1 vccd1 vccd1 _15867_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_153_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15931__A _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17604_ _17493_/A _21151_/A _18894_/B _18703_/A vssd1 vssd1 vccd1 vccd1 _17605_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14816_ _16084_/A _15717_/B _15791_/A _14817_/D vssd1 vssd1 vccd1 vccd1 _14816_/X
+ sky130_fd_sc_hd__and4_1
X_18584_ _19051_/A _20317_/D _19057_/C _19057_/D vssd1 vssd1 vccd1 vccd1 _18584_/X
+ sky130_fd_sc_hd__and4_1
XTAP_3770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15796_ _15796_/A _15796_/B vssd1 vssd1 vccd1 vccd1 _15798_/B sky130_fd_sc_hd__or2_1
XFILLER_0_114_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17535_ _17536_/A _17536_/B _17536_/C vssd1 vssd1 vccd1 vccd1 _17535_/X sky130_fd_sc_hd__a21o_2
X_14747_ _14747_/A _14747_/B vssd1 vssd1 vccd1 vccd1 _14750_/A sky130_fd_sc_hd__xor2_4
XANTENNA__16539__A1 _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11959_ _11960_/A _11960_/B _11960_/C vssd1 vssd1 vccd1 vccd1 _11969_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__19122__B _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14678_ _14677_/B _14825_/B _14677_/A vssd1 vssd1 vccd1 vccd1 _14679_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_15_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17466_ _17466_/A _17466_/B _17466_/C _17466_/D vssd1 vssd1 vccd1 vccd1 _17466_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_74_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15211__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19205_ _19204_/B _19204_/C _19204_/A vssd1 vssd1 vccd1 vccd1 _19206_/C sky130_fd_sc_hd__a21o_1
XANTENNA__18961__B _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16417_ _16328_/A _21784_/Q _16329_/A _16327_/B vssd1 vssd1 vccd1 vccd1 _16421_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13629_ _13475_/A _13475_/C _13475_/B vssd1 vssd1 vccd1 vccd1 _13630_/C sky130_fd_sc_hd__a21bo_1
X_17397_ _17395_/X _17397_/B vssd1 vssd1 vccd1 vccd1 _17398_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_73_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19136_ _19135_/B _19135_/C _19135_/A vssd1 vssd1 vccd1 vccd1 _19136_/Y sky130_fd_sc_hd__a21oi_2
X_16348_ _16348_/A _16348_/B vssd1 vssd1 vccd1 vccd1 _16349_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_82_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18700__A2 _19181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16279_ _16279_/A vssd1 vssd1 vccd1 vccd1 _16293_/A sky130_fd_sc_hd__inv_2
XANTENNA__21099__B _21311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19067_ _19692_/A _19068_/C _20146_/B _19535_/B vssd1 vssd1 vccd1 vccd1 _19070_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14713__C _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18018_ _18018_/A _18018_/B _18018_/C vssd1 vssd1 vccd1 vccd1 _18020_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_11_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18689__A _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout106 _21841_/Q vssd1 vssd1 vccd1 vccd1 _19691_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout117 _21169_/A vssd1 vssd1 vccd1 vccd1 _17739_/D sky130_fd_sc_hd__buf_4
XFILLER_0_61_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout128 _21836_/Q vssd1 vssd1 vccd1 vccd1 _20910_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_129_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout139 _18929_/B vssd1 vssd1 vccd1 vccd1 _20101_/A sky130_fd_sc_hd__buf_4
X_19969_ _20103_/A _21153_/B vssd1 vssd1 vccd1 vccd1 _19970_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18201__B _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19413__B1 _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12530__A _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21931_ _21942_/CLK _21931_/D vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21862_ _21932_/CLK _21862_/D vssd1 vssd1 vccd1 vccd1 hold219/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20813_ _21171_/A _21278_/B _20811_/Y _20938_/A vssd1 vssd1 vccd1 vccd1 _20815_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_78_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19032__B _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14457__A _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17727__B1 _19691_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21793_ _22016_/CLK _21793_/D vssd1 vssd1 vccd1 vccd1 _21793_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_132_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout537_A _15439_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20178__B _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20744_ _20741_/Y _20742_/X _20610_/Y _20612_/Y vssd1 vssd1 vccd1 vccd1 _20744_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19967__B _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14176__B _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18871__B _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20675_ _20801_/A vssd1 vssd1 vccd1 vccd1 _20677_/D sky130_fd_sc_hd__inv_2
XFILLER_0_80_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19686__C _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16391__B _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20922__A _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21227_ _21228_/A _21228_/B _21228_/C vssd1 vssd1 vccd1 vccd1 _21229_/A sky130_fd_sc_hd__o21a_1
Xhold160 hold160/A vssd1 vssd1 vccd1 vccd1 hold160/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 hold171/A vssd1 vssd1 vccd1 vccd1 hold171/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19652__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold182 hold182/A vssd1 vssd1 vccd1 vccd1 hold182/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12143__C _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 hold193/A vssd1 vssd1 vccd1 vccd1 hold193/X sky130_fd_sc_hd__dlygate4sd3_1
X_21158_ _21256_/A _21278_/B vssd1 vssd1 vccd1 vccd1 _21159_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18749__D _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout640 _11041_/A vssd1 vssd1 vccd1 vccd1 fanout640/X sky130_fd_sc_hd__clkbuf_8
X_20109_ _20109_/A _20251_/B vssd1 vssd1 vccd1 vccd1 _20112_/A sky130_fd_sc_hd__nor2_1
X_13980_ _13980_/A _14142_/B _13981_/B vssd1 vssd1 vccd1 vccd1 _14149_/A sky130_fd_sc_hd__or3_1
X_21089_ _21206_/A _21089_/B vssd1 vssd1 vccd1 vccd1 _21090_/B sky130_fd_sc_hd__nor2_1
XTAP_3000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12931_ _12803_/C _12802_/Y _12929_/X _12930_/Y vssd1 vssd1 vccd1 vccd1 _12931_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_3011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13970__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15650_ _15650_/A _15650_/B vssd1 vssd1 vccd1 vccd1 _15689_/A sky130_fd_sc_hd__or2_1
XTAP_3055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12862_ _12862_/A _12989_/B _12862_/C vssd1 vssd1 vccd1 vccd1 _12862_/X sky130_fd_sc_hd__and3_1
XANTENNA__19223__A _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15441__B2 _21735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14601_ _14296_/B _14601_/B _14601_/C vssd1 vssd1 vccd1 vccd1 _14603_/C sky130_fd_sc_hd__and3b_1
X_11813_ _11813_/A _11813_/B _11813_/C vssd1 vssd1 vccd1 vccd1 _11816_/A sky130_fd_sc_hd__nand3_1
XTAP_3099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15581_ _15712_/A _15581_/B vssd1 vssd1 vccd1 vccd1 _15582_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_96_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12793_ _12792_/B _12792_/C _12792_/A vssd1 vssd1 vccd1 vccd1 _12795_/B sky130_fd_sc_hd__a21o_1
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14367__A _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20088__B _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14532_ _14532_/A _14532_/B vssd1 vssd1 vccd1 vccd1 _14551_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17320_ _17316_/X _17317_/Y _17212_/X _17214_/X vssd1 vssd1 vccd1 vccd1 _17356_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11744_ _11744_/A _11744_/B _11744_/C vssd1 vssd1 vccd1 vccd1 _11748_/A sky130_fd_sc_hd__nand3_2
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14463_ _14312_/D _16406_/B _16314_/D _14463_/D vssd1 vssd1 vccd1 vccd1 _14466_/A
+ sky130_fd_sc_hd__and4b_2
X_17251_ _17251_/A _17251_/B _17251_/C vssd1 vssd1 vccd1 vccd1 _17251_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_138_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11675_ _12094_/A _12444_/B _12443_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _11676_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16202_ _16202_/A _16202_/B vssd1 vssd1 vccd1 vccd1 _16206_/A sky130_fd_sc_hd__xnor2_4
X_13414_ _13415_/A _13415_/B vssd1 vssd1 vccd1 vccd1 _13539_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_107_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17182_ _17490_/A _17739_/C _17739_/D _17282_/A vssd1 vssd1 vccd1 vccd1 _17183_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14394_ _14393_/A _14393_/B _14393_/C vssd1 vssd1 vccd1 vccd1 _14395_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_119_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16133_ _16134_/A _16134_/B _16134_/C vssd1 vssd1 vccd1 vccd1 _16133_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_141_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ _13204_/B _13203_/Y _13343_/X _13344_/Y vssd1 vssd1 vccd1 vccd1 _13348_/B
+ sky130_fd_sc_hd__o211a_2
XANTENNA__12037__D _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13530__A2_N _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18694__A1 _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18694__B2 _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16064_ _16064_/A _16064_/B _16064_/C vssd1 vssd1 vccd1 vccd1 _16064_/X sky130_fd_sc_hd__and3_1
XFILLER_0_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13276_ _13427_/A _13275_/C _13275_/A vssd1 vssd1 vccd1 vccd1 _13278_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_121_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15015_ _16087_/A _15653_/C _15112_/D _16092_/D vssd1 vssd1 vccd1 vccd1 _15017_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14180__A1 _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12227_ _12226_/B _12226_/C _12226_/A vssd1 vssd1 vccd1 vccd1 _12228_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__14180__B2 _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19643__B1 _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14830__A _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14461__A1_N _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19823_ _19823_/A _20590_/D _20733_/C _20606_/D vssd1 vssd1 vccd1 vccd1 _20043_/A
+ sky130_fd_sc_hd__nand4_2
X_12158_ _12150_/A _12150_/B _12150_/C vssd1 vssd1 vccd1 vccd1 _12160_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__20734__A2_N _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20270__C _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11109_ _10912_/X hold144/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21703_/D sky130_fd_sc_hd__mux2_1
X_19754_ _19572_/Y _19574_/X _19752_/X _19753_/Y vssd1 vssd1 vccd1 vccd1 _19756_/B
+ sky130_fd_sc_hd__o211ai_4
X_16966_ _16930_/A _16930_/C _16930_/B vssd1 vssd1 vccd1 vccd1 _16982_/B sky130_fd_sc_hd__a21o_1
X_12089_ _12268_/A _12512_/A vssd1 vssd1 vccd1 vccd1 _12091_/B sky130_fd_sc_hd__and2_1
XANTENNA__19946__A1 _19636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18705_ _18705_/A _18705_/B vssd1 vssd1 vccd1 vccd1 _18707_/B sky130_fd_sc_hd__xor2_1
XANTENNA__18956__B _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15917_ _16050_/A vssd1 vssd1 vccd1 vccd1 _15919_/D sky130_fd_sc_hd__inv_2
XANTENNA__19946__B2 _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17860__B _19060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19685_ _19686_/A _21278_/A _20265_/D _19892_/A vssd1 vssd1 vccd1 vccd1 _19685_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12494__A1 _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16897_ _17206_/B _18859_/A _16830_/Y _16832_/B vssd1 vssd1 vccd1 vccd1 _16898_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_56_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12494__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15661__A _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17421__A2 _20249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18636_ _19723_/A _19262_/C _18495_/B _18493_/X vssd1 vssd1 vccd1 vccd1 _18641_/A
+ sky130_fd_sc_hd__a31o_1
X_15848_ _15848_/A _15848_/B vssd1 vssd1 vccd1 vccd1 _15859_/A sky130_fd_sc_hd__or2_1
XANTENNA__14235__A2 _15093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18567_ _18563_/A _18564_/X _18409_/A _18410_/Y vssd1 vssd1 vccd1 vccd1 _18567_/X
+ sky130_fd_sc_hd__o211a_1
X_15779_ _16036_/A _15780_/B vssd1 vssd1 vccd1 vccd1 _15781_/A sky130_fd_sc_hd__and2_1
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13181__A _14712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13994__A1 _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17518_ _17405_/B _17405_/Y _17602_/A _17517_/Y vssd1 vssd1 vccd1 vccd1 _17602_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_86_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18498_ _19123_/A _18498_/B _19872_/C _19972_/C vssd1 vssd1 vccd1 vccd1 _18500_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_28_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17449_ _17557_/B _17924_/B _17670_/B _17557_/A vssd1 vssd1 vccd1 vccd1 _17450_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20460_ _20460_/A _20460_/B vssd1 vssd1 vccd1 vccd1 _20461_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11757__B1 _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19119_ _19439_/A _20242_/C vssd1 vssd1 vccd1 vccd1 _19120_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_15_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20391_ _20391_/A _20559_/B vssd1 vssd1 vccd1 vccd1 _20399_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13761__A4 _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15499__A1 _12291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout118_A _20562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22061_ _22063_/CLK _22061_/D vssd1 vssd1 vccd1 vccd1 hold268/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__12182__B1 _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21012_ _21012_/A _21012_/B _21012_/C vssd1 vssd1 vccd1 vccd1 _21014_/A sky130_fd_sc_hd__or3_1
XFILLER_0_26_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15555__B _15556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout487_A _21747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17660__A2 _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15671__A1 _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15671__B2 _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21914_ _21949_/CLK _21914_/D vssd1 vssd1 vccd1 vccd1 hold100/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__17412__A2 _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21723__D _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21845_ _21845_/CLK _21845_/D vssd1 vssd1 vccd1 vccd1 _21845_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15974__A2 _16396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11604__A _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21776_ _21822_/CLK _21776_/D vssd1 vssd1 vccd1 vccd1 _21776_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_154_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20727_ _20728_/A _20728_/B vssd1 vssd1 vccd1 vccd1 _20727_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_135_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11460_ _21718_/D t2x[3] v1z[3] fanout17/X _11459_/X vssd1 vssd1 vccd1 vccd1 _11460_/X
+ sky130_fd_sc_hd__a221o_1
X_20658_ _20658_/A _20912_/A vssd1 vssd1 vccd1 vccd1 _20660_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_135_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11391_ hold303/X fanout29/X _11390_/X vssd1 vssd1 vccd1 vccd1 _11391_/X sky130_fd_sc_hd__a21o_1
X_20589_ _20589_/A _20589_/B vssd1 vssd1 vccd1 vccd1 _20594_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14353__C _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13130_ _13867_/A _13858_/A _13269_/C _13269_/D vssd1 vssd1 vccd1 vccd1 _13267_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_108_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13061_ _13062_/A _13062_/B _13062_/C vssd1 vssd1 vccd1 vccd1 _13061_/X sky130_fd_sc_hd__and3_1
XANTENNA__18428__A1 _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12012_ _11941_/A _11941_/B _11941_/C vssd1 vssd1 vccd1 vccd1 _12012_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11993__B _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11485__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11920__B1 _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15111__B1 _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16820_ _16820_/A _16820_/B vssd1 vssd1 vccd1 vccd1 _16822_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_136_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout470 _15091_/C vssd1 vssd1 vccd1 vccd1 _14234_/C sky130_fd_sc_hd__clkbuf_8
Xfanout481 _21749_/Q vssd1 vssd1 vccd1 vccd1 _14217_/D sky130_fd_sc_hd__buf_4
Xfanout492 _16409_/A vssd1 vssd1 vccd1 vccd1 _16305_/B sky130_fd_sc_hd__buf_4
X_16751_ _16751_/A _16751_/B vssd1 vssd1 vccd1 vccd1 _16753_/B sky130_fd_sc_hd__xor2_2
X_13963_ _13813_/A _13668_/A _13813_/B vssd1 vssd1 vccd1 vccd1 _13966_/A sky130_fd_sc_hd__a21oi_2
X_15702_ _15435_/A _15838_/B _16314_/D _15702_/D vssd1 vssd1 vccd1 vccd1 _15705_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_88_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12914_ _12913_/B _12913_/C _12913_/A vssd1 vssd1 vccd1 vccd1 _12916_/B sky130_fd_sc_hd__a21o_1
X_19470_ _19318_/A _19318_/B _19317_/A vssd1 vssd1 vccd1 vccd1 _19472_/B sky130_fd_sc_hd__a21oi_2
X_13894_ _14365_/D _13893_/X _13892_/X vssd1 vssd1 vccd1 vccd1 _13896_/A sky130_fd_sc_hd__a21bo_1
X_16682_ _16682_/A _16682_/B _16682_/C vssd1 vssd1 vccd1 vccd1 _16682_/X sky130_fd_sc_hd__or3_2
X_18421_ _18420_/A _18420_/B _18543_/A _18420_/D vssd1 vssd1 vccd1 vccd1 _18421_/X
+ sky130_fd_sc_hd__o22a_1
X_15633_ _15803_/A vssd1 vssd1 vccd1 vccd1 _15635_/D sky130_fd_sc_hd__inv_2
X_12845_ _14138_/A _13975_/B _13258_/C _13258_/D vssd1 vssd1 vccd1 vccd1 _12984_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12779__A2 _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18352_ _18352_/A _18352_/B _18352_/C vssd1 vssd1 vccd1 vccd1 _18355_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_69_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15564_ _15561_/X _15562_/Y _15381_/Y _15386_/B vssd1 vssd1 vccd1 vccd1 _15564_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ _12896_/B _12774_/X _12669_/X _12672_/A vssd1 vssd1 vccd1 vccd1 _12777_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17303_ _17393_/A _17303_/B _17621_/C _17636_/B vssd1 vssd1 vccd1 vccd1 _17393_/B
+ sky130_fd_sc_hd__and4b_1
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14515_ _14365_/C _16406_/A _16404_/A _16173_/A vssd1 vssd1 vccd1 vccd1 _14518_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11727_ _11727_/A _11727_/B _11727_/C vssd1 vssd1 vccd1 vccd1 _11734_/A sky130_fd_sc_hd__nand3_1
X_15495_ _15496_/B _15496_/C _15496_/A vssd1 vssd1 vccd1 vccd1 _15625_/B sky130_fd_sc_hd__a21oi_1
X_18283_ _19487_/B _19382_/B vssd1 vssd1 vccd1 vccd1 _18287_/A sky130_fd_sc_hd__nand2_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16743__C _16743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17234_ _17334_/B _18166_/A _17666_/A _17443_/D vssd1 vssd1 vccd1 vccd1 _17235_/B
+ sky130_fd_sc_hd__and4_1
X_14446_ _14446_/A _14446_/B _14446_/C vssd1 vssd1 vccd1 vccd1 _14913_/C sky130_fd_sc_hd__nor3_2
X_11658_ _12402_/B _12312_/A vssd1 vssd1 vccd1 vccd1 _11662_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20265__C _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14377_ _14228_/B _14230_/A _14375_/X _14376_/Y vssd1 vssd1 vccd1 vccd1 _14379_/B
+ sky130_fd_sc_hd__a211o_1
X_17165_ _17165_/A _17165_/B _17165_/C vssd1 vssd1 vccd1 vccd1 _17169_/A sky130_fd_sc_hd__and3_1
XANTENNA__12400__A1 _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11589_ _13012_/B _12302_/A _11589_/C _11589_/D vssd1 vssd1 vccd1 vccd1 _11591_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__20474__A1 _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16116_ _16113_/Y _16114_/X _15980_/Y _15982_/Y vssd1 vssd1 vccd1 vccd1 _16116_/X
+ sky130_fd_sc_hd__o211a_1
X_13328_ _13327_/B _13327_/C _13327_/A vssd1 vssd1 vccd1 vccd1 _13330_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20474__B2 _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17096_ _17096_/A _17146_/D _17097_/A vssd1 vssd1 vccd1 vccd1 _17096_/X sky130_fd_sc_hd__and3_1
XANTENNA__20562__A _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16047_ _16273_/A _16377_/B _16048_/C _16048_/D vssd1 vssd1 vccd1 vccd1 _16049_/A
+ sky130_fd_sc_hd__a22oi_1
X_13259_ _13858_/B _13258_/C _13258_/D _13860_/A vssd1 vssd1 vccd1 vccd1 _13260_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15806__D _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11395__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21622__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19806_ _19808_/A _19808_/B _19808_/C vssd1 vssd1 vccd1 vccd1 _19809_/A sky130_fd_sc_hd__a21oi_1
X_17998_ _19487_/B _19227_/C _19227_/D _18873_/A vssd1 vssd1 vccd1 vccd1 _17999_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14456__A2 _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21393__A _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19737_ _19737_/A _19737_/B _19737_/C vssd1 vssd1 vccd1 vccd1 _19740_/C sky130_fd_sc_hd__nand3_1
X_16949_ _16956_/A vssd1 vssd1 vccd1 vccd1 _16949_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16487__A _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19668_ _19667_/B _19820_/B _19667_/A vssd1 vssd1 vccd1 vccd1 _19669_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_95_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18619_ _19686_/A _18769_/B vssd1 vssd1 vccd1 vccd1 _18620_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_133_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15956__A2 _21787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19599_ _19441_/A _19441_/C _19441_/B vssd1 vssd1 vccd1 vccd1 _19604_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_48_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21630_ _21682_/CLK _21630_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[93] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_47_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21561_ mstream_o[24] hold43/X _21562_/S vssd1 vssd1 vccd1 vccd1 _22088_/D sky130_fd_sc_hd__mux2_1
X_20512_ _20643_/B vssd1 vssd1 vccd1 vccd1 _20901_/B sky130_fd_sc_hd__inv_2
XFILLER_0_74_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21492_ hold186/X sstream_i[69] _21494_/S vssd1 vssd1 vccd1 vccd1 _22019_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_144_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20443_ _20441_/B _20441_/C _20441_/A vssd1 vssd1 vccd1 vccd1 _20444_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout402_A _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20374_ _19792_/B _20081_/Y _20372_/X _20373_/X vssd1 vssd1 vccd1 vccd1 _20901_/A
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_24_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20191__B _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21718__D _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22044_ _22049_/CLK _22044_/D vssd1 vssd1 vccd1 vccd1 hold237/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18596__B _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10960_ mstream_o[58] _10959_/Y _10992_/S vssd1 vssd1 vccd1 vccd1 _21595_/D sky130_fd_sc_hd__mux2_1
XANTENNA_fanout50_A _11122_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13407__B1 _14663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10891_ hold243/A hold252/A _10886_/A vssd1 vssd1 vccd1 vccd1 _10892_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11681__A2 _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14348__C _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12630_ _12630_/A _12630_/B _12630_/C vssd1 vssd1 vccd1 vccd1 _12631_/A sky130_fd_sc_hd__and3_2
X_21828_ _21829_/CLK _21828_/D vssd1 vssd1 vccd1 vccd1 _21828_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18346__B1 _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12561_ _13173_/C _12780_/A _12780_/B _13155_/A vssd1 vssd1 vccd1 vccd1 _12562_/B
+ sky130_fd_sc_hd__a22oi_1
X_21759_ _22016_/CLK _21759_/D vssd1 vssd1 vccd1 vccd1 _21759_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_54_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14300_ _14913_/A _14296_/B _14288_/A vssd1 vssd1 vccd1 vccd1 _14448_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_0_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11512_ _11511_/X _19382_/B _11521_/S vssd1 vssd1 vccd1 vccd1 _21842_/D sky130_fd_sc_hd__mux2_1
X_15280_ _15281_/A _15281_/B vssd1 vssd1 vccd1 vccd1 _15419_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_135_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12492_ _12497_/B _12492_/B vssd1 vssd1 vccd1 vccd1 _12493_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_81_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14231_ _14231_/A _14231_/B vssd1 vssd1 vccd1 vccd1 _14240_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14383__A1 _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11443_ _11442_/X hold264/X _11470_/S vssd1 vssd1 vccd1 vccd1 _21819_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_0_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15580__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14383__B2 _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14162_ _14162_/A _14162_/B _14162_/C vssd1 vssd1 vccd1 vccd1 _14162_/X sky130_fd_sc_hd__and3_1
XFILLER_0_1_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11374_ _11373_/X _16743_/C _11401_/S vssd1 vssd1 vccd1 vccd1 _21796_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_104_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17321__A1 _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13113_ _13975_/B _14312_/D _13858_/C _13402_/D vssd1 vssd1 vccd1 vccd1 _13113_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_132_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14093_ _14093_/A _14093_/B _14093_/C vssd1 vssd1 vccd1 vccd1 _14095_/B sky130_fd_sc_hd__nand3_1
X_18970_ _18969_/B _18969_/C _18969_/A vssd1 vssd1 vccd1 vccd1 _18972_/B sky130_fd_sc_hd__a21o_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14811__C _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21405__B1 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13044_ _14712_/A _14712_/B _14384_/C _14384_/D vssd1 vssd1 vccd1 vccd1 _13046_/A
+ sky130_fd_sc_hd__and4_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17921_ _17921_/A _17921_/B _17921_/C vssd1 vssd1 vccd1 vccd1 _17923_/A sky130_fd_sc_hd__and3_1
XANTENNA__19890__B _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18787__A _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17852_ _17852_/A _17852_/B _17852_/C vssd1 vssd1 vccd1 vccd1 _17853_/B sky130_fd_sc_hd__and3_1
XANTENNA__19812__A2_N _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16803_ _16868_/A _16917_/C _16968_/C _16734_/B vssd1 vssd1 vccd1 vccd1 _16803_/X
+ sky130_fd_sc_hd__a22o_1
X_17783_ _17913_/B _17781_/X _17666_/X _17669_/A vssd1 vssd1 vccd1 vccd1 _17784_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_156_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14995_ _15768_/A _16418_/A vssd1 vssd1 vccd1 vccd1 _14996_/B sky130_fd_sc_hd__and2_1
XFILLER_0_89_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13724__A _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19377__A2 _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19522_ _19522_/A _19522_/B vssd1 vssd1 vccd1 vccd1 _19524_/B sky130_fd_sc_hd__xnor2_1
X_16734_ _16868_/A _16734_/B _16860_/C _16917_/C vssd1 vssd1 vccd1 vccd1 _16734_/X
+ sky130_fd_sc_hd__and4_1
X_13946_ _13943_/X _13944_/X _13795_/C _13794_/Y vssd1 vssd1 vccd1 vccd1 _13948_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_88_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19453_ _19453_/A _19453_/B vssd1 vssd1 vccd1 vccd1 _19456_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_92_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16665_ _16665_/A _16665_/B _16665_/C vssd1 vssd1 vccd1 vccd1 _16669_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_53_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13877_ _13877_/A _16286_/A _13877_/C _14032_/A vssd1 vssd1 vccd1 vccd1 _14032_/B
+ sky130_fd_sc_hd__nand4_1
X_18404_ _18849_/B _19185_/D _19199_/C _19199_/D vssd1 vssd1 vccd1 vccd1 _18552_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_57_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15616_ _15473_/B _15475_/C _15614_/Y _15615_/X vssd1 vssd1 vccd1 vccd1 _15616_/Y
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__19411__A _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19384_ _19380_/X _19382_/Y _19226_/X _19229_/X vssd1 vssd1 vccd1 vccd1 _19385_/B
+ sky130_fd_sc_hd__a211o_1
X_12828_ fanout9/X _17599_/B vssd1 vssd1 vccd1 vccd1 _12828_/Y sky130_fd_sc_hd__nor2_1
X_16596_ _16597_/A _16597_/B vssd1 vssd1 vccd1 vccd1 _17217_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__12059__B _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18335_ _18787_/A _18787_/B _19546_/D _19906_/C vssd1 vssd1 vccd1 vccd1 _18481_/A
+ sky130_fd_sc_hd__and4_1
X_15547_ _15547_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15558_/A sky130_fd_sc_hd__or2_1
XANTENNA__11424__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ _12759_/A _12759_/B vssd1 vssd1 vccd1 vccd1 _12762_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_16_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18266_ _18267_/A _18267_/B vssd1 vssd1 vccd1 vccd1 _18266_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15478_ _15475_/Y _15476_/X _15295_/A _15341_/X vssd1 vssd1 vccd1 vccd1 _15478_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_114_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17217_ _17217_/A _17217_/B _17217_/C vssd1 vssd1 vccd1 vccd1 _17219_/C sky130_fd_sc_hd__nand3_1
XANTENNA__18468__A2_N _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15571__B1 _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14429_ _14430_/A _14430_/B vssd1 vssd1 vccd1 vccd1 _14429_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18197_ _19438_/A _19438_/B _19092_/C _19262_/C vssd1 vssd1 vccd1 vccd1 _18197_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_114_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17148_ _17150_/A _17150_/B _17149_/A _17149_/B vssd1 vssd1 vccd1 vccd1 _17148_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_141_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout8 fanout8/A vssd1 vssd1 vccd1 vccd1 fanout8/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__10935__A1 _10934_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17079_ _17078_/A _17077_/Y _17038_/X _17060_/Y vssd1 vssd1 vccd1 vccd1 _17081_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_110_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20090_ _20091_/B _20091_/A vssd1 vssd1 vccd1 vccd1 _20386_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_0_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19008__D _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11360__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout185_A _21825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17032__A2_N _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20992_ _20992_/A _21096_/B vssd1 vssd1 vccd1 vccd1 _20994_/B sky130_fd_sc_hd__or2_1
XANTENNA__14449__B _14449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15929__A2 _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout352_A _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21613_ _21906_/CLK _21613_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[76] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_36_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout617_A _21717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21544_ mstream_o[7] hold19/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22071_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_47_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17551__A1 _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21475_ hold166/X sstream_i[52] _21481_/S vssd1 vssd1 vccd1 vccd1 _22002_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20426_ _20616_/B _20426_/B vssd1 vssd1 vccd1 vccd1 _20441_/A sky130_fd_sc_hd__and2_1
XFILLER_0_132_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20357_ _20165_/Y _20211_/Y _20355_/Y _20356_/X vssd1 vssd1 vccd1 vccd1 _20357_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_101_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout98_A _21842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11090_ _11043_/X hold13/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21684_/D sky130_fd_sc_hd__mux2_1
XANTENNA__20930__A _21842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20288_ _20288_/A _20427_/B vssd1 vssd1 vccd1 vccd1 _20290_/B sky130_fd_sc_hd__or2_1
X_22027_ _22038_/CLK _22027_/D vssd1 vssd1 vccd1 vccd1 hold312/A sky130_fd_sc_hd__dfxtp_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18400__A _21791_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16814__B1 _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 hold75/A vssd1 vssd1 vccd1 vccd1 hold75/X sky130_fd_sc_hd__dlygate4sd3_1
X_13800_ _13800_/A _13800_/B _13800_/C _13800_/D vssd1 vssd1 vccd1 vccd1 _13800_/X
+ sky130_fd_sc_hd__or4_2
Xhold86 hold86/A vssd1 vssd1 vccd1 vccd1 hold86/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 hold97/A vssd1 vssd1 vccd1 vccd1 hold97/X sky130_fd_sc_hd__dlygate4sd3_1
X_14780_ _14780_/A _14780_/B vssd1 vssd1 vccd1 vccd1 _14782_/B sky130_fd_sc_hd__xnor2_1
X_11992_ _11992_/A _11992_/B vssd1 vssd1 vccd1 vccd1 _11994_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_39_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13731_ _13732_/A _13732_/B _13732_/C vssd1 vssd1 vccd1 vccd1 _13734_/B sky130_fd_sc_hd__a21o_1
X_10943_ hold263/A hold273/A vssd1 vssd1 vccd1 vccd1 _10945_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16450_ _16456_/A _16456_/B vssd1 vssd1 vccd1 vccd1 _16493_/A sky130_fd_sc_hd__nand2b_1
X_10874_ _10880_/B _10874_/B vssd1 vssd1 vccd1 vccd1 _10874_/Y sky130_fd_sc_hd__nor2_4
X_13662_ _13662_/A _13662_/B vssd1 vssd1 vccd1 vccd1 _13964_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__20377__A _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16593__A2 _16813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20690__A1_N _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15401_ _15402_/A _15402_/B vssd1 vssd1 vccd1 vccd1 _15600_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_38_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12613_ _12505_/A _12505_/B _12503_/A vssd1 vssd1 vccd1 vccd1 _12615_/B sky130_fd_sc_hd__o21ai_2
X_16381_ _16345_/A _16345_/B _16301_/A vssd1 vssd1 vccd1 vccd1 _16382_/B sky130_fd_sc_hd__a21oi_1
X_13593_ _15514_/B _14365_/D _14212_/C _15514_/A vssd1 vssd1 vccd1 vccd1 _13593_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_13_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18120_ _18120_/A _18120_/B vssd1 vssd1 vccd1 vccd1 _18122_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15332_ _15332_/A _15332_/B _15332_/C vssd1 vssd1 vccd1 vccd1 _15334_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_109_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12544_ _12544_/A _12544_/B _12544_/C vssd1 vssd1 vccd1 vccd1 _12544_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13710__C _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18051_ _18049_/Y _18185_/A _19692_/A _18789_/A vssd1 vssd1 vccd1 vccd1 _18185_/B
+ sky130_fd_sc_hd__and4bb_1
X_15263_ _16196_/B _16369_/A _15264_/C _15264_/D vssd1 vssd1 vccd1 vccd1 _15267_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_81_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12475_ _12475_/A _12475_/B _12475_/C _12475_/D vssd1 vssd1 vccd1 vccd1 _12475_/Y
+ sky130_fd_sc_hd__nor4_4
XFILLER_0_41_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17002_ _17002_/A _17002_/B _17002_/C vssd1 vssd1 vccd1 vccd1 _17002_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_35_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12326__C _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20429__A1 _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14214_ _14537_/A _14365_/D vssd1 vssd1 vccd1 vccd1 _14215_/B sky130_fd_sc_hd__and2_1
XFILLER_0_112_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12906__A2 _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20429__B2 _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11426_ _11447_/A1 hold296/A fanout48/X hold130/A vssd1 vssd1 vccd1 vccd1 _11426_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15194_ _15195_/A _15195_/B vssd1 vssd1 vccd1 vccd1 _15194_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_6 _11319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14145_ _14146_/A _14146_/B vssd1 vssd1 vccd1 vccd1 _14317_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_10_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11357_ _11124_/A hold224/X _11126_/B hold213/X vssd1 vssd1 vccd1 vccd1 _11357_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19109__C _19753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__A1 _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14076_ _14557_/B _14077_/B _14077_/C _14231_/A vssd1 vssd1 vccd1 vccd1 _14076_/X
+ sky130_fd_sc_hd__a22o_1
X_18953_ _18950_/X _19106_/B _18795_/X _18798_/A vssd1 vssd1 vccd1 vccd1 _18954_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ _12858_/C _11287_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21773_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_123_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11884__D _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12342__B _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ _13027_/A _13148_/B _13027_/C vssd1 vssd1 vccd1 vccd1 _13029_/B sky130_fd_sc_hd__nand3_4
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17904_ _17904_/A _17904_/B _17904_/C vssd1 vssd1 vccd1 vccd1 _18026_/A sky130_fd_sc_hd__nand3_1
X_18884_ _18881_/Y _18882_/Y _18719_/Y _18721_/Y vssd1 vssd1 vccd1 vccd1 _18885_/D
+ sky130_fd_sc_hd__a211oi_2
X_17835_ hold96/X fanout7/X _11553_/Y vssd1 vssd1 vccd1 vccd1 _17835_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19125__B _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17766_ _17765_/B _17765_/C _17765_/A vssd1 vssd1 vccd1 vccd1 _17768_/B sky130_fd_sc_hd__a21o_1
X_14978_ _15076_/B _16380_/B _16173_/B _15076_/A vssd1 vssd1 vccd1 vccd1 _14981_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19505_ _19664_/B _20671_/B _19372_/X _19373_/X fanout96/X vssd1 vssd1 vccd1 vccd1
+ _19510_/A sky130_fd_sc_hd__a32o_1
X_16717_ _16682_/X _16713_/Y _16711_/X _16708_/Y vssd1 vssd1 vccd1 vccd1 _16718_/C
+ sky130_fd_sc_hd__a211o_1
X_13929_ _13928_/B _13928_/C _13928_/A vssd1 vssd1 vccd1 vccd1 _13931_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_107_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17697_ _17693_/X _17695_/Y _17580_/C _17580_/Y vssd1 vssd1 vccd1 vccd1 _17698_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22073__RESET_B fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19436_ _19436_/A _19436_/B vssd1 vssd1 vccd1 vccd1 _19449_/A sky130_fd_sc_hd__xor2_4
XANTENNA__21390__B _21390_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16648_ _16648_/A _16648_/B _16648_/C vssd1 vssd1 vccd1 vccd1 _16653_/A sky130_fd_sc_hd__nand3_4
XFILLER_0_53_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17781__A1 _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19367_ _19368_/B _19368_/A vssd1 vssd1 vccd1 vccd1 _19483_/A sky130_fd_sc_hd__and2b_1
XANTENNA__21314__C1 _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16579_ _17211_/B _16578_/B _16578_/C vssd1 vssd1 vccd1 vccd1 _16580_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_45_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20668__A1 _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18318_ _19535_/A _18622_/B _19089_/B _18319_/B vssd1 vssd1 vccd1 vccd1 _18320_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20668__B2 _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13620__C _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19298_ _19299_/A _19299_/B vssd1 vssd1 vccd1 vccd1 _19298_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_5_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14347__A1 _14659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14347__B2 _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18249_ _18394_/A _18245_/B _18240_/X vssd1 vssd1 vccd1 vccd1 _18390_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_44_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17596__A _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12358__B1 _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21260_ _21260_/A _21260_/B vssd1 vssd1 vccd1 vccd1 _21266_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20211_ _20212_/A _20212_/B vssd1 vssd1 vccd1 vccd1 _20211_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_64_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13570__A2 _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21191_ _21191_/A _21191_/B vssd1 vssd1 vccd1 vccd1 _21193_/A sky130_fd_sc_hd__nor2_1
XANTENNA_fanout100_A _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12533__A _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20840__A1 _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20142_ _20142_/A _20142_/B vssd1 vssd1 vccd1 vccd1 _20157_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_0_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19589__A2 _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20073_ _20224_/A _20073_/B vssd1 vssd1 vccd1 vccd1 _20075_/B sky130_fd_sc_hd__and2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16037__B1_N _15907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11333__B2 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout567_A _12403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11097__A0 _11059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20975_ _20845_/D _21293_/B _21853_/Q _20975_/D vssd1 vssd1 vccd1 vccd1 _21095_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_135_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19051__A _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14195__A _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12427__B _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21527_ hold286/X sstream_i[104] _21528_/S vssd1 vssd1 vccd1 vccd1 _22054_/D sky130_fd_sc_hd__mux2_1
XANTENNA__21725__RESET_B _21329_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15535__B1 _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12260_ _12268_/A _12269_/C _12249_/C _12249_/D vssd1 vssd1 vccd1 vccd1 _12264_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21458_ hold196/X sstream_i[35] _21494_/S vssd1 vssd1 vccd1 vccd1 _21985_/D sky130_fd_sc_hd__mux2_1
X_11211_ hold214/X _11122_/X fanout48/X hold245/A vssd1 vssd1 vccd1 vccd1 _11211_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16560__D _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20409_ _20256_/A _20256_/B _20260_/B vssd1 vssd1 vccd1 vccd1 _20446_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_142_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12191_ _12191_/A _12191_/B vssd1 vssd1 vccd1 vccd1 _12193_/B sky130_fd_sc_hd__xnor2_1
X_21389_ hold174/X _21390_/B _21387_/Y _21388_/X vssd1 vssd1 vccd1 vccd1 _21937_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11572__A1 _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11142_ hold255/X _11126_/A fanout45/X hold186/X vssd1 vssd1 vccd1 vccd1 _11142_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13258__B _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12162__B _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15950_ _15784_/B _15823_/X _15948_/Y _15949_/X vssd1 vssd1 vccd1 vccd1 _15999_/A
+ sky130_fd_sc_hd__a211oi_4
X_11073_ _10886_/Y hold68/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21668_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19226__A _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11324__A1 _11323_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14901_ _14901_/A _14901_/B vssd1 vssd1 vccd1 vccd1 _14904_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__16569__B _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15881_ _15878_/Y _15879_/X _15743_/Y _15745_/Y vssd1 vssd1 vccd1 vccd1 _15881_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17620_ _17619_/A _21056_/A _17739_/D _17619_/B vssd1 vssd1 vccd1 vccd1 _17620_/Y
+ sky130_fd_sc_hd__a22oi_1
X_14832_ _14831_/B _15029_/B _14831_/A vssd1 vssd1 vccd1 vccd1 _14833_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13705__C _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14089__B hold313/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11088__A0 _10988_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17551_ _17915_/A _19587_/B _17915_/D _19587_/A vssd1 vssd1 vccd1 vccd1 _17551_/Y
+ sky130_fd_sc_hd__a22oi_1
X_14763_ _14627_/A _14627_/B _14630_/A vssd1 vssd1 vccd1 vccd1 _14906_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_86_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11975_ _11901_/X _11972_/Y _11982_/A _11971_/A vssd1 vssd1 vccd1 vccd1 _11976_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_58_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16502_ _16498_/X _16500_/Y _16471_/A _16474_/A vssd1 vssd1 vccd1 vccd1 _16503_/C
+ sky130_fd_sc_hd__a211oi_1
X_13714_ _13714_/A _13714_/B vssd1 vssd1 vccd1 vccd1 _13716_/B sky130_fd_sc_hd__or2_1
XANTENNA__19752__A2 _19753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10926_ _10926_/A _10926_/B vssd1 vssd1 vccd1 vccd1 _10926_/X sky130_fd_sc_hd__xor2_4
X_17482_ _17483_/A _17483_/B _17483_/C _17483_/D vssd1 vssd1 vccd1 vccd1 _17594_/A
+ sky130_fd_sc_hd__a31o_2
X_14694_ _16418_/A _14693_/X _14692_/X vssd1 vssd1 vccd1 vccd1 _14696_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_156_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19221_ _19373_/B _20462_/D _19221_/C vssd1 vssd1 vccd1 vccd1 _19221_/X sky130_fd_sc_hd__and3_1
XFILLER_0_67_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16433_ _16433_/A _16433_/B vssd1 vssd1 vccd1 vccd1 _16434_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13645_ _13491_/C _13490_/Y _13643_/X _13644_/Y vssd1 vssd1 vccd1 vccd1 _13648_/C
+ sky130_fd_sc_hd__o211a_2
X_10857_ _10857_/A _10857_/B vssd1 vssd1 vccd1 vccd1 _10859_/C sky130_fd_sc_hd__nand2_1
XANTENNA__19896__A _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18008__C _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19152_ _19152_/A _19152_/B _19152_/C vssd1 vssd1 vccd1 vccd1 _19154_/A sky130_fd_sc_hd__and3_1
X_16364_ _10984_/Y fanout5/X _16362_/Y _12291_/B _16363_/X vssd1 vssd1 vccd1 vccd1
+ _16364_/X sky130_fd_sc_hd__a221o_1
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13576_ _13732_/A _13576_/B vssd1 vssd1 vccd1 vccd1 _13578_/B sky130_fd_sc_hd__and2_1
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18103_ hold63/X fanout7/X _18101_/X _11547_/X _18102_/Y vssd1 vssd1 vccd1 vccd1
+ _18103_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_13_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11260__A0 _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15315_ _15315_/A _15315_/B vssd1 vssd1 vccd1 vccd1 _15334_/A sky130_fd_sc_hd__xnor2_1
X_19083_ _19083_/A _19083_/B vssd1 vssd1 vccd1 vccd1 _19143_/A sky130_fd_sc_hd__xor2_1
X_12527_ _12604_/A _12526_/C _12526_/A vssd1 vssd1 vccd1 vccd1 _12587_/B sky130_fd_sc_hd__o21a_1
X_16295_ _16372_/A _16295_/B vssd1 vssd1 vccd1 vccd1 _16297_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_14_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18034_ _21087_/D _18319_/B _18622_/B _20583_/A vssd1 vssd1 vccd1 vccd1 _18035_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15246_ _15246_/A vssd1 vssd1 vccd1 vccd1 _15246_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_140_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12458_ _12458_/A _12785_/B _13034_/D _14386_/B vssd1 vssd1 vccd1 vccd1 _12460_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_124_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16470__D _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11409_ hold281/A fanout28/X _11408_/X vssd1 vssd1 vccd1 vccd1 _11409_/X sky130_fd_sc_hd__a21o_1
X_15177_ _15177_/A _15177_/B _15177_/C vssd1 vssd1 vccd1 vccd1 _15179_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_50_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12389_ _11909_/B _12388_/B _11907_/A vssd1 vssd1 vccd1 vccd1 _12390_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__12353__A _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__A1 _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11563__B2 _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14128_ _12291_/B _14126_/X _14127_/X vssd1 vssd1 vccd1 vccd1 _14128_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_10_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19985_ _19983_/Y _20122_/B _19885_/B _19884_/Y vssd1 vssd1 vccd1 vccd1 _19985_/Y
+ sky130_fd_sc_hd__a211oi_1
X_14059_ _15373_/A _14873_/B _14217_/D _14859_/A vssd1 vssd1 vccd1 vccd1 _14062_/B
+ sky130_fd_sc_hd__a22o_1
X_18936_ _18936_/A _18936_/B _18936_/C vssd1 vssd1 vccd1 vccd1 _18938_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_20_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18867_ _18745_/A _18744_/B _18742_/X vssd1 vssd1 vccd1 vccd1 _18867_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17818_ _17815_/X _17816_/Y _17693_/C _17694_/X vssd1 vssd1 vccd1 vccd1 _17819_/C
+ sky130_fd_sc_hd__o211ai_2
X_18798_ _18798_/A _18798_/B vssd1 vssd1 vccd1 vccd1 _18807_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11079__A0 _10934_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17749_ _17749_/A _17749_/B _17749_/C vssd1 vssd1 vccd1 vccd1 _17750_/C sky130_fd_sc_hd__nand3_1
X_20760_ _20757_/X _20758_/Y _20623_/X _20627_/C vssd1 vssd1 vccd1 vccd1 _20760_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14017__B1 _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14727__B _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19419_ _19416_/Y _19417_/X _19264_/D _19266_/B vssd1 vssd1 vccd1 vccd1 _19420_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_134_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15765__B1 _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20691_ _20808_/A _21046_/B _21171_/A _20691_/D vssd1 vssd1 vccd1 vccd1 _20808_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_91_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12528__A _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout148_A _19092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11251__B1 _11250_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout315_A _21792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21312_ _21230_/A _21230_/B _21229_/A vssd1 vssd1 vccd1 vccd1 _21318_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_103_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13976__A1_N _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold320 hold320/A vssd1 vssd1 vccd1 vccd1 hold320/X sky130_fd_sc_hd__dlygate4sd3_1
X_21243_ _21243_/A _21243_/B vssd1 vssd1 vccd1 vccd1 _21244_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_13_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold331 hold331/A vssd1 vssd1 vccd1 vccd1 hold331/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14181__C _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21174_ _21174_/A _21174_/B vssd1 vssd1 vccd1 vccd1 _21175_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_1_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19691__D _19691_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20125_ _20125_/A _20125_/B vssd1 vssd1 vccd1 vccd1 _20161_/A sky130_fd_sc_hd__and2_1
XFILLER_0_110_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11306__A1 _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21369__A2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19431__A1 _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20056_ _20053_/X _20054_/Y _19828_/B _19830_/B vssd1 vssd1 vccd1 vccd1 _20056_/Y
+ sky130_fd_sc_hd__o211ai_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold262_A hold262/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13525__C _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16796__A2 _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_204 hold270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_215 hold275/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_226 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_237 hold309/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13822__A _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_248 hold262/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _11741_/A _11741_/C _11741_/B vssd1 vssd1 vccd1 vccd1 _11761_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_138_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_259 hold262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20958_ _20960_/B vssd1 vssd1 vccd1 vccd1 _20958_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_67_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14637__B _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11691_ _11691_/A _11691_/B vssd1 vssd1 vccd1 vccd1 _11699_/A sky130_fd_sc_hd__xnor2_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20889_ _20886_/X _20887_/Y _20750_/A _20753_/A vssd1 vssd1 vccd1 vccd1 _20889_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13430_ _13306_/B _13306_/Y _13428_/Y _13429_/X vssd1 vssd1 vccd1 vccd1 _13430_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_76_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20655__A _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19866__D _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13361_ _13361_/A _13512_/A _13361_/C vssd1 vssd1 vccd1 vccd1 _13363_/A sky130_fd_sc_hd__or3_1
XFILLER_0_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18170__A1 _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17667__C _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15100_ _15097_/X _15238_/B _14998_/X _15001_/X vssd1 vssd1 vccd1 vccd1 _15101_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__18170__B2 _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_774 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12312_ _12312_/A _13258_/C _12313_/A vssd1 vssd1 vccd1 vccd1 _12312_/X sky130_fd_sc_hd__and3_1
X_16080_ _16079_/B _16079_/C _16079_/A vssd1 vssd1 vccd1 vccd1 _16080_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_122_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13292_ _13292_/A _13292_/B vssd1 vssd1 vccd1 vccd1 _13302_/A sky130_fd_sc_hd__and2_1
XANTENNA__21057__A1 _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11488__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15031_ _15931_/B _16328_/A _16326_/A _15931_/A vssd1 vssd1 vccd1 vccd1 _15034_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13269__A _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12243_ _12226_/A _12226_/C _12226_/B vssd1 vssd1 vccd1 vccd1 _12256_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11545__A1 _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12174_ _12128_/B _12131_/Y _12169_/X _12172_/X vssd1 vssd1 vccd1 vccd1 _12174_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20390__A _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11125_ _11124_/A _11126_/A _11126_/B _21422_/A vssd1 vssd1 vccd1 vccd1 _11348_/S
+ sky130_fd_sc_hd__o31a_4
X_19770_ _19617_/A _19617_/B _19615_/X vssd1 vssd1 vccd1 vccd1 _19772_/B sky130_fd_sc_hd__a21oi_2
X_16982_ _16982_/A _16982_/B _16982_/C vssd1 vssd1 vccd1 vccd1 _16994_/A sky130_fd_sc_hd__and3_2
X_18721_ _18559_/A _18560_/Y _18719_/Y _18720_/X vssd1 vssd1 vccd1 vccd1 _18721_/Y
+ sky130_fd_sc_hd__a211oi_4
X_15933_ _16056_/A _16391_/B _15933_/C _15933_/D vssd1 vssd1 vccd1 vccd1 _16056_/B
+ sky130_fd_sc_hd__and4b_1
X_11056_ _11055_/Y hold65/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21657_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18652_ _18652_/A _19123_/B _19972_/C _21258_/B vssd1 vssd1 vccd1 vccd1 _18653_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__19973__A2 _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15864_ _15861_/Y _15862_/X _15721_/Y _15723_/Y vssd1 vssd1 vccd1 vccd1 _15864_/X
+ sky130_fd_sc_hd__o211a_1
X_17603_ _17825_/A _17603_/B vssd1 vssd1 vccd1 vccd1 _17698_/A sky130_fd_sc_hd__or2_1
X_14815_ _16196_/A _15791_/A _14817_/D _16374_/A vssd1 vssd1 vccd1 vccd1 _14820_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15931__B _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18583_ _19051_/A _19057_/C _19057_/D _20317_/D vssd1 vssd1 vccd1 vccd1 _18583_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_153_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15795_ _15795_/A _15921_/B vssd1 vssd1 vccd1 vccd1 _15798_/A sky130_fd_sc_hd__or2_1
XFILLER_0_87_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14828__A _16173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17534_ _17534_/A _17534_/B vssd1 vssd1 vccd1 vccd1 _17536_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14746_ _14746_/A _14746_/B vssd1 vssd1 vccd1 vccd1 _14747_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_8_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16539__A2 _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11958_ _11958_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _11960_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10909_ _10909_/A vssd1 vssd1 vccd1 vccd1 _10911_/C sky130_fd_sc_hd__inv_2
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17465_ _17466_/A _17466_/B _17466_/C _17466_/D vssd1 vssd1 vccd1 vccd1 _17465_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_156_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14677_ _14677_/A _14677_/B _14825_/B vssd1 vssd1 vccd1 vccd1 _14679_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_156_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11889_ _11889_/A _11889_/B _11889_/C vssd1 vssd1 vccd1 vccd1 _11889_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_104_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19204_ _19204_/A _19204_/B _19204_/C vssd1 vssd1 vccd1 vccd1 _19206_/B sky130_fd_sc_hd__nand3_1
X_16416_ _16416_/A _16416_/B vssd1 vssd1 vccd1 vccd1 _16422_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13628_ _13627_/B _13627_/C _13627_/A vssd1 vssd1 vccd1 vccd1 _13630_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_104_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20334__A2_N _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17396_ _17621_/C _17739_/C _17739_/D _17504_/C vssd1 vssd1 vccd1 vccd1 _17397_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19135_ _19135_/A _19135_/B _19135_/C vssd1 vssd1 vccd1 vccd1 _19135_/X sky130_fd_sc_hd__and3_1
X_16347_ _16347_/A _16347_/B _16347_/C vssd1 vssd1 vccd1 vccd1 _16349_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_137_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13559_ _13867_/A _13858_/A _14354_/C _14663_/D vssd1 vssd1 vccd1 vccd1 _13714_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_14_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18035__A _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12981__B1 _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19066_ _19087_/B _19089_/B _18928_/X _18929_/X _18773_/B vssd1 vssd1 vccd1 vccd1
+ _19071_/A sky130_fd_sc_hd__a32o_1
X_16278_ _16278_/A _16278_/B vssd1 vssd1 vccd1 vccd1 _16279_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_129_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21099__C _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11398__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18017_ _18018_/A _18018_/B _18018_/C vssd1 vssd1 vccd1 vccd1 _18017_/X sky130_fd_sc_hd__and3_1
X_15229_ _15892_/A _15632_/B _15370_/B _16391_/B vssd1 vssd1 vccd1 vccd1 _15407_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__17874__A _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11536__A1 _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18689__B _18689_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21396__A _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout107 _21267_/A vssd1 vssd1 vccd1 vccd1 _20797_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout118 _20562_/B vssd1 vssd1 vccd1 vccd1 _21169_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__17672__B1 _18789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout129 _20103_/A vssd1 vssd1 vccd1 vccd1 _18769_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_61_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19968_ _19874_/B _19967_/X _19966_/X vssd1 vssd1 vccd1 vccd1 _19970_/A sky130_fd_sc_hd__a21bo_1
X_18919_ _18919_/A _18919_/B _18919_/C vssd1 vssd1 vccd1 vccd1 _19049_/B sky130_fd_sc_hd__or3_1
XANTENNA__19413__A1 _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19413__B2 _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19899_ _19691_/X _19694_/X _19897_/X _19898_/Y vssd1 vssd1 vccd1 vccd1 _19899_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12530__B _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21930_ _21948_/CLK _21930_/D vssd1 vssd1 vccd1 vccd1 hold150/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14789__A1 _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21861_ _21932_/CLK hold108/X vssd1 vssd1 vccd1 vccd1 hold107/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout265_A _19531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20812_ _21056_/A _21169_/A _21256_/B hold264/A vssd1 vssd1 vccd1 vccd1 _20938_/A
+ sky130_fd_sc_hd__and4_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21792_ _21974_/CLK _21792_/D vssd1 vssd1 vccd1 vccd1 _21792_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__17727__A1 _21795_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14457__B _14774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17727__B2 _19337_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20178__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20743_ _20610_/Y _20612_/Y _20741_/Y _20742_/X vssd1 vssd1 vccd1 vccd1 _20743_/Y
+ sky130_fd_sc_hd__a211oi_2
XANTENNA_fanout432_A _21762_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20731__B1 _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19967__C _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14176__C _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18871__C _19053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20674_ _20797_/A _21258_/A _21153_/B _21264_/B vssd1 vssd1 vccd1 vccd1 _20801_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_135_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21039__A1 _21040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11527__A1 _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20922__B _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12724__B1 _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold150 hold150/A vssd1 vssd1 vccd1 vccd1 hold150/X sky130_fd_sc_hd__dlygate4sd3_1
X_21226_ _21226_/A _21226_/B vssd1 vssd1 vccd1 vccd1 _21228_/C sky130_fd_sc_hd__xnor2_2
Xhold161 hold161/A vssd1 vssd1 vccd1 vccd1 hold161/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 hold172/A vssd1 vssd1 vccd1 vccd1 hold172/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19652__B2 _19493_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold183 hold183/A vssd1 vssd1 vccd1 vccd1 hold183/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12143__D _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold194 hold194/A vssd1 vssd1 vccd1 vccd1 hold194/X sky130_fd_sc_hd__dlygate4sd3_1
X_21157_ _21258_/B _21156_/X _21155_/X vssd1 vssd1 vccd1 vccd1 _21159_/A sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout80_A _21847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout630 _21806_/Q vssd1 vssd1 vccd1 vccd1 _17657_/A sky130_fd_sc_hd__buf_8
XANTENNA__22105__RESET_B _11089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout641 _11041_/A vssd1 vssd1 vccd1 vccd1 fanout641/X sky130_fd_sc_hd__clkbuf_8
X_20108_ _20105_/Y _20251_/A _20249_/A _20242_/D vssd1 vssd1 vccd1 vccd1 _20251_/B
+ sky130_fd_sc_hd__and4bb_1
X_21088_ _21087_/D _21293_/B _21261_/B _20975_/D vssd1 vssd1 vccd1 vccd1 _21089_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__15454__D _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12930_ _12929_/B _12929_/C _12929_/A vssd1 vssd1 vccd1 vccd1 _12930_/Y sky130_fd_sc_hd__o21ai_2
X_20039_ _20039_/A _20039_/B vssd1 vssd1 vccd1 vccd1 _20041_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ _13554_/B _12402_/B _12989_/A _12860_/D vssd1 vssd1 vccd1 vccd1 _12862_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19223__B _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14600_ _14288_/A _14445_/A _14913_/C vssd1 vssd1 vccd1 vccd1 _14603_/B sky130_fd_sc_hd__a21oi_2
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ _11781_/A _11781_/C _11781_/B vssd1 vssd1 vccd1 vccd1 _11813_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_150_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15580_ _15435_/A _21788_/Q _16374_/B _15439_/D vssd1 vssd1 vccd1 vccd1 _15581_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ _12792_/A _12792_/B _12792_/C vssd1 vssd1 vccd1 vccd1 _12795_/A sky130_fd_sc_hd__nand3_2
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14367__B _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14531_ _14531_/A _14531_/B vssd1 vssd1 vccd1 vccd1 _14584_/A sky130_fd_sc_hd__xor2_4
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _11732_/A _11732_/C _11732_/B vssd1 vssd1 vccd1 vccd1 _11744_/C sky130_fd_sc_hd__a21o_1
XANTENNA__20722__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17250_ _17251_/A _17251_/B _17251_/C vssd1 vssd1 vccd1 vccd1 _17250_/X sky130_fd_sc_hd__and3_1
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14462_ _14462_/A _14462_/B vssd1 vssd1 vccd1 vccd1 _14467_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11674_ _12223_/A _12877_/B vssd1 vssd1 vccd1 vccd1 _11763_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_153_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16201_ _16201_/A _16201_/B vssd1 vssd1 vccd1 vccd1 _16202_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_36_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13413_ _13413_/A _13413_/B vssd1 vssd1 vccd1 vccd1 _13415_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17181_ _17490_/A _17282_/A _17739_/C _17739_/D vssd1 vssd1 vccd1 vccd1 _17183_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_3_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14393_ _14393_/A _14393_/B _14393_/C vssd1 vssd1 vccd1 vccd1 _14532_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16132_ _16132_/A _16132_/B vssd1 vssd1 vccd1 vccd1 _16134_/C sky130_fd_sc_hd__or2_1
XFILLER_0_109_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13344_ _13343_/A _13343_/B _13343_/C _13343_/D vssd1 vssd1 vccd1 vccd1 _13344_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_51_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18694__A2 _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16063_ _16171_/B vssd1 vssd1 vccd1 vccd1 _16064_/C sky130_fd_sc_hd__inv_2
X_13275_ _13275_/A _13427_/A _13275_/C vssd1 vssd1 vccd1 vccd1 _13427_/B sky130_fd_sc_hd__nand3_2
XANTENNA__11518__A1 _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15014_ _15010_/Y _15012_/X _14887_/B _14889_/A vssd1 vssd1 vccd1 vccd1 _15014_/Y
+ sky130_fd_sc_hd__a211oi_1
X_12226_ _12226_/A _12226_/B _12226_/C vssd1 vssd1 vccd1 vccd1 _12256_/A sky130_fd_sc_hd__and3_1
XFILLER_0_20_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19643__A1 _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19643__B2 _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14830__B _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12157_ _12157_/A _12197_/A vssd1 vssd1 vccd1 vccd1 _12160_/B sky130_fd_sc_hd__xor2_1
X_19822_ _19823_/A _20733_/C _20606_/D _20590_/D vssd1 vssd1 vccd1 vccd1 _19825_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19117__C _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11108_ _10903_/Y hold17/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21702_/D sky130_fd_sc_hd__mux2_1
XANTENNA__20270__D _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16965_ _16946_/A _16946_/C _16946_/B vssd1 vssd1 vccd1 vccd1 _16965_/Y sky130_fd_sc_hd__o21ai_1
X_12088_ _12261_/A _12269_/B _12639_/A _12530_/A vssd1 vssd1 vccd1 vccd1 _12091_/A
+ sky130_fd_sc_hd__nand4_2
X_19753_ _20650_/A _19753_/B _19753_/C _19753_/D vssd1 vssd1 vccd1 vccd1 _19753_/Y
+ sky130_fd_sc_hd__nand4_4
X_15916_ _16380_/A _15916_/B _16377_/B _16414_/B vssd1 vssd1 vccd1 vccd1 _16050_/A
+ sky130_fd_sc_hd__and4_1
X_11039_ mstream_o[113] hold283/X _11039_/S vssd1 vssd1 vccd1 vccd1 hold284/A sky130_fd_sc_hd__mux2_1
XANTENNA__19946__A2 _15070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18704_ _18705_/A _18705_/B vssd1 vssd1 vccd1 vccd1 _18866_/B sky130_fd_sc_hd__or2_1
XFILLER_0_95_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19414__A _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19684_ _19554_/A _19554_/B _19554_/C _19556_/X vssd1 vssd1 vccd1 vccd1 _19719_/A
+ sky130_fd_sc_hd__a31o_1
X_16896_ _16896_/A _16896_/B vssd1 vssd1 vccd1 vccd1 _16901_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18635_ _18787_/A _19732_/B _18640_/B _19092_/C _18487_/B vssd1 vssd1 vccd1 vccd1
+ _18644_/A sky130_fd_sc_hd__a41o_1
XANTENNA__15661__B _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15847_ _15847_/A _15847_/B vssd1 vssd1 vccd1 vccd1 _15867_/A sky130_fd_sc_hd__or2_1
XFILLER_0_91_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18566_ _18409_/A _18410_/Y _18563_/A _18564_/X vssd1 vssd1 vccd1 vccd1 _18566_/X
+ sky130_fd_sc_hd__a211o_1
X_15778_ _15778_/A _15778_/B vssd1 vssd1 vccd1 vccd1 _15780_/B sky130_fd_sc_hd__xor2_1
XTAP_3590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13181__B _14712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17517_ _17514_/A _17515_/Y _17426_/X _17429_/Y vssd1 vssd1 vccd1 vccd1 _17517_/Y
+ sky130_fd_sc_hd__o211ai_4
X_14729_ _15217_/A _15510_/B _14729_/C _14854_/A vssd1 vssd1 vccd1 vccd1 _14854_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_24_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13994__A2 _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18497_ _19445_/A _19874_/B vssd1 vssd1 vccd1 vccd1 _18500_/A sky130_fd_sc_hd__and2_1
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17448_ _17557_/A _17557_/B _17924_/B _17670_/B vssd1 vssd1 vccd1 vccd1 _17450_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_7_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17379_ _17379_/A _17379_/B _17479_/B vssd1 vssd1 vccd1 vccd1 _17483_/A sky130_fd_sc_hd__or3_1
XFILLER_0_43_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12954__B1 _11057_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19118_ _20242_/D _19117_/X _19116_/X vssd1 vssd1 vccd1 vccd1 _19120_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__11710__A _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20390_ _20910_/A _21278_/B _20390_/C _20559_/A vssd1 vssd1 vccd1 vccd1 _20559_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_42_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15499__A2 _21399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19049_ _18919_/B _19049_/B vssd1 vssd1 vccd1 vccd1 _19083_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_63_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11509__A1 _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_22060_ _22063_/CLK _22060_/D vssd1 vssd1 vccd1 vccd1 hold306/A sky130_fd_sc_hd__dfxtp_4
XFILLER_0_26_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21011_ _21008_/Y _21009_/X _20877_/B _20880_/B vssd1 vssd1 vccd1 vccd1 _21012_/C
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__16448__A1 _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout382_A _21773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15671__A2 _14698_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21913_ _21945_/CLK _21913_/D vssd1 vssd1 vccd1 vccd1 hold145/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11693__B1 _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21844_ _21845_/CLK _21844_/D vssd1 vssd1 vccd1 vccd1 _21844_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_78_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11604__B _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21775_ _21809_/CLK _21775_/D vssd1 vssd1 vccd1 vccd1 _21775_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_72_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19570__B1 _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15187__A1 _15046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20726_ _20726_/A _20726_/B vssd1 vssd1 vccd1 vccd1 _20728_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20657_ _20657_/A _20916_/A vssd1 vssd1 vccd1 vccd1 _20912_/A sky130_fd_sc_hd__or2_4
XFILLER_0_18_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11390_ _11124_/A hold250/X fanout45/X hold123/X vssd1 vssd1 vccd1 vccd1 _11390_/X
+ sky130_fd_sc_hd__a22o_1
X_20588_ _20588_/A _20588_/B vssd1 vssd1 vccd1 vccd1 _20589_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_33_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19873__A1 _21833_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13060_ _13059_/A _13059_/B _13059_/C vssd1 vssd1 vccd1 vccd1 _13062_/C sky130_fd_sc_hd__a21o_1
XANTENNA__18428__A2 _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16439__A1 _10988_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12011_ _12011_/A _12011_/B _12011_/C vssd1 vssd1 vccd1 vccd1 _12011_/Y sky130_fd_sc_hd__nand3_2
X_21209_ _21209_/A _21209_/B vssd1 vssd1 vccd1 vccd1 _21216_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13370__B1 _11063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17019__A _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15173__A2_N _15174_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout460 _16369_/B vssd1 vssd1 vccd1 vccd1 _14557_/D sky130_fd_sc_hd__buf_4
Xfanout471 _15091_/C vssd1 vssd1 vccd1 vccd1 _16266_/C sky130_fd_sc_hd__clkbuf_8
XANTENNA__15762__A _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout482 _21748_/Q vssd1 vssd1 vccd1 vccd1 _14391_/B sky130_fd_sc_hd__clkbuf_8
X_16750_ _16751_/A _16751_/B vssd1 vssd1 vccd1 vccd1 _16773_/A sky130_fd_sc_hd__nand2_1
Xfanout493 _21746_/Q vssd1 vssd1 vccd1 vccd1 _16409_/A sky130_fd_sc_hd__buf_4
X_13962_ _13962_/A _13962_/B vssd1 vssd1 vccd1 vccd1 _14291_/A sky130_fd_sc_hd__xor2_4
X_15701_ _15701_/A _15701_/B vssd1 vssd1 vccd1 vccd1 _15706_/A sky130_fd_sc_hd__xnor2_2
X_12913_ _12913_/A _12913_/B _12913_/C vssd1 vssd1 vccd1 vccd1 _12916_/A sky130_fd_sc_hd__nand3_1
X_16681_ _16682_/A _16682_/B _16682_/C vssd1 vssd1 vccd1 vccd1 _16681_/Y sky130_fd_sc_hd__nor3_1
X_13893_ _14365_/A _14384_/A _14212_/B vssd1 vssd1 vccd1 vccd1 _13893_/X sky130_fd_sc_hd__and3_1
XFILLER_0_115_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18420_ _18420_/A _18420_/B _18543_/A _18420_/D vssd1 vssd1 vccd1 vccd1 _18543_/B
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_154_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15632_ _15892_/A _15632_/B _16177_/B _16380_/B vssd1 vssd1 vccd1 vccd1 _15803_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ _12844_/A _12844_/B vssd1 vssd1 vccd1 vccd1 _12855_/A sky130_fd_sc_hd__or2_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18351_ _18498_/B _19874_/B _19872_/C _18652_/A vssd1 vssd1 vccd1 vccd1 _18352_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15563_ _15381_/Y _15386_/B _15561_/X _15562_/Y vssd1 vssd1 vccd1 vccd1 _15563_/Y
+ sky130_fd_sc_hd__a211oi_4
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12775_ _12669_/X _12672_/A _12896_/B _12774_/X vssd1 vssd1 vccd1 vccd1 _12775_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_96_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17302_ _17619_/A _17300_/C _17520_/D _17619_/B vssd1 vssd1 vccd1 vccd1 _17303_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14514_ _14385_/A _14387_/B _14385_/B vssd1 vssd1 vccd1 vccd1 _14519_/A sky130_fd_sc_hd__a21bo_1
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18282_ _18282_/A _18282_/B vssd1 vssd1 vccd1 vccd1 _18292_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11726_ _12458_/A _13173_/C _12357_/C _13155_/A vssd1 vssd1 vccd1 vccd1 _11727_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15494_ _15204_/A _15352_/Y _15492_/Y _15205_/X _15353_/X vssd1 vssd1 vccd1 vccd1
+ _15496_/C sky130_fd_sc_hd__a221oi_2
XFILLER_0_84_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17233_ _17334_/B _17666_/A _17443_/D _18166_/A vssd1 vssd1 vccd1 vccd1 _17235_/A
+ sky130_fd_sc_hd__a22oi_2
X_14445_ _14445_/A vssd1 vssd1 vccd1 vccd1 _14447_/A sky130_fd_sc_hd__inv_2
XANTENNA__16743__D _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11657_ _13012_/B _12268_/B _11649_/B _11648_/B vssd1 vssd1 vccd1 vccd1 _11664_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17164_ _16916_/Y _16961_/B _16961_/Y _17006_/Y _17163_/X vssd1 vssd1 vccd1 vccd1
+ _17164_/X sky130_fd_sc_hd__a32o_1
XANTENNA__20265__D _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14376_ _14375_/B _14375_/C _14375_/A vssd1 vssd1 vccd1 vccd1 _14376_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12400__A2 _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11588_ _11588_/A vssd1 vssd1 vccd1 vccd1 _11589_/D sky130_fd_sc_hd__inv_2
XFILLER_0_12_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16115_ _15980_/Y _15982_/Y _16113_/Y _16114_/X vssd1 vssd1 vccd1 vccd1 _16115_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_80_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13327_ _13327_/A _13327_/B _13327_/C vssd1 vssd1 vccd1 vccd1 _13330_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_12_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20474__A2 _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17095_ _17096_/A _17146_/D vssd1 vssd1 vccd1 vccd1 _17097_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_40_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19409__A _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18313__A _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20562__B _20562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16046_ _16165_/A vssd1 vssd1 vccd1 vccd1 _16048_/D sky130_fd_sc_hd__inv_2
XFILLER_0_126_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13258_ _13858_/B _13860_/A _13258_/C _13258_/D vssd1 vssd1 vccd1 vccd1 _13411_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_23_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12209_ _12168_/X _12176_/Y _12207_/B _12206_/Y vssd1 vssd1 vccd1 vccd1 _12209_/X
+ sky130_fd_sc_hd__a211o_1
X_13189_ _13188_/B _13188_/C _13188_/A vssd1 vssd1 vccd1 vccd1 _13191_/B sky130_fd_sc_hd__a21o_1
XANTENNA__20319__A1_N _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19805_ _19647_/A _19647_/B _19645_/B vssd1 vssd1 vccd1 vccd1 _19808_/C sky130_fd_sc_hd__o21ai_1
X_17997_ _19487_/B _18873_/A _19227_/C _19227_/D vssd1 vssd1 vccd1 vccd1 _17999_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__16768__A _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16948_ _16946_/A _16945_/Y _16947_/X _16890_/Y vssd1 vssd1 vccd1 vccd1 _16956_/A
+ sky130_fd_sc_hd__o211ai_4
X_19736_ _19735_/B _19849_/B _19735_/A vssd1 vssd1 vccd1 vccd1 _19737_/C sky130_fd_sc_hd__a21o_1
XANTENNA__16487__B _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16879_ _16816_/B _16879_/B vssd1 vssd1 vccd1 vccd1 _16881_/B sky130_fd_sc_hd__and2b_1
X_19667_ _19667_/A _19667_/B _19820_/B vssd1 vssd1 vccd1 vccd1 _19669_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_56_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18618_ _18618_/A _18618_/B vssd1 vssd1 vccd1 vccd1 _18620_/A sky130_fd_sc_hd__nand2_1
X_19598_ _19598_/A _19598_/B vssd1 vssd1 vccd1 vccd1 _19606_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17599__A _19636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18549_ _18550_/A _18550_/B vssd1 vssd1 vccd1 vccd1 _18707_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_47_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21560_ mstream_o[23] hold54/X _21562_/S vssd1 vssd1 vccd1 vccd1 _22087_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_74_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20511_ _20509_/Y _20511_/B vssd1 vssd1 vccd1 vccd1 _20643_/B sky130_fd_sc_hd__and2b_2
XFILLER_0_144_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21491_ hold165/X sstream_i[68] _21494_/S vssd1 vssd1 vccd1 vccd1 _22018_/D sky130_fd_sc_hd__mux2_1
XANTENNA_fanout228_A _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20442_ _20444_/A vssd1 vssd1 vccd1 vccd1 _20442_/Y sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_41_clk_i _21822_/CLK vssd1 vssd1 vccd1 vccd1 _21829_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20373_ _20079_/A _20224_/X _20372_/X _20080_/X _20226_/B vssd1 vssd1 vccd1 vccd1
+ _20373_/X sky130_fd_sc_hd__o221a_1
XFILLER_0_113_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout597_A _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20191__C _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22043_ _22049_/CLK _22043_/D vssd1 vssd1 vccd1 vccd1 hold236/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18596__C _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13407__A1 _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13407__B2 _21734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ _10890_/A _10899_/A vssd1 vssd1 vccd1 vccd1 _10892_/A sky130_fd_sc_hd__or2_2
XFILLER_0_156_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21827_ _21829_/CLK _21827_/D vssd1 vssd1 vccd1 vccd1 _21827_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_78_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12560_ _13173_/C _13155_/A _12780_/A _12780_/B vssd1 vssd1 vccd1 vccd1 _12562_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_93_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21758_ _22016_/CLK _21758_/D vssd1 vssd1 vccd1 vccd1 _21758_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11511_ _11224_/A t2x[20] v1z[20] fanout21/X _11510_/X vssd1 vssd1 vccd1 vccd1 _11511_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20709_ _20836_/B _20708_/C _20708_/A vssd1 vssd1 vccd1 vccd1 _20710_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12491_ _12496_/B _12388_/Y _12497_/A _12391_/A vssd1 vssd1 vccd1 vccd1 _12492_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_0_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21689_ _22080_/CLK _21689_/D vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14230_ _14230_/A _14230_/B vssd1 vssd1 vccd1 vccd1 _14264_/A sky130_fd_sc_hd__and2_1
XFILLER_0_18_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14383__A2 _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11442_ hold236/A fanout28/X _11441_/X vssd1 vssd1 vccd1 vccd1 _11442_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_34_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15580__B2 _15439_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14161_ _14160_/B _14160_/C _14160_/A vssd1 vssd1 vccd1 vccd1 _14162_/C sky130_fd_sc_hd__a21o_1
XANTENNA__19229__A _19230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11373_ hold179/X fanout29/X _11372_/X vssd1 vssd1 vccd1 vccd1 _11373_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18133__A _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17321__A2 _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13112_ _13112_/A _13112_/B vssd1 vssd1 vccd1 vccd1 _13213_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14092_ _13928_/A _13928_/B _13928_/C vssd1 vssd1 vccd1 vccd1 _14093_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21405__A1 _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13043_ _14716_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _13047_/A sky130_fd_sc_hd__nand2_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17920_ _18047_/B _17919_/C _17919_/A vssd1 vssd1 vccd1 vccd1 _17921_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12181__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13894__A1 _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19890__C _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15159__A_N _21733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18787__B _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17851_ _17852_/A _17852_/B _17852_/C vssd1 vssd1 vccd1 vccd1 _18095_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_79_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16802_ _16870_/A _17013_/C vssd1 vssd1 vccd1 vccd1 _16805_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_156_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17782_ _17666_/X _17669_/A _17913_/B _17781_/X vssd1 vssd1 vccd1 vccd1 _17782_/X
+ sky130_fd_sc_hd__o211a_1
X_14994_ _14994_/A _14994_/B vssd1 vssd1 vccd1 vccd1 _14996_/A sky130_fd_sc_hd__nand2_1
Xfanout290 _17874_/A vssd1 vssd1 vccd1 vccd1 _19487_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16733_ _16868_/A _17129_/B _16917_/C vssd1 vssd1 vccd1 vccd1 _16733_/X sky130_fd_sc_hd__and3_1
XANTENNA__18034__B1 _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19521_ _19521_/A _19521_/B vssd1 vssd1 vccd1 vccd1 _19522_/B sky130_fd_sc_hd__xnor2_1
X_13945_ _13795_/C _13794_/Y _13943_/X _13944_/X vssd1 vssd1 vccd1 vccd1 _13948_/C
+ sky130_fd_sc_hd__o211a_2
XANTENNA__13724__B _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19452_ _19452_/A _19452_/B vssd1 vssd1 vccd1 vccd1 _19453_/B sky130_fd_sc_hd__xnor2_4
X_16664_ _16639_/A _16639_/C _16639_/B vssd1 vssd1 vccd1 vccd1 _16665_/C sky130_fd_sc_hd__a21o_1
X_13876_ _13877_/A _16286_/A _13877_/C _14032_/A vssd1 vssd1 vccd1 vccd1 _13878_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20392__A1 _20249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20838__A _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15615_ _15612_/Y _15613_/X _15475_/A _15475_/Y vssd1 vssd1 vccd1 vccd1 _15615_/X
+ sky130_fd_sc_hd__o211a_1
X_18403_ _18849_/B _19199_/C _19199_/D _19185_/D vssd1 vssd1 vccd1 vccd1 _18403_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_147_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19383_ _19226_/X _19229_/X _19380_/X _19382_/Y vssd1 vssd1 vccd1 vccd1 _19383_/X
+ sky130_fd_sc_hd__o211a_1
X_12827_ _12827_/A _12827_/B vssd1 vssd1 vccd1 vccd1 _17599_/B sky130_fd_sc_hd__xnor2_4
X_16595_ _16595_/A _16595_/B vssd1 vssd1 vccd1 vccd1 _16597_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_69_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18337__A1 _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18334_ _18787_/B _19546_/D _19906_/C _18787_/A vssd1 vssd1 vccd1 vccd1 _18338_/C
+ sky130_fd_sc_hd__a22o_1
X_15546_ _15727_/B _15546_/B vssd1 vssd1 vccd1 vccd1 _15561_/A sky130_fd_sc_hd__and2_1
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12758_ _13155_/C _12756_/X _12757_/X vssd1 vssd1 vccd1 vccd1 _12759_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_29_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21341__B1 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18265_ _18265_/A _18265_/B vssd1 vssd1 vccd1 vccd1 _18267_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_38_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11709_ _11709_/A _11747_/A vssd1 vssd1 vccd1 vccd1 _11716_/A sky130_fd_sc_hd__nor2_1
X_15477_ _15295_/A _15341_/X _15475_/Y _15476_/X vssd1 vssd1 vccd1 vccd1 _15477_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_84_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15020__B1 _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12356__A _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12689_ _12578_/B _12578_/Y _12686_/X _12688_/Y vssd1 vssd1 vccd1 vccd1 _12692_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_154_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17216_ _17217_/A _17217_/B _17217_/C vssd1 vssd1 vccd1 vccd1 _17297_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_142_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14428_ _14264_/A _14264_/C _14264_/B vssd1 vssd1 vccd1 vccd1 _14430_/B sky130_fd_sc_hd__a21bo_2
XFILLER_0_115_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15571__A1 _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18196_ _19723_/A _18640_/B vssd1 vssd1 vccd1 vccd1 _18200_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17147_ _17089_/B _17145_/X _17146_/X vssd1 vssd1 vccd1 vccd1 _17150_/B sky130_fd_sc_hd__a21bo_1
X_14359_ _14355_/X _14357_/Y _14181_/X _14184_/X vssd1 vssd1 vccd1 vccd1 _14360_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout9 fanout9/A vssd1 vssd1 vccd1 vccd1 fanout9/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15386__B _15386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17078_ _17078_/A _17078_/B _17078_/C vssd1 vssd1 vccd1 vccd1 _17078_/X sky130_fd_sc_hd__or3_1
XFILLER_0_12_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16029_ _16029_/A _16029_/B vssd1 vssd1 vccd1 vccd1 _16031_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_126_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _21822_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_110_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13915__A _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19719_ _19719_/A _19719_/B _19719_/C vssd1 vssd1 vccd1 vccd1 _19721_/A sky130_fd_sc_hd__and3_1
X_20991_ _21096_/A _21311_/B _20991_/C _20991_/D vssd1 vssd1 vccd1 vccd1 _21096_/B
+ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout178_A _17443_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21612_ _21906_/CLK _21612_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[75] sky130_fd_sc_hd__dfrtp_4
XANTENNA__20135__A1 _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21332__B1 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21543_ mstream_o[6] hold16/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22070_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout512_A _21741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19491__A1_N _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21474_ hold142/X sstream_i[51] _21481_/S vssd1 vssd1 vccd1 vccd1 _22001_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_121_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20425_ _20425_/A _20425_/B vssd1 vssd1 vccd1 vccd1 _20426_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_132_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20356_ _20355_/C _20355_/B _20354_/Y vssd1 vssd1 vccd1 vccd1 _20356_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20287_ _20427_/A _21305_/A _21171_/A _20287_/D vssd1 vssd1 vccd1 vccd1 _20427_/B
+ sky130_fd_sc_hd__and4b_1
XANTENNA__13876__A1 _13877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20930__B _21815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22026_ _22038_/CLK _22026_/D vssd1 vssd1 vccd1 vccd1 hold303/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18400__B _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16814__A1 _16813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__21776__CLK _21822_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16814__B2 _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 hold76/A vssd1 vssd1 vccd1 vccd1 hold76/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 hold87/A vssd1 vssd1 vccd1 vccd1 hold87/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold98 hold98/A vssd1 vssd1 vccd1 vccd1 hold98/X sky130_fd_sc_hd__dlygate4sd3_1
X_11991_ _12094_/A _12094_/B _12639_/A _12530_/A vssd1 vssd1 vccd1 vccd1 _11992_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_98_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13730_ _13732_/A _13732_/B _13732_/C vssd1 vssd1 vccd1 vccd1 _13730_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10942_ mstream_o[55] _10941_/X _10992_/S vssd1 vssd1 vccd1 vccd1 _21592_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_129_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13661_ _13662_/A _13662_/B vssd1 vssd1 vccd1 vccd1 _13668_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_85_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10873_ _10873_/A _10873_/B _10873_/C vssd1 vssd1 vccd1 vccd1 _10874_/B sky130_fd_sc_hd__and3_1
XFILLER_0_97_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15400_ _15400_/A _15400_/B vssd1 vssd1 vccd1 vccd1 _15402_/B sky130_fd_sc_hd__or2_1
XFILLER_0_94_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12612_ _12728_/B _12612_/B vssd1 vssd1 vccd1 vccd1 _12615_/A sky130_fd_sc_hd__or2_1
X_16380_ _16380_/A _16380_/B vssd1 vssd1 vccd1 vccd1 _16382_/A sky130_fd_sc_hd__nand2_1
X_13592_ _13592_/A _13592_/B vssd1 vssd1 vccd1 vccd1 _13602_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15331_ _15179_/X _15331_/B vssd1 vssd1 vccd1 vccd1 _15332_/C sky130_fd_sc_hd__and2b_1
XFILLER_0_38_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17967__A _17967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12543_ _12544_/A _12544_/B _12544_/C vssd1 vssd1 vccd1 vccd1 _12543_/X sky130_fd_sc_hd__a21o_4
XFILLER_0_136_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13710__D _14663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18050_ _18787_/A _18787_/B _19089_/B _18773_/B vssd1 vssd1 vccd1 vccd1 _18185_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__12607__C _21776_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15262_ _15400_/A vssd1 vssd1 vccd1 vccd1 _15264_/D sky130_fd_sc_hd__inv_2
XFILLER_0_124_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12474_ _12470_/X _12472_/Y _12370_/B _12370_/Y vssd1 vssd1 vccd1 vccd1 _12475_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__20393__A _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17001_ _16946_/X _16965_/Y _16994_/A _16994_/Y vssd1 vssd1 vccd1 vccd1 _17002_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_124_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14213_ _14213_/A _14213_/B vssd1 vssd1 vccd1 vccd1 _14215_/A sky130_fd_sc_hd__nand2_1
XANTENNA__20429__A2 _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11425_ _11424_/X _21040_/A _11470_/S vssd1 vssd1 vccd1 vccd1 _21813_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_22_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12326__D _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14391__A _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15193_ _15056_/A _15056_/B _15054_/Y vssd1 vssd1 vccd1 vccd1 _15195_/B sky130_fd_sc_hd__a21boi_2
XANTENNA_7 _11319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14144_ _14144_/A _14144_/B vssd1 vssd1 vccd1 vccd1 _14146_/B sky130_fd_sc_hd__xor2_1
X_11356_ _11355_/X _17146_/D _11401_/S vssd1 vssd1 vccd1 vccd1 _21790_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_50_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19109__D _19751_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11590__A2 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14075_ _14848_/A _14557_/A _14234_/C _15001_/B vssd1 vssd1 vccd1 vccd1 _14231_/A
+ sky130_fd_sc_hd__nand4_2
X_18952_ _18795_/X _18798_/A _18950_/X _19106_/B vssd1 vssd1 vccd1 vccd1 _18952_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11287_ fanout58/X v0z[15] fanout17/X _11286_/X vssd1 vssd1 vccd1 vccd1 _11287_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ _13148_/A _13025_/C _13025_/A vssd1 vssd1 vccd1 vccd1 _13027_/C sky130_fd_sc_hd__a21o_1
XANTENNA__18255__B1 _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17903_ _17765_/A _17765_/C _17765_/B vssd1 vssd1 vccd1 vccd1 _17904_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18883_ _18719_/Y _18721_/Y _18881_/Y _18882_/Y vssd1 vssd1 vccd1 vccd1 _19006_/A
+ sky130_fd_sc_hd__o211a_1
X_17834_ _19636_/A _17834_/B vssd1 vssd1 vccd1 vccd1 _17834_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17207__A _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14977_ _14716_/A _14848_/C _14712_/X vssd1 vssd1 vccd1 vccd1 _15218_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_88_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17765_ _17765_/A _17765_/B _17765_/C vssd1 vssd1 vccd1 vccd1 _17768_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_89_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19504_ _19504_/A _19504_/B vssd1 vssd1 vccd1 vccd1 _19512_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13928_ _13928_/A _13928_/B _13928_/C vssd1 vssd1 vccd1 vccd1 _13931_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_77_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16716_ _16721_/A _16716_/B vssd1 vssd1 vccd1 vccd1 _16718_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_57_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13173__C _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17696_ _17580_/C _17580_/Y _17693_/X _17695_/Y vssd1 vssd1 vccd1 vccd1 _17698_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_88_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16647_ _16629_/A _16629_/B _16629_/C vssd1 vssd1 vccd1 vccd1 _16648_/C sky130_fd_sc_hd__a21o_1
X_19435_ _19433_/X _19435_/B vssd1 vssd1 vccd1 vccd1 _19436_/B sky130_fd_sc_hd__and2b_1
XANTENNA__10853__A1 _10852_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13859_ _13859_/A _13859_/B vssd1 vssd1 vccd1 vccd1 _13861_/A sky130_fd_sc_hd__nor2_1
XANTENNA__14566__A _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17781__A2 _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20287__B _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16578_ _17211_/B _16578_/B _16578_/C vssd1 vssd1 vccd1 vccd1 _17199_/A sky130_fd_sc_hd__nand3_1
X_19366_ _19366_/A _19366_/B vssd1 vssd1 vccd1 vccd1 _19368_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15529_ _15529_/A _15529_/B vssd1 vssd1 vccd1 vccd1 _15567_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20668__A2 _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18317_ _19695_/A _18624_/A vssd1 vssd1 vccd1 vccd1 _18321_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19297_ _19135_/A _19135_/C _19135_/B vssd1 vssd1 vccd1 vccd1 _19299_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__13620__D _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21399__A _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18248_ hold122/X _18247_/Y fanout2/X vssd1 vssd1 vccd1 vccd1 _21895_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_4_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14347__A2 _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17596__B _21343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12358__A1 _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18179_ _18179_/A _18179_/B vssd1 vssd1 vccd1 vccd1 _18181_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19286__A2 _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20210_ _20210_/A _20210_/B vssd1 vssd1 vccd1 vccd1 _20212_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11030__A1 hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21190_ _21291_/A _21296_/A _21286_/B _21296_/B vssd1 vssd1 vccd1 vccd1 _21191_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_12_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18494__B1 _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12533__B _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20141_ _20142_/A _20142_/B vssd1 vssd1 vccd1 vccd1 _20343_/B sky130_fd_sc_hd__or2_1
XFILLER_0_99_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18246__B1 _13369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20072_ _20072_/A _20072_/B _20072_/C vssd1 vssd1 vccd1 vccd1 _20073_/B sky130_fd_sc_hd__nand3_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout295_A _21796_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16659__C _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout462_A _21754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20974_ _20974_/A _21091_/A vssd1 vssd1 vccd1 vccd1 _20978_/A sky130_fd_sc_hd__or2_1
XANTENNA__17221__A1 _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19051__B _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15783__A1 _15907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14195__B _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12427__C _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15535__A1 _15916_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21526_ hold309/X sstream_i[103] _21528_/S vssd1 vssd1 vccd1 vccd1 _22053_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_8_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_133_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21102__A _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19277__A2 _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21457_ hold209/X sstream_i[34] _21489_/S vssd1 vssd1 vccd1 vccd1 _21984_/D sky130_fd_sc_hd__mux2_1
X_11210_ _15098_/B _11209_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21753_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12190_ _12223_/A _12269_/C _12191_/A vssd1 vssd1 vccd1 vccd1 _12199_/B sky130_fd_sc_hd__and3_1
X_20408_ _20408_/A _20408_/B vssd1 vssd1 vccd1 vccd1 _20450_/A sky130_fd_sc_hd__nand2_1
X_21388_ _21420_/S _14918_/Y _21403_/S vssd1 vssd1 vccd1 vccd1 _21388_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_32_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20941__A _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15299__B1 _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12443__B _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11572__A2 _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11141_ _12214_/C _11140_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21730_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19029__A2 _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19507__A _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20339_ _20340_/A _20340_/B vssd1 vssd1 vccd1 vccd1 _20339_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13258__C _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11072_ _10881_/X hold24/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21667_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18788__A1 _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14900_ _14900_/A _14900_/B vssd1 vssd1 vccd1 vccd1 _14901_/B sky130_fd_sc_hd__xnor2_1
X_22009_ _22013_/CLK _22009_/D vssd1 vssd1 vccd1 vccd1 hold161/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__16569__C _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15880_ _15743_/Y _15745_/Y _15878_/Y _15879_/X vssd1 vssd1 vccd1 vccd1 _16011_/A
+ sky130_fd_sc_hd__a211oi_4
X_14831_ _14831_/A _14831_/B _15029_/B vssd1 vssd1 vccd1 vccd1 _14833_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13705__D _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14089__C hold319/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17550_ _17550_/A _17550_/B vssd1 vssd1 vccd1 vccd1 _17570_/A sky130_fd_sc_hd__xor2_2
X_14762_ hold83/X _14761_/X fanout4/A vssd1 vssd1 vccd1 vccd1 hold84/A sky130_fd_sc_hd__mux2_1
X_11974_ _11901_/X _11972_/Y _11982_/A _11971_/A vssd1 vssd1 vccd1 vccd1 _11977_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__20388__A _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16501_ _16471_/A _16474_/A _16498_/X _16500_/Y vssd1 vssd1 vccd1 vccd1 _17197_/A
+ sky130_fd_sc_hd__o211a_2
X_13713_ _13713_/A _13713_/B vssd1 vssd1 vccd1 vccd1 _13716_/A sky130_fd_sc_hd__nor2_1
X_10925_ _10924_/A _10924_/B _10926_/A vssd1 vssd1 vccd1 vccd1 _10925_/Y sky130_fd_sc_hd__o21bai_1
X_17481_ _17593_/A _17481_/B vssd1 vssd1 vccd1 vccd1 _17483_/D sky130_fd_sc_hd__xor2_1
X_14693_ _15892_/A _15632_/B _16326_/A vssd1 vssd1 vccd1 vccd1 _14693_/X sky130_fd_sc_hd__and3_1
XANTENNA__14386__A _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13290__A _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16432_ _16432_/A _16432_/B vssd1 vssd1 vccd1 vccd1 _16433_/B sky130_fd_sc_hd__xnor2_1
X_19220_ _19373_/B _18732_/C _19221_/C _20462_/D vssd1 vssd1 vccd1 vccd1 _19220_/X
+ sky130_fd_sc_hd__a22o_1
X_13644_ _13643_/A _13643_/B _13643_/C _13643_/D vssd1 vssd1 vccd1 vccd1 _13644_/Y
+ sky130_fd_sc_hd__o22ai_4
X_10856_ _10857_/B vssd1 vssd1 vccd1 vccd1 _10866_/A sky130_fd_sc_hd__inv_2
XANTENNA__19896__B _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19151_ _19148_/X _19149_/Y _18985_/Y _18987_/X vssd1 vssd1 vccd1 vccd1 _19152_/C
+ sky130_fd_sc_hd__o211ai_2
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16363_ _16363_/A hold195/A vssd1 vssd1 vccd1 vccd1 _16363_/X sky130_fd_sc_hd__and2_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ _13572_/X _13720_/B _13437_/D _13439_/A vssd1 vssd1 vccd1 vccd1 _13576_/B
+ sky130_fd_sc_hd__o211ai_1
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18008__D _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18102_ _19636_/A _21355_/B vssd1 vssd1 vccd1 vccd1 _18102_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_27_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18712__A1 _19337_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15314_ _15314_/A _15314_/B vssd1 vssd1 vccd1 vccd1 _15315_/B sky130_fd_sc_hd__xnor2_1
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19082_ _19082_/A _19082_/B vssd1 vssd1 vccd1 vccd1 _19083_/B sky130_fd_sc_hd__nand2_1
X_12526_ _12526_/A _12604_/A _12526_/C vssd1 vssd1 vccd1 vccd1 _12604_/B sky130_fd_sc_hd__nor3_1
X_16294_ _16294_/A _16294_/B vssd1 vssd1 vccd1 vccd1 _16295_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_125_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18405__A2_N _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18033_ _21087_/D _19379_/B _18319_/B _18622_/B vssd1 vssd1 vccd1 vccd1 _18175_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15245_ _15247_/B _15247_/A vssd1 vssd1 vccd1 vccd1 _15246_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_125_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12457_ _13173_/C _12784_/A vssd1 vssd1 vccd1 vccd1 _12460_/A sky130_fd_sc_hd__and2_1
XFILLER_0_124_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11408_ _11447_/A1 hold295/A fanout47/X hold162/A vssd1 vssd1 vccd1 vccd1 _11408_/X
+ sky130_fd_sc_hd__a22o_1
X_15176_ _15175_/B _15316_/B _15175_/A vssd1 vssd1 vccd1 vccd1 _15177_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12388_ _12035_/A _12388_/B vssd1 vssd1 vccd1 vccd1 _12388_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__12353__B _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11563__A2 _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20283__B1 _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__A1 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14127_ _16363_/A hold191/A _10874_/Y fanout5/X vssd1 vssd1 vccd1 vccd1 _14127_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11339_ _21407_/S v0z[28] fanout20/X _11338_/X vssd1 vssd1 vccd1 vccd1 _11339_/X
+ sky130_fd_sc_hd__a31o_2
XANTENNA__19417__A _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19984_ _19984_/A _19984_/B _20126_/B _19984_/D vssd1 vssd1 vccd1 vccd1 _20122_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_120_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14058_ _15373_/B _14218_/B vssd1 vssd1 vccd1 vccd1 _14062_/A sky130_fd_sc_hd__and2_1
X_18935_ _18936_/B _18936_/C _18936_/A vssd1 vssd1 vccd1 vccd1 _18938_/A sky130_fd_sc_hd__a21o_1
X_13009_ _13097_/B _13009_/B vssd1 vssd1 vccd1 vccd1 _13072_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16479__C _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18866_ _18866_/A _18866_/B _18866_/C vssd1 vssd1 vccd1 vccd1 _18885_/B sky130_fd_sc_hd__and3_1
XFILLER_0_27_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17817_ _17693_/C _17694_/X _17815_/X _17816_/Y vssd1 vssd1 vccd1 vccd1 _17819_/B
+ sky130_fd_sc_hd__a211o_2
X_18797_ _19723_/A _19753_/B _18794_/Y _18795_/X vssd1 vssd1 vccd1 vccd1 _18798_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_94_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21535__A0 hold277/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17748_ _17749_/A _17749_/B _17749_/C vssd1 vssd1 vccd1 vccd1 _17750_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_89_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14017__A1 _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14017__B2 _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17679_ _17678_/B _17678_/C _17678_/A vssd1 vssd1 vccd1 vccd1 _17681_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_76_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19418_ _19264_/D _19266_/B _19416_/Y _19417_/X vssd1 vssd1 vccd1 vccd1 _19563_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15765__A1 _15892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20690_ _21171_/A _21046_/B _20688_/Y _20808_/A vssd1 vssd1 vccd1 vccd1 _20692_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__15765__B2 _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13313__A2_N _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12528__B _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19349_ _20026_/B _19223_/B _19220_/X _19221_/X fanout96/X vssd1 vssd1 vccd1 vccd1
+ _19354_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11251__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21311_ _21311_/A _21311_/B vssd1 vssd1 vccd1 vccd1 _21319_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout210_A _21815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout308_A _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21242_ _21095_/A _21094_/Y _21093_/B vssd1 vssd1 vccd1 vccd1 _21243_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_4_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold310 hold310/A vssd1 vssd1 vccd1 vccd1 hold310/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 hold321/A vssd1 vssd1 vccd1 vccd1 hold321/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 hold332/A vssd1 vssd1 vccd1 vccd1 hold332/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19972__D _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21173_ _21172_/B _21172_/C _21172_/A vssd1 vssd1 vccd1 vccd1 _21174_/B sky130_fd_sc_hd__a21oi_1
X_20124_ _20124_/A _20124_/B vssd1 vssd1 vccd1 vccd1 _20163_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20055_ _19828_/B _19830_/B _20053_/X _20054_/Y vssd1 vssd1 vccd1 vccd1 _20203_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19431__A2 _19751_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13525__D _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21526__A0 hold309/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_205 hold270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_216 hold275/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_227 hold290/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_238 hold309/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_249 hold262/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20957_ _20822_/Y _20824_/X _20955_/X _20956_/Y vssd1 vssd1 vccd1 vccd1 _20960_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11490__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17013__C _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11690_ _11688_/X _11690_/B vssd1 vssd1 vccd1 vccd1 _11691_/B sky130_fd_sc_hd__and2b_1
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20888_ _20750_/A _20753_/A _20886_/X _20887_/Y vssd1 vssd1 vccd1 vccd1 _20888_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20655__B _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11242__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13360_ _13509_/B _13358_/X _13218_/B _13218_/Y vssd1 vssd1 vccd1 vccd1 _13361_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11242__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18170__A2 _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12990__A1 _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12311_ _12312_/A _13258_/C vssd1 vssd1 vccd1 vccd1 _12313_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_133_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21509_ hold305/X sstream_i[86] _21510_/S vssd1 vssd1 vccd1 vccd1 _22036_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12990__B2 _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13291_ _14027_/A _14537_/A _13290_/C _13290_/D vssd1 vssd1 vccd1 vccd1 _13292_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_1_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_786 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12454__A _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15030_ _15768_/A _14873_/B _14870_/X _14871_/X _16268_/B vssd1 vssd1 vccd1 vccd1
+ _15035_/A sky130_fd_sc_hd__a32o_1
XANTENNA__14192__B1 _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21057__A2 _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12242_ _12267_/A _12242_/B _12269_/C _12269_/D vssd1 vssd1 vccd1 vccd1 _12258_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_121_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13269__B _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20671__A _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20027__A1_N _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12173_ _12169_/X _12172_/X _12128_/B _12131_/Y vssd1 vssd1 vccd1 vccd1 _12173_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_130_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20390__B _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11124_ _11124_/A _11126_/B vssd1 vssd1 vccd1 vccd1 _11124_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_101_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16981_ _16980_/B _16980_/C _16980_/A vssd1 vssd1 vccd1 vccd1 _16982_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_101_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18720_ _18720_/A _18720_/B _18720_/C vssd1 vssd1 vccd1 vccd1 _18720_/X sky130_fd_sc_hd__and3_1
X_15932_ _15933_/C _16391_/B _15930_/Y _16056_/A vssd1 vssd1 vccd1 vccd1 _15934_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_11055_ _11055_/A _11055_/B vssd1 vssd1 vccd1 vccd1 _11055_/Y sky130_fd_sc_hd__xnor2_4
X_15863_ _15721_/Y _15723_/Y _15861_/Y _15862_/X vssd1 vssd1 vccd1 vccd1 _15863_/Y
+ sky130_fd_sc_hd__a211oi_2
X_18651_ _19123_/B _19972_/C _21258_/B _18652_/A vssd1 vssd1 vccd1 vccd1 _18653_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14814_ _14814_/A _14814_/B vssd1 vssd1 vccd1 vccd1 _14824_/A sky130_fd_sc_hd__xor2_2
X_17602_ _17602_/A _17602_/B _17602_/C vssd1 vssd1 vccd1 vccd1 _17603_/B sky130_fd_sc_hd__and3_1
X_15794_ _16369_/A _16040_/C _15794_/C _15794_/D vssd1 vssd1 vccd1 vccd1 _15921_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_8_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18582_ _18582_/A _18582_/B vssd1 vssd1 vccd1 vccd1 _18592_/A sky130_fd_sc_hd__nand2_1
XTAP_3750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15931__C _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14828__B _14828_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14745_ _14746_/A _14746_/B vssd1 vssd1 vccd1 vccd1 _14745_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_87_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17533_ _17534_/A _17534_/B vssd1 vssd1 vccd1 vccd1 _17533_/X sky130_fd_sc_hd__and2_2
XTAP_3794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11957_ _12015_/A _12015_/B vssd1 vssd1 vccd1 vccd1 _11957_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_129_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18933__A1 _19092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18933__B2 _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10908_ _10908_/A _10908_/B vssd1 vssd1 vccd1 vccd1 _10909_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11481__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17464_ _17460_/X _17462_/Y _17351_/B _17351_/Y vssd1 vssd1 vccd1 vccd1 _17466_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_156_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14676_ _15808_/C _16406_/A _14676_/C _14825_/A vssd1 vssd1 vccd1 vccd1 _14825_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__11481__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11888_ _11889_/A _11889_/B _11889_/C vssd1 vssd1 vccd1 vccd1 _11899_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_74_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16415_ _16261_/X _16298_/B _15907_/A _16151_/B vssd1 vssd1 vccd1 vccd1 _16416_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_95_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19203_ _19202_/B _19348_/B _19202_/A vssd1 vssd1 vccd1 vccd1 _19204_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13627_ _13627_/A _13627_/B _13627_/C vssd1 vssd1 vccd1 vccd1 _13630_/A sky130_fd_sc_hd__nand3_1
X_10839_ _10815_/B _11057_/B _10815_/A vssd1 vssd1 vccd1 vccd1 _11059_/A sky130_fd_sc_hd__a21bo_1
X_17395_ _17621_/C _17504_/C _17739_/C _17739_/D vssd1 vssd1 vccd1 vccd1 _17395_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_156_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16346_ _16347_/A _16347_/B _16347_/C vssd1 vssd1 vccd1 vccd1 _16349_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_15_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11233__A1 _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19134_ _19133_/A _19133_/B _19133_/C vssd1 vssd1 vccd1 vccd1 _19135_/C sky130_fd_sc_hd__a21o_1
X_13558_ _13867_/A _14354_/C _14663_/D _13858_/A vssd1 vssd1 vccd1 vccd1 _13558_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__11233__B2 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12981__A1 _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18035__B _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19065_ _19065_/A _19065_/B vssd1 vssd1 vccd1 vccd1 _19073_/A sky130_fd_sc_hd__nand2_1
X_12509_ _12402_/A _12402_/B _12405_/B _12403_/X vssd1 vssd1 vccd1 vccd1 _12519_/A
+ sky130_fd_sc_hd__a31o_1
X_16277_ _16277_/A _16277_/B vssd1 vssd1 vccd1 vccd1 _16278_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12981__B2 _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13489_ _13485_/X _13487_/Y _13338_/B _13338_/Y vssd1 vssd1 vccd1 vccd1 _13491_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21099__D _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15228_ _15632_/B _16414_/B _16391_/B _15892_/A vssd1 vssd1 vccd1 vccd1 _15231_/C
+ sky130_fd_sc_hd__a22o_1
X_18016_ _17878_/A _17878_/C _17878_/B vssd1 vssd1 vccd1 vccd1 _18018_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_11_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17874__B _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19110__A1 _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15159_ _21733_/Q _15838_/B _16314_/D _15159_/D vssd1 vssd1 vccd1 vccd1 _15162_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_11_957 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout108 _19692_/C vssd1 vssd1 vccd1 vccd1 _19227_/C sky130_fd_sc_hd__buf_4
XANTENNA__17672__A1 _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout119 _20146_/B vssd1 vssd1 vccd1 vccd1 _19238_/C sky130_fd_sc_hd__buf_4
X_19967_ _20101_/A _20101_/B _21264_/B vssd1 vssd1 vccd1 vccd1 _19967_/X sky130_fd_sc_hd__and3_1
X_18918_ _18917_/A _18917_/B _18917_/C vssd1 vssd1 vccd1 vccd1 _18919_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__19413__A2 _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19898_ _19898_/A _19898_/B _19898_/C vssd1 vssd1 vccd1 vccd1 _19898_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_98_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18849_ _18849_/A _18849_/B _21848_/Q _19013_/C vssd1 vssd1 vccd1 vccd1 _19017_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__14789__A2 _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21860_ _21932_/CLK _21860_/D vssd1 vssd1 vccd1 vccd1 hold221/A sky130_fd_sc_hd__dfxtp_1
X_20811_ _20814_/D vssd1 vssd1 vccd1 vccd1 _20811_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout160_A _21829_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21791_ _21974_/CLK _21791_/D vssd1 vssd1 vccd1 vccd1 _21791_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_77_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17727__A2 _19692_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout258_A _21803_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14457__C _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11472__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20178__D _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20742_ _20742_/A _20742_/B _20742_/C vssd1 vssd1 vccd1 vccd1 _20742_/X sky130_fd_sc_hd__and3_1
XANTENNA__20731__A1 _20991_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20731__B2 _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18871__D _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20673_ _21258_/A _21153_/B _21264_/B _20797_/A vssd1 vssd1 vccd1 vccd1 _20677_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21039__A2 _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15910__A1 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20922__C _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold140 hold140/A vssd1 vssd1 vccd1 vccd1 hold140/X sky130_fd_sc_hd__dlygate4sd3_1
X_21225_ _21225_/A _21225_/B vssd1 vssd1 vccd1 vccd1 _21226_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12724__B2 _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19057__A _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold151 hold151/A vssd1 vssd1 vccd1 vccd1 hold151/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold162 hold162/A vssd1 vssd1 vccd1 vccd1 hold162/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 hold173/A vssd1 vssd1 vccd1 vccd1 hold173/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 hold184/A vssd1 vssd1 vccd1 vccd1 hold184/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 hold195/A vssd1 vssd1 vccd1 vccd1 hold195/X sky130_fd_sc_hd__dlygate4sd3_1
X_21156_ _21267_/A _21841_/Q _21256_/B vssd1 vssd1 vccd1 vccd1 _21156_/X sky130_fd_sc_hd__and3_1
XFILLER_0_106_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout620 _21717_/Q vssd1 vssd1 vccd1 vccd1 _11039_/S sky130_fd_sc_hd__buf_4
Xfanout631 _21776_/Q vssd1 vssd1 vccd1 vccd1 _13258_/C sky130_fd_sc_hd__clkbuf_8
X_20107_ _20249_/A _20242_/D _20105_/Y _20251_/A vssd1 vssd1 vccd1 vccd1 _20109_/A
+ sky130_fd_sc_hd__o2bb2a_1
Xfanout642 _21329_/B1 vssd1 vssd1 vccd1 vccd1 _11041_/A sky130_fd_sc_hd__clkbuf_4
X_21087_ _20975_/D _21293_/B _21853_/Q _21087_/D vssd1 vssd1 vccd1 vccd1 _21206_/A
+ sky130_fd_sc_hd__and4b_2
XANTENNA_fanout73_A _21849_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20038_ _20039_/A _20039_/B vssd1 vssd1 vccd1 vccd1 _20222_/A sky130_fd_sc_hd__and2_1
XFILLER_0_137_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12860_ _13554_/B _13573_/D _12989_/A _12860_/D vssd1 vssd1 vccd1 vccd1 _12989_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_73_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19168__A1 _17841_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _11810_/B _11810_/C _11810_/A vssd1 vssd1 vccd1 vccd1 _11813_/B sky130_fd_sc_hd__a21bo_1
XTAP_3079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ _12790_/A _12790_/B _12790_/C vssd1 vssd1 vccd1 vccd1 _12792_/C sky130_fd_sc_hd__a21o_1
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21989_ _22020_/CLK _21989_/D vssd1 vssd1 vccd1 vccd1 hold182/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14530_ _14530_/A _14530_/B vssd1 vssd1 vccd1 vccd1 _14531_/B sky130_fd_sc_hd__nor2_2
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11463__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11742_ _11741_/B _11741_/C _11741_/A vssd1 vssd1 vccd1 vccd1 _11744_/B sky130_fd_sc_hd__a21bo_1
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13271__C _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20722__B2 _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14461_ _16084_/C _14306_/X _14309_/A _14309_/B vssd1 vssd1 vccd1 vccd1 _14462_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_83_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11673_ _12094_/A _12094_/B _12444_/B _12443_/A vssd1 vssd1 vccd1 vccd1 _11673_/X
+ sky130_fd_sc_hd__and4_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16200_ _16200_/A _16309_/B vssd1 vssd1 vccd1 vccd1 _16202_/A sky130_fd_sc_hd__or2_2
XFILLER_0_3_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13412_ _13413_/B _13413_/A vssd1 vssd1 vccd1 vccd1 _13539_/A sky130_fd_sc_hd__nand2b_1
X_17180_ _17636_/B _17490_/A _16571_/B _16569_/X vssd1 vssd1 vccd1 vccd1 _17187_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_0_64_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14392_ _14220_/A _14220_/C _14220_/B vssd1 vssd1 vccd1 vccd1 _14393_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_119_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16131_ _16128_/Y _16129_/X _15999_/A _15999_/Y vssd1 vssd1 vccd1 vccd1 _16132_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_148_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12963__A1 _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13343_ _13343_/A _13343_/B _13343_/C _13343_/D vssd1 vssd1 vccd1 vccd1 _13343_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_49_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16062_ _16171_/A _16369_/B _16286_/A _16062_/D vssd1 vssd1 vccd1 vccd1 _16171_/B
+ sky130_fd_sc_hd__and4b_1
X_13274_ _13416_/B _13273_/C _13273_/A vssd1 vssd1 vccd1 vccd1 _13275_/C sky130_fd_sc_hd__o21ai_1
X_15013_ _14887_/B _14889_/A _15010_/Y _15012_/X vssd1 vssd1 vccd1 vccd1 _15013_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_20_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13912__B1 _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12225_ _12219_/A _12219_/B _12219_/C vssd1 vssd1 vccd1 vccd1 _12226_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_121_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19643__A2 _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19821_ _20721_/D _20671_/B _19685_/X _19686_/X _21278_/A vssd1 vssd1 vccd1 vccd1
+ _19826_/A sky130_fd_sc_hd__a32o_1
X_12156_ _12157_/A _12197_/A vssd1 vssd1 vccd1 vccd1 _12156_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_20_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11107_ _10892_/Y hold32/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21701_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19752_ _21833_/Q _19753_/B _19753_/C _19753_/D vssd1 vssd1 vccd1 vccd1 _19752_/X
+ sky130_fd_sc_hd__a22o_1
X_16964_ _16956_/A _16956_/C _16956_/B vssd1 vssd1 vccd1 vccd1 _16964_/X sky130_fd_sc_hd__a21o_1
X_12087_ _12040_/A _12040_/C _12040_/B vssd1 vssd1 vccd1 vccd1 _12093_/B sky130_fd_sc_hd__a21o_1
X_18703_ _18703_/A _19185_/B vssd1 vssd1 vccd1 vccd1 _18705_/B sky130_fd_sc_hd__nand2_1
X_15915_ _16371_/A _16377_/B _16414_/B _16380_/A vssd1 vssd1 vccd1 vccd1 _15919_/C
+ sky130_fd_sc_hd__a22o_1
X_11038_ mstream_o[112] hold277/X _11039_/S vssd1 vssd1 vccd1 vccd1 _21649_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19414__B _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19683_ _19683_/A _19683_/B vssd1 vssd1 vccd1 vccd1 _19773_/A sky130_fd_sc_hd__xnor2_1
X_16895_ _16896_/A _16896_/B vssd1 vssd1 vccd1 vccd1 _16895_/X sky130_fd_sc_hd__and2b_1
XANTENNA__20410__B1 _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18634_ _18631_/X _18632_/Y _18472_/Y _18474_/X vssd1 vssd1 vccd1 vccd1 _18669_/B
+ sky130_fd_sc_hd__o211a_1
X_15846_ _15846_/A _15846_/B vssd1 vssd1 vccd1 vccd1 _15847_/B sky130_fd_sc_hd__and2_1
XFILLER_0_8_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18565_ _18409_/A _18410_/Y _18563_/A _18564_/X vssd1 vssd1 vccd1 vccd1 _18565_/Y
+ sky130_fd_sc_hd__a211oi_1
X_15777_ _15778_/B _15778_/A vssd1 vssd1 vccd1 vccd1 _15777_/Y sky130_fd_sc_hd__nand2b_1
XTAP_3580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12989_ _12989_/A _12989_/B vssd1 vssd1 vccd1 vccd1 _12997_/A sky130_fd_sc_hd__nand2_1
XTAP_3591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17516_ _17426_/X _17429_/Y _17514_/A _17515_/Y vssd1 vssd1 vccd1 vccd1 _17602_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_8_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11454__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19430__A _19430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14728_ _14859_/A _15510_/B _14729_/C _14854_/A vssd1 vssd1 vccd1 vccd1 _14730_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13181__C _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13994__A3 _14477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20713__A1 _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18496_ _18496_/A _18496_/B vssd1 vssd1 vccd1 vccd1 _18505_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20713__B2 _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14659_ _14659_/A _15788_/B vssd1 vssd1 vccd1 vccd1 _14660_/B sky130_fd_sc_hd__nand2_1
X_17447_ _19445_/A _17915_/D vssd1 vssd1 vccd1 vccd1 _17450_/A sky130_fd_sc_hd__and2_1
XFILLER_0_28_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17378_ _21142_/A _21340_/B vssd1 vssd1 vccd1 vccd1 _17378_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_83_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12954__A1 _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11757__A2 _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19117_ _19587_/A _19587_/B _20249_/B vssd1 vssd1 vccd1 vccd1 _19117_/X sky130_fd_sc_hd__and3_1
XANTENNA__11710__B _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16329_ _16329_/A _16329_/B vssd1 vssd1 vccd1 vccd1 _16331_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12954__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19048_ _19048_/A _19048_/B vssd1 vssd1 vccd1 vccd1 _19148_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_152_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21010_ _20877_/B _20880_/B _21008_/Y _21009_/X vssd1 vssd1 vccd1 vccd1 _21012_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12182__A2 _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15309__A2_N _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13131__A1 _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13131__B2 _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15408__B1 _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout375_A _14828_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21912_ _21945_/CLK _21912_/D vssd1 vssd1 vccd1 vccd1 hold226/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11693__A1 _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11693__B2 _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21843_ _21845_/CLK _21843_/D vssd1 vssd1 vccd1 vccd1 _21843_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_136_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout542_A _21735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21774_ _21789_/CLK _21774_/D vssd1 vssd1 vccd1 vccd1 _21774_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__11604__C _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19570__A1 _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19570__B2 _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20725_ _20594_/A _20593_/A _20593_/B _20589_/B _20589_/A vssd1 vssd1 vccd1 vccd1
+ _20726_/B sky130_fd_sc_hd__o32ai_4
XFILLER_0_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15187__A2 _15050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19337__A_N _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20656_ _20656_/A _20656_/B vssd1 vssd1 vccd1 vccd1 _20658_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20587_ _20587_/A _20719_/B vssd1 vssd1 vccd1 vccd1 _20589_/A sky130_fd_sc_hd__or2_2
XANTENNA__17333__B1 _17443_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19873__A2 _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13370__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ _11999_/A _11999_/C _11999_/B vssd1 vssd1 vccd1 vccd1 _12011_/C sky130_fd_sc_hd__a21o_1
XANTENNA__16439__A2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21208_ _21208_/A _21208_/B vssd1 vssd1 vccd1 vccd1 _21218_/A sky130_fd_sc_hd__or2_1
XANTENNA__13370__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17019__B _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11920__A2 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21139_ _21026_/B _21027_/A _21138_/X _21025_/B _21137_/Y vssd1 vssd1 vccd1 vccd1
+ _21141_/A sky130_fd_sc_hd__a221oi_1
Xfanout450 _14248_/A vssd1 vssd1 vccd1 vccd1 _12269_/A sky130_fd_sc_hd__buf_2
Xfanout461 _16369_/B vssd1 vssd1 vccd1 vccd1 _15368_/D sky130_fd_sc_hd__buf_4
XANTENNA__19389__A1 _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout472 _15091_/C vssd1 vssd1 vccd1 vccd1 _16377_/B sky130_fd_sc_hd__buf_2
XANTENNA__19389__B2 _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13961_ _13962_/A _13962_/B vssd1 vssd1 vccd1 vccd1 _14290_/B sky130_fd_sc_hd__and2b_1
Xfanout483 _21748_/Q vssd1 vssd1 vccd1 vccd1 _14873_/B sky130_fd_sc_hd__buf_4
XANTENNA__14659__A _14659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout494 _21745_/Q vssd1 vssd1 vccd1 vccd1 _14386_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__14870__A1 _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15700_ _15700_/A _15700_/B vssd1 vssd1 vccd1 vccd1 _15701_/B sky130_fd_sc_hd__nor2_2
X_12912_ _14087_/A _14391_/B _13913_/C _14089_/A vssd1 vssd1 vccd1 vccd1 _12913_/C
+ sky130_fd_sc_hd__a22o_1
X_16680_ _16680_/A _16680_/B vssd1 vssd1 vccd1 vccd1 _16682_/C sky130_fd_sc_hd__xnor2_1
X_13892_ _14365_/A _14212_/B _14365_/D _14384_/A vssd1 vssd1 vccd1 vccd1 _13892_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20943__A1 _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15631_ _15632_/B _16177_/B _16286_/B _15892_/A vssd1 vssd1 vccd1 vccd1 _15635_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12843_ _13394_/A _13997_/C _12839_/X _12841_/Y vssd1 vssd1 vccd1 vccd1 _12844_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15562_ _15561_/B _15561_/C _15561_/A vssd1 vssd1 vccd1 vccd1 _15562_/Y sky130_fd_sc_hd__a21oi_2
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18350_ _18652_/A _18498_/B _19874_/B _19872_/C vssd1 vssd1 vccd1 vccd1 _18352_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_51_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ _13018_/B _21766_/Q _12896_/A _12773_/D vssd1 vssd1 vccd1 vccd1 _12774_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14513_ _14513_/A _14513_/B vssd1 vssd1 vccd1 vccd1 _14521_/A sky130_fd_sc_hd__nand2_1
X_17301_ _17393_/A vssd1 vssd1 vccd1 vccd1 _17301_/Y sky130_fd_sc_hd__inv_2
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11725_ _12458_/A _13173_/C _12357_/C _13155_/A vssd1 vssd1 vccd1 vccd1 _11727_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_68_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15493_ _14916_/A _14916_/B _15492_/A _15207_/Y _15492_/B vssd1 vssd1 vccd1 vccd1
+ _15496_/B sky130_fd_sc_hd__a2111o_1
X_18281_ _18849_/B _19223_/B _18281_/C _18281_/D vssd1 vssd1 vccd1 vccd1 _18282_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_12_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12907__A _14712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14444_ _14446_/A _14446_/B _14446_/C vssd1 vssd1 vccd1 vccd1 _14445_/A sky130_fd_sc_hd__o21ai_2
X_17232_ _17434_/B _18058_/A vssd1 vssd1 vccd1 vccd1 _17236_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_154_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11656_ _11799_/A _11799_/B _11655_/A vssd1 vssd1 vccd1 vccd1 _11670_/A sky130_fd_sc_hd__o21ai_2
Xfanout90 _21844_/Q vssd1 vssd1 vccd1 vccd1 _18894_/B sky130_fd_sc_hd__buf_4
XFILLER_0_117_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17163_ _17050_/X _17162_/X _17007_/X vssd1 vssd1 vccd1 vccd1 _17163_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14375_ _14375_/A _14375_/B _14375_/C vssd1 vssd1 vccd1 vccd1 _14375_/X sky130_fd_sc_hd__and3_1
XFILLER_0_25_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11587_ _12319_/C _12420_/D _12511_/A _12268_/B vssd1 vssd1 vccd1 vccd1 _11588_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__12400__A3 _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16114_ _16114_/A _16114_/B _16114_/C vssd1 vssd1 vccd1 vccd1 _16114_/X sky130_fd_sc_hd__and3_1
X_13326_ _14087_/A _14234_/C _15370_/B _14089_/A vssd1 vssd1 vccd1 vccd1 _13327_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17875__A1 _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17094_ _17094_/A _17094_/B vssd1 vssd1 vccd1 vccd1 _17097_/A sky130_fd_sc_hd__nor2_1
XANTENNA__19409__B _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18313__B _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16045_ _16380_/A _16371_/A _16414_/B _16391_/B vssd1 vssd1 vccd1 vccd1 _16165_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__20562__C _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13257_ _13257_/A _13257_/B vssd1 vssd1 vccd1 vccd1 _13266_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12642__A _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12208_ _12207_/B _12206_/Y _12168_/X _12176_/Y vssd1 vssd1 vccd1 vccd1 _12208_/X
+ sky130_fd_sc_hd__o211a_1
X_13188_ _13188_/A _13188_/B _13188_/C vssd1 vssd1 vccd1 vccd1 _13191_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_23_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__22067__RESET_B fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19804_ _20032_/D _20841_/B _19804_/C _19804_/D vssd1 vssd1 vccd1 vccd1 _19808_/B
+ sky130_fd_sc_hd__nand4_2
X_12139_ _12139_/A _12139_/B _12139_/C vssd1 vssd1 vccd1 vccd1 _12185_/A sky130_fd_sc_hd__nand3_1
X_17996_ _18849_/A _19382_/B vssd1 vssd1 vccd1 vccd1 _17999_/A sky130_fd_sc_hd__and2_1
XANTENNA__16768__B _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19735_ _19735_/A _19735_/B _19849_/B vssd1 vssd1 vccd1 vccd1 _19737_/B sky130_fd_sc_hd__nand3_1
X_16947_ _16890_/A _16890_/C _16890_/B vssd1 vssd1 vccd1 vccd1 _16947_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13473__A _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16487__C _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19666_ _20026_/B _20193_/D _19666_/C _19820_/A vssd1 vssd1 vccd1 vccd1 _19820_/B
+ sky130_fd_sc_hd__nand4_2
X_16878_ _16989_/C _17123_/C _16815_/C _16815_/D vssd1 vssd1 vccd1 vccd1 _16879_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18617_ _18617_/A vssd1 vssd1 vccd1 vccd1 _18618_/B sky130_fd_sc_hd__inv_2
X_15829_ _16203_/D _16092_/D _15829_/C _16084_/D vssd1 vssd1 vccd1 vccd1 _15959_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__12089__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19597_ _19597_/A _19597_/B vssd1 vssd1 vccd1 vccd1 _19609_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_59_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18548_ _18548_/A _18548_/B vssd1 vssd1 vccd1 vccd1 _18550_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17599__B _17599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21631__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18479_ _18323_/X _18325_/X _18477_/Y _18478_/X vssd1 vssd1 vccd1 vccd1 _18516_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_118_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11721__A _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20510_ _20639_/B _20508_/X _20363_/A _20367_/A vssd1 vssd1 vccd1 vccd1 _20511_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_142_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21490_ hold192/X sstream_i[67] _21490_/S vssd1 vssd1 vccd1 vccd1 _22017_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20441_ _20441_/A _20441_/B _20441_/C vssd1 vssd1 vccd1 vccd1 _20444_/A sky130_fd_sc_hd__and3_1
XFILLER_0_144_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout123_A _20689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20372_ _20372_/A _20372_/B vssd1 vssd1 vccd1 vccd1 _20372_/X sky130_fd_sc_hd__or2_1
XFILLER_0_67_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16024__A fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22042_ _22049_/CLK _22042_/D vssd1 vssd1 vccd1 vccd1 hold245/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__21414__A2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20191__D _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout492_A _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18596__D _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11115__A0 _10950_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14479__A _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21719__RESET_B _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13407__A2 _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19070__A _19379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21826_ _21829_/CLK _21826_/D vssd1 vssd1 vccd1 vccd1 _21826_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_149_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout36_A _21490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18346__A2 _19868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21757_ _22063_/CLK _21757_/D vssd1 vssd1 vccd1 vccd1 hold313/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_66_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21350__A1 _21407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11510_ _21723_/D t1y[20] t0x[20] _11223_/A vssd1 vssd1 vccd1 vccd1 _11510_/X sky130_fd_sc_hd__a22o_1
XANTENNA__18113__A2_N _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20708_ _20708_/A _20836_/B _20708_/C vssd1 vssd1 vccd1 vccd1 _20710_/A sky130_fd_sc_hd__or3_1
XFILLER_0_19_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12490_ _12708_/B _12490_/B vssd1 vssd1 vccd1 vccd1 _12497_/B sky130_fd_sc_hd__xor2_4
XANTENNA__20944__A _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21688_ _22069_/CLK _21688_/D vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout2_A fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11441_ _11447_/A1 hold175/A fanout49/X hold180/A vssd1 vssd1 vccd1 vccd1 _11441_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20639_ _20639_/A _20639_/B vssd1 vssd1 vccd1 vccd1 _20641_/B sky130_fd_sc_hd__or2_2
XFILLER_0_151_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16860__C _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14160_ _14160_/A _14160_/B _14160_/C vssd1 vssd1 vccd1 vccd1 _14162_/B sky130_fd_sc_hd__nand3_2
X_11372_ _11124_/A hold231/X fanout45/X hold204/X vssd1 vssd1 vccd1 vccd1 _11372_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19229__B _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13111_ _13111_/A _13111_/B vssd1 vssd1 vccd1 vccd1 _13112_/B sky130_fd_sc_hd__xor2_2
XANTENNA__18133__B _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1138 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14091_ _14090_/B _14090_/C _14090_/A vssd1 vssd1 vccd1 vccd1 _14093_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_131_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13042_ _13042_/A _13042_/B vssd1 vssd1 vccd1 vccd1 _13062_/A sky130_fd_sc_hd__nor2_1
XANTENNA__12181__B _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19890__D _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17850_ _17850_/A _17850_/B vssd1 vssd1 vccd1 vccd1 _17852_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__18787__C _21040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16801_ _16800_/A _16800_/C _16800_/B vssd1 vssd1 vccd1 vccd1 _16806_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11106__A0 _10886_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17781_ _20583_/A _18789_/A _17913_/A _17780_/D vssd1 vssd1 vccd1 vccd1 _17781_/X
+ sky130_fd_sc_hd__a22o_1
X_14993_ _14993_/A _15892_/B _16268_/B _16266_/C vssd1 vssd1 vccd1 vccd1 _14994_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__14389__A _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout280 _19644_/A vssd1 vssd1 vccd1 vccd1 _20178_/D sky130_fd_sc_hd__clkbuf_8
Xfanout291 _17874_/A vssd1 vssd1 vccd1 vccd1 _19810_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__18034__A1 _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19520_ _19521_/A _19521_/B vssd1 vssd1 vccd1 vccd1 _19520_/Y sky130_fd_sc_hd__nor2_1
X_16732_ _17096_/A _16968_/C vssd1 vssd1 vccd1 vccd1 _16737_/A sky130_fd_sc_hd__nand2_1
XANTENNA__18034__B2 _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__A1 _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13944_ _13943_/A _13943_/B _13941_/X _13942_/Y vssd1 vssd1 vccd1 vccd1 _13944_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_89_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19451_ _19452_/B _19452_/A vssd1 vssd1 vccd1 vccd1 _19451_/X sky130_fd_sc_hd__and2b_1
X_13875_ _21741_/Q _13875_/B _14516_/A _14365_/C vssd1 vssd1 vccd1 vccd1 _14032_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_88_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16663_ _16662_/B _16662_/C _16662_/A vssd1 vssd1 vccd1 vccd1 _16665_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__20392__A2 _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20838__B _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18402_ _18402_/A _18402_/B vssd1 vssd1 vccd1 vccd1 _18411_/A sky130_fd_sc_hd__or2_1
X_15614_ _15475_/A _15475_/Y _15612_/Y _15613_/X vssd1 vssd1 vccd1 vccd1 _15614_/Y
+ sky130_fd_sc_hd__a211oi_4
X_12826_ _12957_/B _12710_/B _12825_/X vssd1 vssd1 vccd1 vccd1 _12827_/B sky130_fd_sc_hd__o21a_2
X_19382_ _19382_/A _19382_/B _19382_/C _19382_/D vssd1 vssd1 vccd1 vccd1 _19382_/Y
+ sky130_fd_sc_hd__nand4_1
X_16594_ _16592_/X _16594_/B vssd1 vssd1 vccd1 vccd1 _16595_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_96_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18337__A2 _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18333_ _19723_/A _18640_/B _18199_/B _18197_/X vssd1 vssd1 vccd1 vccd1 _18341_/A
+ sky130_fd_sc_hd__a31o_1
X_15545_ _15545_/A _15545_/B vssd1 vssd1 vccd1 vccd1 _15546_/B sky130_fd_sc_hd__nand2_1
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ _14024_/B _13155_/C _13155_/D _13013_/A vssd1 vssd1 vccd1 vccd1 _12757_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21341__A1 _21349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12637__A _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11708_ _11709_/A _11707_/Y _12223_/A _12443_/A vssd1 vssd1 vccd1 vccd1 _11747_/A
+ sky130_fd_sc_hd__and4bb_1
X_15476_ _15475_/A _15475_/B _15475_/C _15475_/D vssd1 vssd1 vccd1 vccd1 _15476_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18264_ _18265_/A _18265_/B vssd1 vssd1 vccd1 vccd1 _18264_/X sky130_fd_sc_hd__or2_1
XFILLER_0_44_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12688_ _12687_/B _12687_/C _12687_/A vssd1 vssd1 vccd1 vccd1 _12688_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_126_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12356__B _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14427_ _14427_/A _14427_/B vssd1 vssd1 vccd1 vccd1 _14430_/A sky130_fd_sc_hd__xnor2_4
X_17215_ _17215_/A _17215_/B vssd1 vssd1 vccd1 vccd1 _17217_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11639_ _12528_/B _12020_/A _13155_/D _12619_/A vssd1 vssd1 vccd1 vccd1 _11640_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__15571__A2 _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18195_ _18195_/A _18195_/B vssd1 vssd1 vccd1 vccd1 _18215_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_154_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14358_ _14181_/X _14184_/X _14355_/X _14357_/Y vssd1 vssd1 vccd1 vccd1 _14358_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17146_ _17146_/A _17146_/B _17146_/C _17146_/D vssd1 vssd1 vccd1 vccd1 _17146_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_13_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13468__A _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13309_ _13184_/A _13183_/B _13183_/A vssd1 vssd1 vccd1 vccd1 _13316_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17077_ _17078_/A _17078_/B _17078_/C vssd1 vssd1 vccd1 vccd1 _17077_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_40_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14289_ _14289_/A _14289_/B vssd1 vssd1 vccd1 vccd1 _14913_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__16520__A1 _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16520__B2 _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16028_ _16028_/A _16028_/B vssd1 vssd1 vccd1 vccd1 _16029_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20604__B1 _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13915__B _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17979_ _17980_/A _17980_/B _17980_/C vssd1 vssd1 vccd1 vccd1 _18120_/A sky130_fd_sc_hd__o21ai_2
X_19718_ _19715_/Y _19716_/X _19580_/X _19585_/A vssd1 vssd1 vccd1 vccd1 _19719_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_137_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20990_ _21291_/A _21311_/B _20988_/Y _21096_/A vssd1 vssd1 vccd1 vccd1 _20992_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19649_ _19649_/A _19649_/B vssd1 vssd1 vccd1 vccd1 _19654_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_133_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21611_ _21934_/CLK _21611_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[74] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20135__A2 _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21332__A1 _21407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout338_A _15174_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1015 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21542_ mstream_o[5] hold15/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22069_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_30_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21473_ hold162/X sstream_i[50] _21481_/S vssd1 vssd1 vccd1 vccd1 _22000_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout505_A _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20424_ _20425_/A _20425_/B vssd1 vssd1 vccd1 vccd1 _20616_/B sky130_fd_sc_hd__or2_1
XFILLER_0_71_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20355_ _20354_/Y _20355_/B _20355_/C vssd1 vssd1 vccd1 vccd1 _20355_/Y sky130_fd_sc_hd__nand3b_4
XFILLER_0_144_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11336__A0 _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17792__B _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20286_ _21839_/Q _21305_/A _20284_/Y _20427_/A vssd1 vssd1 vccd1 vccd1 _20288_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13876__A2 _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16689__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22025_ _22038_/CLK _22025_/D vssd1 vssd1 vccd1 vccd1 hold261/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__15078__A1 _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18400__C _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16814__A2 _17063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20004__A _20689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold66 hold66/A vssd1 vssd1 vccd1 vccd1 hold66/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 hold77/A vssd1 vssd1 vccd1 vccd1 hold77/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 hold88/A vssd1 vssd1 vccd1 vccd1 hold88/X sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ _12094_/A _12639_/A _12530_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _11992_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_98_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold99 hold99/A vssd1 vssd1 vccd1 vccd1 hold99/X sky130_fd_sc_hd__dlygate4sd3_1
X_10941_ _10945_/B _10941_/B vssd1 vssd1 vccd1 vccd1 _10941_/X sky130_fd_sc_hd__and2_2
XFILLER_0_39_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21571__A1 _11048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13660_ _13813_/A _13660_/B vssd1 vssd1 vccd1 vccd1 _13662_/B sky130_fd_sc_hd__and2_2
X_10872_ _10873_/A _10873_/B _10873_/C vssd1 vssd1 vccd1 vccd1 _10880_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_112_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12611_ _13983_/B _14018_/C _12610_/C _12610_/D vssd1 vssd1 vccd1 vccd1 _12612_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_156_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21809_ _21809_/CLK _21809_/D vssd1 vssd1 vccd1 vccd1 _21809_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13591_ _13875_/B _14537_/A _13591_/C _13591_/D vssd1 vssd1 vccd1 vccd1 _13592_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_13_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18052__A2_N _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12457__A _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15330_ _15327_/Y _15328_/X _15177_/B _15179_/B vssd1 vssd1 vccd1 vccd1 _15332_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12542_ _12542_/A _12542_/B vssd1 vssd1 vccd1 vccd1 _12544_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20674__A _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15768__A _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15261_ _15791_/A _16371_/A _16305_/B _16399_/A vssd1 vssd1 vccd1 vccd1 _15400_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_151_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12473_ _12370_/B _12370_/Y _12470_/X _12472_/Y vssd1 vssd1 vccd1 vccd1 _12475_/C
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__12607__D _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20393__B _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14212_ _14384_/A _14212_/B _14212_/C _14212_/D vssd1 vssd1 vccd1 vccd1 _14213_/B
+ sky130_fd_sc_hd__nand4_1
X_17000_ _17005_/A _17000_/B vssd1 vssd1 vccd1 vccd1 _17002_/B sky130_fd_sc_hd__nand2_1
X_11424_ hold233/A fanout29/X _11423_/X vssd1 vssd1 vccd1 vccd1 _11424_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_152_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15192_ _15192_/A _15192_/B vssd1 vssd1 vccd1 vccd1 _15195_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__14761__B1 _10903_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14391__B _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_8 _11331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18697__A2_N _19181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14143_ _14144_/A _14144_/B vssd1 vssd1 vccd1 vccd1 _14317_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11355_ hold200/X fanout29/X _11354_/X vssd1 vssd1 vccd1 vccd1 _11355_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_105_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11300__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14074_ _14557_/A _14234_/C _15001_/B _14848_/A vssd1 vssd1 vccd1 vccd1 _14077_/C
+ sky130_fd_sc_hd__a22o_1
X_18951_ _19732_/B _19866_/C _18951_/C _19106_/A vssd1 vssd1 vccd1 vccd1 _19106_/B
+ sky130_fd_sc_hd__nand4_2
X_11286_ _11493_/A1 t1x[15] v2z[15] _11507_/B2 _11285_/X vssd1 vssd1 vccd1 vccd1 _11286_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__11327__B1 _11326_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ _13025_/A _13148_/A _13025_/C vssd1 vssd1 vccd1 vccd1 _13148_/B sky130_fd_sc_hd__nand3_2
XANTENNA__18255__A1 _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17902_ _17901_/B _17901_/C _17901_/A vssd1 vssd1 vccd1 vccd1 _17904_/B sky130_fd_sc_hd__a21o_1
XANTENNA__18255__B2 _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18882_ _18878_/X _18879_/Y _18716_/A _18717_/Y vssd1 vssd1 vccd1 vccd1 _18882_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_20_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17833_ _20770_/B _21349_/B vssd1 vssd1 vccd1 vccd1 _17833_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17207__B _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18007__A1 _18008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18007__B2 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19703__A _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17764_ _19892_/A _18319_/B _18622_/B _19823_/A vssd1 vssd1 vccd1 vccd1 _17765_/C
+ sky130_fd_sc_hd__a22o_1
X_14976_ _14976_/A _14976_/B vssd1 vssd1 vccd1 vccd1 _14984_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_107_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_40_clk_i _21822_/CLK vssd1 vssd1 vccd1 vccd1 _21789_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19503_ _19386_/A _19385_/B _19383_/X vssd1 vssd1 vccd1 vccd1 _19503_/Y sky130_fd_sc_hd__a21oi_1
X_16715_ _16715_/A _16715_/B _16715_/C vssd1 vssd1 vccd1 vccd1 _16716_/B sky130_fd_sc_hd__and3_1
X_13927_ _14248_/A _21759_/Q _15234_/C _14250_/B vssd1 vssd1 vccd1 vccd1 _13928_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_89_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13173__D _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17695_ _17718_/B _17694_/B _17693_/C _17693_/D vssd1 vssd1 vccd1 vccd1 _17695_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XANTENNA__18319__A _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_44_clk_i_A _21822_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17223__A _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19434_ _19433_/B _19598_/B _19433_/A vssd1 vssd1 vccd1 vccd1 _19435_/B sky130_fd_sc_hd__a21o_1
X_16646_ _16645_/B _16645_/C _16645_/A vssd1 vssd1 vccd1 vccd1 _16648_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13858_ _13858_/A _13858_/B _13858_/C _16414_/A vssd1 vssd1 vccd1 vccd1 _13859_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__14566__B _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20287__C _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19365_ _19365_/A _19365_/B vssd1 vssd1 vccd1 vccd1 _19366_/B sky130_fd_sc_hd__xnor2_1
X_12809_ _12837_/B _12808_/B _12807_/C _12807_/D vssd1 vssd1 vccd1 vccd1 _12809_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
X_16577_ _16522_/A _16522_/B _16522_/C vssd1 vssd1 vccd1 vccd1 _16578_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_130_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13789_ _13790_/A _13790_/B _13790_/C vssd1 vssd1 vccd1 vccd1 _13789_/X sky130_fd_sc_hd__and3_1
XFILLER_0_85_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18316_ _18316_/A _18316_/B vssd1 vssd1 vccd1 vccd1 _18326_/A sky130_fd_sc_hd__and2_1
X_15528_ _15529_/A _15529_/B vssd1 vssd1 vccd1 vccd1 _15528_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_139_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19296_ _19296_/A _19296_/B vssd1 vssd1 vccd1 vccd1 _19299_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_115_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15678__A _15678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18247_ _20770_/B _21358_/B _18246_/X vssd1 vssd1 vccd1 vccd1 _18247_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_154_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15459_ _15459_/A _15459_/B vssd1 vssd1 vccd1 vccd1 _15461_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21399__B _21399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13555__A1 _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18178_ _18179_/A _18179_/B vssd1 vssd1 vccd1 vccd1 _18178_/X sky130_fd_sc_hd__and2_2
XFILLER_0_13_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17893__A _18008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17129_ _17144_/A _17129_/B _17146_/C _17146_/D vssd1 vssd1 vccd1 vccd1 _17130_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_13_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11210__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20179__A2_N _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20140_ _20140_/A _20140_/B vssd1 vssd1 vccd1 vccd1 _20142_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_111_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18246__B2 _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20071_ _20072_/A _20072_/B _20072_/C vssd1 vssd1 vccd1 vccd1 _20224_/A sky130_fd_sc_hd__a21o_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19994__A1 _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16659__D _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout288_A _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20973_ _20972_/B _20973_/B vssd1 vssd1 vccd1 vccd1 _21091_/A sky130_fd_sc_hd__and2b_1
XANTENNA_fanout455_A _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20478__B _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17221__A2 _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19051__C _19051_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout622_A _21822_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21525_ hold275/X sstream_i[102] _21528_/S vssd1 vssd1 vccd1 vccd1 _22052_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_118_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12427__D _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21102__B _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21456_ hold213/X sstream_i[33] _21489_/S vssd1 vssd1 vccd1 vccd1 _21983_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18485__A1 _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20407_ _20407_/A _20407_/B vssd1 vssd1 vccd1 vccd1 _20408_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_102_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21387_ _21420_/S _21387_/B vssd1 vssd1 vccd1 vccd1 _21387_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15299__A1 _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15299__B2 _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20941__B _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11140_ hold177/X fanout23/X _11139_/X vssd1 vssd1 vccd1 vccd1 _11140_/X sky130_fd_sc_hd__a21o_1
X_20338_ _20338_/A _20338_/B vssd1 vssd1 vccd1 vccd1 _20340_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__19507__B _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13258__D _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11071_ _10874_/Y hold10/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21666_/D sky130_fd_sc_hd__mux2_1
X_20269_ _20416_/B _20270_/C _20924_/A _20416_/A vssd1 vssd1 vccd1 vccd1 _20273_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19226__C _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22008_ _22013_/CLK _22008_/D vssd1 vssd1 vccd1 vccd1 hold178/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__18788__A2 _18789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16569__D _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14830_ _15808_/C _16404_/A _14830_/C _15029_/A vssd1 vssd1 vccd1 vccd1 _15029_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_76_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20669__A _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14761_ _21720_/Q hold169/A _10903_/Y fanout6/X _14760_/Y vssd1 vssd1 vccd1 vccd1
+ _14761_/X sky130_fd_sc_hd__a221o_1
X_11973_ _11971_/A _11982_/A _11972_/Y _11901_/X vssd1 vssd1 vccd1 vccd1 _11976_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13571__A _13877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16500_ _17493_/A _17739_/C _17739_/D _17387_/A vssd1 vssd1 vccd1 vccd1 _16500_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__20388__B _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13712_ _13709_/Y _13710_/X _13858_/A _16273_/A vssd1 vssd1 vccd1 vccd1 _13713_/B
+ sky130_fd_sc_hd__and4bb_1
X_10924_ _10924_/A _10924_/B vssd1 vssd1 vccd1 vccd1 _10926_/B sky130_fd_sc_hd__nor2_2
X_14692_ _15632_/B _16326_/A _16418_/A _15892_/A vssd1 vssd1 vccd1 vccd1 _14692_/X
+ sky130_fd_sc_hd__a22o_1
X_17480_ _17590_/A _17593_/B vssd1 vssd1 vccd1 vccd1 _17481_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_129_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14386__B _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16431_ _16431_/A _16431_/B vssd1 vssd1 vccd1 vccd1 _16432_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13290__B _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13643_ _13643_/A _13643_/B _13643_/C _13643_/D vssd1 vssd1 vccd1 vccd1 _13643_/X
+ sky130_fd_sc_hd__or4_2
X_10855_ hold29/A hold22/A vssd1 vssd1 vccd1 vccd1 _10857_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_116_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16882__A _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19150_ _18985_/Y _18987_/X _19148_/X _19149_/Y vssd1 vssd1 vccd1 vccd1 _19152_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13574_ _13437_/D _13439_/A _13572_/X _13720_/B vssd1 vssd1 vccd1 vccd1 _13732_/A
+ sky130_fd_sc_hd__a211o_1
X_16362_ _16362_/A _16362_/B vssd1 vssd1 vccd1 vccd1 _16362_/Y sky130_fd_sc_hd__xnor2_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18101_ _18101_/A _18243_/B vssd1 vssd1 vccd1 vccd1 _18101_/X sky130_fd_sc_hd__xor2_4
XANTENNA__18712__A2 _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15313_ _15314_/A _15314_/B vssd1 vssd1 vccd1 vccd1 _15313_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12525_ _12522_/Y _12523_/X _12436_/X _12439_/Y vssd1 vssd1 vccd1 vccd1 _12526_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16293_ _16293_/A _16293_/B vssd1 vssd1 vccd1 vccd1 _16294_/B sky130_fd_sc_hd__and2_1
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19081_ _19078_/X _19079_/Y _18944_/B _18946_/A vssd1 vssd1 vccd1 vccd1 _19082_/B
+ sky130_fd_sc_hd__o211ai_1
X_18032_ _18032_/A _18032_/B vssd1 vssd1 vccd1 vccd1 _18040_/A sky130_fd_sc_hd__xnor2_1
X_15244_ _15244_/A _15244_/B vssd1 vssd1 vccd1 vccd1 _15247_/B sky130_fd_sc_hd__xnor2_2
X_12456_ _12456_/A _12456_/B vssd1 vssd1 vccd1 vccd1 _12465_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_140_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ _11406_/X _17915_/A _11446_/S vssd1 vssd1 vccd1 vccd1 _21807_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_140_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15175_ _15175_/A _15175_/B _15316_/B vssd1 vssd1 vccd1 vccd1 _15177_/B sky130_fd_sc_hd__or3_2
XFILLER_0_50_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12387_ _12708_/A _12387_/B vssd1 vssd1 vccd1 vccd1 _12496_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12353__C _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20283__A1 _20562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14126_ _14126_/A _14126_/B vssd1 vssd1 vccd1 vccd1 _14126_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_1_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11338_ _11544_/A1 t1x[28] v2z[28] _11543_/B2 _11337_/X vssd1 vssd1 vccd1 vccd1 _11338_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__20283__B2 _20689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12760__A2 _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19983_ _19984_/A _19984_/B _20126_/B _19984_/D vssd1 vssd1 vccd1 vccd1 _19983_/Y
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__19417__B _19868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14057_ _14057_/A _14057_/B vssd1 vssd1 vccd1 vccd1 _14066_/A sky130_fd_sc_hd__xor2_1
X_18934_ _20088_/A _19092_/A _19092_/C _19262_/C vssd1 vssd1 vccd1 vccd1 _18936_/C
+ sky130_fd_sc_hd__nand4_2
X_11269_ _11325_/A1 t2y[11] t0y[11] _11498_/A1 vssd1 vssd1 vccd1 vccd1 _11269_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13008_ _13097_/A _13006_/Y _12866_/Y _12869_/X vssd1 vssd1 vccd1 vccd1 _13009_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__16479__D _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18865_ _18866_/A _18866_/B _18866_/C vssd1 vssd1 vccd1 vccd1 _19159_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_118_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11720__B1 _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17816_ _17852_/B _17815_/B _17815_/C _17815_/D vssd1 vssd1 vccd1 vccd1 _17816_/Y
+ sky130_fd_sc_hd__a22oi_2
X_18796_ _18794_/Y _18795_/X _19723_/A _19753_/B vssd1 vssd1 vccd1 vccd1 _18798_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_118_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17747_ _17749_/A _17749_/B _17749_/C vssd1 vssd1 vccd1 vccd1 _17747_/Y sky130_fd_sc_hd__a21oi_1
X_14959_ _14793_/B _14795_/B _14956_/X _14957_/Y vssd1 vssd1 vccd1 vccd1 _14959_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17678_ _17678_/A _17678_/B _17678_/C vssd1 vssd1 vccd1 vccd1 _17681_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_134_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14017__A2 _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19417_ _20650_/A _19868_/B _19417_/C _19417_/D vssd1 vssd1 vccd1 vccd1 _19417_/X
+ sky130_fd_sc_hd__and4_2
XANTENNA__14727__D _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16629_ _16629_/A _16629_/B _16629_/C vssd1 vssd1 vccd1 vccd1 _16648_/A sky130_fd_sc_hd__nand3_2
XANTENNA__12097__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12528__C _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19348_ _19348_/A _19348_/B vssd1 vssd1 vccd1 vccd1 _19356_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19279_ _19430_/A _19951_/B _19751_/C _20242_/C vssd1 vssd1 vccd1 vccd1 _19427_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_5_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21310_ _21310_/A _21310_/B vssd1 vssd1 vccd1 vccd1 _21320_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13528__B2 _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold300 hold300/A vssd1 vssd1 vccd1 vccd1 hold300/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21241_ _21239_/Y _21241_/B vssd1 vssd1 vccd1 vccd1 _21243_/A sky130_fd_sc_hd__and2b_1
Xhold311 hold311/A vssd1 vssd1 vccd1 vccd1 hold311/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout203_A _21817_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold322 hold322/A vssd1 vssd1 vccd1 vccd1 hold322/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold333 hold333/A vssd1 vssd1 vccd1 vccd1 hold333/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21172_ _21172_/A _21172_/B _21172_/C vssd1 vssd1 vccd1 vccd1 _21174_/A sky130_fd_sc_hd__and3_1
XFILLER_0_29_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20123_ _20124_/A _20124_/B vssd1 vssd1 vccd1 vccd1 _20123_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_141_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12560__A _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20054_ _20186_/B _20053_/C _20053_/A vssd1 vssd1 vccd1 vccd1 _20054_/Y sky130_fd_sc_hd__a21oi_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout572_A _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_206 hold270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_217 hold277/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_228 hold290/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_239 hold309/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20956_ _20953_/A _20954_/Y _20784_/A _20785_/Y vssd1 vssd1 vccd1 vccd1 _20956_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__13822__C _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18393__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20887_ _21016_/B _20885_/Y _20755_/A _20755_/Y vssd1 vssd1 vccd1 vccd1 _20887_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17013__D _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12310_ _12310_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12313_/A sky130_fd_sc_hd__xor2_2
X_21508_ hold280/X sstream_i[85] _21510_/S vssd1 vssd1 vccd1 vccd1 _22035_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13290_ _14027_/A _14537_/A _13290_/C _13290_/D vssd1 vssd1 vccd1 vccd1 _13292_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12990__A2 _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12454__B _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14192__A1 _21743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12241_ _12241_/A _12241_/B vssd1 vssd1 vccd1 vccd1 _12241_/X sky130_fd_sc_hd__or2_1
XFILLER_0_122_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14192__B2 _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21439_ hold282/X sstream_i[16] _21442_/S vssd1 vssd1 vccd1 vccd1 _21966_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13269__C _13269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20671__B _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16469__B1 _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12172_ _12169_/X _12172_/B _12175_/A vssd1 vssd1 vccd1 vccd1 _12172_/X sky130_fd_sc_hd__and3b_1
X_11123_ _11123_/A hold1/A vssd1 vssd1 vccd1 vccd1 _11123_/X sky130_fd_sc_hd__or2_1
XFILLER_0_130_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16980_ _16980_/A _16980_/B _16980_/C vssd1 vssd1 vccd1 vccd1 _17028_/A sky130_fd_sc_hd__nand3_1
X_15931_ _15931_/A _15931_/B _16369_/B _16177_/B vssd1 vssd1 vccd1 vccd1 _16056_/A
+ sky130_fd_sc_hd__and4_1
X_11054_ _11053_/X hold86/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21656_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18795__C _19751_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18650_ _19445_/A _19872_/C vssd1 vssd1 vccd1 vccd1 _18653_/A sky130_fd_sc_hd__and2_1
X_15862_ _15862_/A _15862_/B _15862_/C vssd1 vssd1 vccd1 vccd1 _15862_/X sky130_fd_sc_hd__and3_1
XFILLER_0_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17601_ _17602_/A _17602_/B _17602_/C vssd1 vssd1 vccd1 vccd1 _17825_/A sky130_fd_sc_hd__a21oi_2
X_14813_ _14813_/A _15788_/B vssd1 vssd1 vccd1 vccd1 _14814_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_99_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18581_ _18873_/A _19223_/B _18581_/C _18581_/D vssd1 vssd1 vccd1 vccd1 _18582_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_3740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15793_ _16369_/A _16040_/C _15794_/C _15794_/D vssd1 vssd1 vccd1 vccd1 _15795_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__14397__A _14398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14828__C _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17532_ _17532_/A _17532_/B vssd1 vssd1 vccd1 vccd1 _17534_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_153_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14744_ _14584_/A _14584_/B _14582_/Y vssd1 vssd1 vccd1 vccd1 _14746_/B sky130_fd_sc_hd__a21boi_4
XTAP_3784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11956_ _11956_/A _11956_/B vssd1 vssd1 vccd1 vccd1 _12015_/B sky130_fd_sc_hd__xor2_1
XTAP_3795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10907_ _10908_/B vssd1 vssd1 vccd1 vccd1 _10917_/A sky130_fd_sc_hd__inv_2
X_17463_ _17351_/B _17351_/Y _17460_/X _17462_/Y vssd1 vssd1 vccd1 vccd1 _17466_/C
+ sky130_fd_sc_hd__a211oi_4
X_14675_ _15808_/C _16406_/A _14676_/C _14825_/A vssd1 vssd1 vccd1 vccd1 _14677_/B
+ sky130_fd_sc_hd__a22o_1
X_11887_ _11887_/A _11887_/B vssd1 vssd1 vccd1 vccd1 _11889_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19202_ _19202_/A _19202_/B _19348_/B vssd1 vssd1 vccd1 vccd1 _19204_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_67_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16414_ _16414_/A _16414_/B vssd1 vssd1 vccd1 vccd1 _16416_/A sky130_fd_sc_hd__nand2_1
X_13626_ _14087_/A _15098_/B _14557_/D _14089_/A vssd1 vssd1 vccd1 vccd1 _13627_/C
+ sky130_fd_sc_hd__a22o_1
X_10838_ _10836_/B _11055_/A _10817_/Y vssd1 vssd1 vccd1 vccd1 _11057_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_156_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17394_ _17490_/A _17741_/B vssd1 vssd1 vccd1 vccd1 _17398_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13560__A1_N _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19133_ _19133_/A _19133_/B _19133_/C vssd1 vssd1 vccd1 vccd1 _19135_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_55_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16345_ _16345_/A _16345_/B vssd1 vssd1 vccd1 vccd1 _16347_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_55_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13557_ _13557_/A _13557_/B vssd1 vssd1 vccd1 vccd1 _13567_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19894__B1 _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12981__A2 _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19064_ _19064_/A _19064_/B vssd1 vssd1 vccd1 vccd1 _19078_/A sky130_fd_sc_hd__xnor2_1
X_12508_ _12606_/A _12508_/B vssd1 vssd1 vccd1 vccd1 _12522_/A sky130_fd_sc_hd__or2_1
X_16276_ _16277_/A _16277_/B vssd1 vssd1 vccd1 vccd1 _16276_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_125_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13488_ _13338_/B _13338_/Y _13485_/X _13487_/Y vssd1 vssd1 vccd1 vccd1 _13491_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_124_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14183__A1 _14659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18015_ _18014_/B _18014_/C _18014_/A vssd1 vssd1 vccd1 vccd1 _18018_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_23_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15227_ _15218_/A _15080_/B _15215_/B _15085_/C vssd1 vssd1 vccd1 vccd1 _15244_/A
+ sky130_fd_sc_hd__a31o_1
X_12439_ _12331_/X _12333_/X _12436_/X _12437_/Y vssd1 vssd1 vccd1 vccd1 _12439_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_120_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19110__A2 _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15158_ _15156_/X _15158_/B vssd1 vssd1 vccd1 vccd1 _15163_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_2_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14109_ _14132_/B _14109_/B _14107_/X _14108_/Y vssd1 vssd1 vccd1 vccd1 _14109_/X
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_1_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15089_ _14984_/A _14984_/C _14984_/B vssd1 vssd1 vccd1 vccd1 _15103_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_120_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout109 _19692_/C vssd1 vssd1 vccd1 vccd1 _19057_/C sky130_fd_sc_hd__buf_2
XANTENNA__17672__A2 _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19966_ _20101_/B _19866_/D _19874_/B _20101_/A vssd1 vssd1 vccd1 vccd1 _19966_/X
+ sky130_fd_sc_hd__a22o_1
X_18917_ _18917_/A _18917_/B _18917_/C vssd1 vssd1 vccd1 vccd1 _18919_/B sky130_fd_sc_hd__and3_1
XFILLER_0_38_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19897_ _19898_/A _19898_/B _19898_/C vssd1 vssd1 vccd1 vccd1 _19897_/X sky130_fd_sc_hd__a21o_1
X_18848_ _18849_/A _19201_/B _19013_/C _18849_/B vssd1 vssd1 vccd1 vccd1 _18848_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__18621__A1 _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18621__B2 _19092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18779_ _18925_/A _18778_/C _18778_/A vssd1 vssd1 vccd1 vccd1 _18780_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_89_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20810_ _20562_/B _21256_/B hold264/A _21056_/A vssd1 vssd1 vccd1 vccd1 _20814_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11724__A _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21790_ _21963_/CLK _21790_/D vssd1 vssd1 vccd1 vccd1 _21790_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_72_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20741_ _20742_/A _20742_/B _20742_/C vssd1 vssd1 vccd1 vccd1 _20741_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA_fanout153_A _19092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20731__A2 _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13749__A1 _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17411__A _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20672_ _20672_/A _20858_/B vssd1 vssd1 vccd1 vccd1 _20683_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout320_A _21791_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16027__A _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout418_A _21765_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19637__B1 _21384_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14770__A _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21224_ _21275_/B _21222_/Y _21109_/Y _21111_/Y vssd1 vssd1 vccd1 vccd1 _21225_/B
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__12724__A2 _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 hold130/A vssd1 vssd1 vccd1 vccd1 hold130/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20922__D _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold141 hold141/A vssd1 vssd1 vccd1 vccd1 hold141/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19057__B _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold152 hold152/A vssd1 vssd1 vccd1 vccd1 hold152/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__B1 _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold163 hold163/A vssd1 vssd1 vccd1 vccd1 hold163/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold174 hold174/A vssd1 vssd1 vccd1 vccd1 hold174/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 hold185/A vssd1 vssd1 vccd1 vccd1 hold185/X sky130_fd_sc_hd__dlygate4sd3_1
X_21155_ _21841_/Q _21256_/B _21258_/B _21267_/A vssd1 vssd1 vccd1 vccd1 _21155_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12290__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout610 _21718_/Q vssd1 vssd1 vccd1 vccd1 _21723_/D sky130_fd_sc_hd__buf_4
Xhold196 hold196/A vssd1 vssd1 vccd1 vccd1 hold196/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout621 _17146_/A vssd1 vssd1 vccd1 vccd1 _17141_/A sky130_fd_sc_hd__buf_4
X_20106_ _21831_/Q _21832_/Q _20249_/B _20247_/C vssd1 vssd1 vccd1 vccd1 _20251_/A
+ sky130_fd_sc_hd__and4_1
Xfanout632 _21776_/Q vssd1 vssd1 vccd1 vccd1 _14354_/C sky130_fd_sc_hd__buf_4
Xfanout643 _21329_/B1 vssd1 vssd1 vccd1 vccd1 fanout643/X sky130_fd_sc_hd__clkbuf_8
X_21086_ _21086_/A _21086_/B vssd1 vssd1 vccd1 vccd1 _21090_/A sky130_fd_sc_hd__xnor2_2
X_20037_ _19807_/X _19814_/B _19809_/B vssd1 vssd1 vccd1 vccd1 _20039_/B sky130_fd_sc_hd__a21o_1
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout66_A _20841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11810_ _11810_/A _11810_/B _11810_/C vssd1 vssd1 vccd1 vccd1 _11848_/A sky130_fd_sc_hd__nand3_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ _12790_/A _12790_/B _12790_/C vssd1 vssd1 vccd1 vccd1 _12792_/B sky130_fd_sc_hd__nand3_1
XANTENNA__17179__A1 _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21988_ _22020_/CLK _21988_/D vssd1 vssd1 vccd1 vccd1 hold204/A sky130_fd_sc_hd__dfxtp_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _11741_/A _11741_/B _11741_/C vssd1 vssd1 vccd1 vccd1 _11761_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_96_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20939_ _20910_/A _21171_/B _20911_/A _20776_/A vssd1 vssd1 vccd1 vccd1 _20946_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13271__D _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19335__A1_N _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14460_ _14460_/A _14460_/B vssd1 vssd1 vccd1 vccd1 _14462_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_3_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11672_ _11672_/A _11672_/B vssd1 vssd1 vccd1 vccd1 _11805_/A sky130_fd_sc_hd__xor2_1
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13411_ _13411_/A _13411_/B vssd1 vssd1 vccd1 vccd1 _13413_/B sky130_fd_sc_hd__and2_1
XFILLER_0_154_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14391_ _15375_/A _14391_/B _14391_/C _14391_/D vssd1 vssd1 vccd1 vccd1 _14393_/B
+ sky130_fd_sc_hd__nand4_4
XANTENNA__11215__A2 _11126_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20563__A2_N _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16130_ _15999_/A _15999_/Y _16128_/Y _16129_/X vssd1 vssd1 vccd1 vccd1 _16132_/A
+ sky130_fd_sc_hd__o211a_1
X_13342_ _13343_/A _13343_/B _13343_/C _13343_/D vssd1 vssd1 vccd1 vccd1 _13342_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_91_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12963__A2 _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16061_ _16286_/A _16369_/B _16062_/D _16060_/Y vssd1 vssd1 vccd1 vccd1 _16064_/B
+ sky130_fd_sc_hd__a22o_1
X_13273_ _13273_/A _13416_/B _13273_/C vssd1 vssd1 vccd1 vccd1 _13427_/A sky130_fd_sc_hd__or3_2
XFILLER_0_51_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15012_ _15012_/A _15012_/B _15012_/C _15012_/D vssd1 vssd1 vccd1 vccd1 _15012_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__13912__A1 _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12224_ _12224_/A _12224_/B vssd1 vssd1 vccd1 vccd1 _12226_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__13912__B2 _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17103__A1 _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19820_ _19820_/A _19820_/B vssd1 vssd1 vccd1 vccd1 _19828_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17991__A _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12155_ _12229_/A _12155_/B _12269_/C _12269_/D vssd1 vssd1 vccd1 vccd1 _12197_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_20_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16862__B1 _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ _10886_/Y hold73/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21700_/D sky130_fd_sc_hd__mux2_1
X_19751_ _19972_/A _20394_/B _19751_/C _19872_/C vssd1 vssd1 vccd1 vccd1 _19753_/D
+ sky130_fd_sc_hd__nand4_4
X_16963_ _16961_/B _16961_/C _16961_/A vssd1 vssd1 vccd1 vccd1 _16963_/X sky130_fd_sc_hd__a21o_1
X_12086_ _12050_/A _12050_/C _12050_/B vssd1 vssd1 vccd1 vccd1 _12102_/B sky130_fd_sc_hd__a21o_1
X_18702_ _18702_/A _18702_/B vssd1 vssd1 vccd1 vccd1 _18705_/A sky130_fd_sc_hd__xor2_1
X_15914_ _15914_/A _16102_/B vssd1 vssd1 vccd1 vccd1 _15925_/A sky130_fd_sc_hd__nand2_1
X_11037_ mstream_o[111] hold268/X _11039_/S vssd1 vssd1 vccd1 vccd1 _21648_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19682_ _19683_/A _19683_/B vssd1 vssd1 vccd1 vccd1 _19798_/B sky130_fd_sc_hd__and2b_1
X_16894_ _16894_/A _16894_/B vssd1 vssd1 vccd1 vccd1 _16896_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19414__C _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20410__A1 _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18633_ _18472_/Y _18474_/X _18631_/X _18632_/Y vssd1 vssd1 vccd1 vccd1 _18669_/A
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__20410__B2 _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15845_ _15846_/A _15846_/B vssd1 vssd1 vccd1 vccd1 _15847_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_95_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18564_ _18564_/A _18564_/B _18564_/C vssd1 vssd1 vccd1 vccd1 _18564_/X sky130_fd_sc_hd__and3_1
X_15776_ _15776_/A _15776_/B vssd1 vssd1 vccd1 vccd1 _15778_/B sky130_fd_sc_hd__nand2_1
XTAP_3570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12988_ _12988_/A _12988_/B vssd1 vssd1 vccd1 vccd1 _13002_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17515_ _17513_/B _17513_/C _17513_/A vssd1 vssd1 vccd1 vccd1 _17515_/Y sky130_fd_sc_hd__a21oi_2
X_14727_ _15076_/A _15076_/B _15368_/D _15234_/C vssd1 vssd1 vccd1 vccd1 _14854_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_129_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18495_ _18493_/X _18495_/B vssd1 vssd1 vccd1 vccd1 _18496_/B sky130_fd_sc_hd__and2b_1
X_11939_ _11940_/A _11940_/B vssd1 vssd1 vccd1 vccd1 _11960_/B sky130_fd_sc_hd__nand2_1
XANTENNA__19430__B _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13181__D _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13994__A4 _14635_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17446_ _17446_/A _17446_/B vssd1 vssd1 vccd1 vccd1 _17455_/A sky130_fd_sc_hd__xnor2_2
X_14658_ _15653_/C _14657_/X _14656_/X vssd1 vssd1 vccd1 vccd1 _14660_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_89_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13609_ _14848_/A _14873_/B _13470_/B _13468_/X vssd1 vssd1 vccd1 vccd1 _13616_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_83_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17377_ hold134/X _17376_/X fanout3/X vssd1 vssd1 vccd1 vccd1 hold135/A sky130_fd_sc_hd__mux2_1
XFILLER_0_156_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14589_ _14435_/A _14435_/B _14433_/X vssd1 vssd1 vccd1 vccd1 _14591_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19116_ _19587_/B _20242_/D _20249_/B _19587_/A vssd1 vssd1 vccd1 vccd1 _19116_/X
+ sky130_fd_sc_hd__a22o_1
X_16328_ _16328_/A _16328_/B vssd1 vssd1 vccd1 vccd1 _16329_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_125_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14156__A1 _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19047_ _19048_/A _19048_/B vssd1 vssd1 vccd1 vccd1 _19047_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_152_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16259_ hold128/X _16258_/X fanout1/X vssd1 vssd1 vccd1 vccd1 hold129/A sky130_fd_sc_hd__mux2_1
XFILLER_0_112_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11719__A _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19949_ _19841_/A _19838_/X _19839_/Y _19842_/X vssd1 vssd1 vccd1 vccd1 _20070_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13131__A2 _13269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15852__C _16396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15408__A1 _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15408__B2 _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21911_ _21945_/CLK _21911_/D vssd1 vssd1 vccd1 vccd1 hold276/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__11693__A2 _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout270_A _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout368_A _15916_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21842_ _21845_/CLK _21842_/D vssd1 vssd1 vccd1 vccd1 _21842_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_78_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11445__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21773_ _21789_/CLK _21773_/D vssd1 vssd1 vccd1 vccd1 _21773_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_37_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11604__D _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout535_A _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14919__B1 _10912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20724_ _20724_/A _20724_/B vssd1 vssd1 vccd1 vccd1 _20726_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__19570__A2 _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20655_ _20910_/A _21258_/B vssd1 vssd1 vccd1 vccd1 _20656_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20586_ _20721_/D _21291_/B _20586_/C _20586_/D vssd1 vssd1 vccd1 vccd1 _20719_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__17333__A1 _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17333__B2 _17334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19068__A _19692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19086__A1 _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19086__B2 _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21207_ _21207_/A _21207_/B vssd1 vssd1 vccd1 vccd1 _21220_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11629__A _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17019__C _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21138_ _21138_/A _21138_/B vssd1 vssd1 vccd1 vccd1 _21138_/X sky130_fd_sc_hd__or2_1
Xfanout440 _14572_/A vssd1 vssd1 vccd1 vccd1 _12268_/A sky130_fd_sc_hd__buf_4
Xfanout451 _14248_/A vssd1 vssd1 vccd1 vccd1 _14089_/A sky130_fd_sc_hd__buf_4
Xfanout462 _21754_/Q vssd1 vssd1 vccd1 vccd1 _16369_/B sky130_fd_sc_hd__clkbuf_8
Xfanout473 _21751_/Q vssd1 vssd1 vccd1 vccd1 _15091_/C sky130_fd_sc_hd__buf_4
X_13960_ _13960_/A _13960_/B vssd1 vssd1 vccd1 vccd1 _13962_/B sky130_fd_sc_hd__xnor2_2
X_21069_ _21069_/A _21069_/B vssd1 vssd1 vccd1 vccd1 _21069_/Y sky130_fd_sc_hd__nor2_1
Xfanout484 _21748_/Q vssd1 vssd1 vccd1 vccd1 _16326_/A sky130_fd_sc_hd__buf_4
Xfanout495 _21745_/Q vssd1 vssd1 vccd1 vccd1 _14212_/C sky130_fd_sc_hd__buf_4
XANTENNA__14870__A2 _14217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14659__B _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ _14089_/A _14087_/A _14391_/B _13913_/C vssd1 vssd1 vccd1 vccd1 _12913_/B
+ sky130_fd_sc_hd__nand4_1
X_13891_ _13770_/A _13769_/B _13767_/X vssd1 vssd1 vccd1 vccd1 _13906_/A sky130_fd_sc_hd__a21o_1
XANTENNA__20943__A2 _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15630_ _15511_/A _15670_/B _15519_/B _15518_/B _15518_/A vssd1 vssd1 vccd1 vccd1
+ _15645_/A sky130_fd_sc_hd__a32o_2
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19531__A _19531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12842_ _12839_/X _12842_/B _13394_/A _13997_/C vssd1 vssd1 vccd1 vccd1 _12844_/A
+ sky130_fd_sc_hd__and4b_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14083__B1 _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20677__A _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15561_ _15561_/A _15561_/B _15561_/C vssd1 vssd1 vccd1 vccd1 _15561_/X sky130_fd_sc_hd__and3_1
XFILLER_0_96_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ _13018_/B _21766_/Q _12896_/A _12773_/D vssd1 vssd1 vccd1 vccd1 _12896_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_150_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17300_ _17619_/A _17619_/B _17300_/C _17520_/D vssd1 vssd1 vccd1 vccd1 _17393_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_57_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14512_ _14512_/A _14512_/B vssd1 vssd1 vccd1 vccd1 _14526_/A sky130_fd_sc_hd__xnor2_2
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18280_ _18849_/B _19223_/B _18281_/C _18281_/D vssd1 vssd1 vccd1 vccd1 _18282_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ _12784_/A _13155_/B vssd1 vssd1 vccd1 vccd1 _11727_/A sky130_fd_sc_hd__and2_1
X_15492_ _15492_/A _15492_/B vssd1 vssd1 vccd1 vccd1 _15492_/Y sky130_fd_sc_hd__nor2_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12907__B _14712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17231_ _17231_/A _17231_/B vssd1 vssd1 vccd1 vccd1 _17251_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_138_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14443_ _14443_/A _14443_/B vssd1 vssd1 vccd1 vccd1 _14446_/C sky130_fd_sc_hd__xor2_2
X_11655_ _11655_/A _11655_/B vssd1 vssd1 vccd1 vccd1 _11799_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout80 _21847_/Q vssd1 vssd1 vccd1 vccd1 _20606_/D sky130_fd_sc_hd__buf_4
Xfanout91 _21844_/Q vssd1 vssd1 vccd1 vccd1 _21301_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17162_ _17117_/Y _17159_/X _17160_/Y _17161_/X vssd1 vssd1 vccd1 vccd1 _17162_/X
+ sky130_fd_sc_hd__a211o_1
X_14374_ _14373_/A _14373_/B _14373_/C vssd1 vssd1 vccd1 vccd1 _14375_/C sky130_fd_sc_hd__a21o_1
X_11586_ _12319_/C _12511_/A _12402_/A _12420_/D vssd1 vssd1 vccd1 vccd1 _11589_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10947__A1 _10946_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16113_ _16114_/A _16114_/B _16114_/C vssd1 vssd1 vccd1 vccd1 _16113_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__21301__A _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12400__A4 _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13325_ _14089_/A _14087_/A _14234_/C _15370_/B vssd1 vssd1 vccd1 vccd1 _13327_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_134_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17875__A2 _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17093_ _17144_/A _17129_/B _17145_/B _17146_/C vssd1 vssd1 vccd1 vccd1 _17094_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_49_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19409__C _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16044_ _16371_/A _16414_/B _21753_/Q _16380_/A vssd1 vssd1 vccd1 vccd1 _16048_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18313__C _18929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20562__D _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13256_ _14312_/D _13997_/C vssd1 vssd1 vccd1 vccd1 _13257_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13897__B1 _14218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12642__B _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17088__B1 _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12207_ _12207_/A _12207_/B _12207_/C vssd1 vssd1 vccd1 vccd1 _12207_/X sky130_fd_sc_hd__or3_1
X_13187_ _14087_/A _14077_/B _14234_/C _14089_/A vssd1 vssd1 vccd1 vccd1 _13188_/C
+ sky130_fd_sc_hd__a22o_1
X_12138_ _12261_/A _12530_/A _12512_/A _12269_/B vssd1 vssd1 vccd1 vccd1 _12139_/C
+ sky130_fd_sc_hd__a22o_1
X_19803_ _20032_/D _20841_/B _19804_/C _19804_/D vssd1 vssd1 vccd1 vccd1 _19808_/A
+ sky130_fd_sc_hd__a22o_1
X_17995_ _17995_/A _17995_/B vssd1 vssd1 vccd1 vccd1 _18005_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16946_ _16946_/A _16946_/B _16946_/C vssd1 vssd1 vccd1 vccd1 _16946_/X sky130_fd_sc_hd__or3_1
X_12069_ _12063_/A _12063_/B _12056_/X vssd1 vssd1 vccd1 vccd1 _12073_/A sky130_fd_sc_hd__a21o_1
X_19734_ _20088_/A _20242_/D _19734_/C _19849_/A vssd1 vssd1 vccd1 vccd1 _19849_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__12321__B1 _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13473__B _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19665_ _20026_/B _20193_/D _19666_/C _19820_/A vssd1 vssd1 vccd1 vccd1 _19667_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16877_ _17096_/A _17013_/D _16867_/X _16868_/X _17013_/C vssd1 vssd1 vccd1 vccd1
+ _16881_/A sky130_fd_sc_hd__a32o_1
XANTENNA__11675__A2 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20395__B1 _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18616_ _19535_/A _19695_/A _18929_/B _18616_/D vssd1 vssd1 vccd1 vccd1 _18617_/A
+ sky130_fd_sc_hd__and4_1
X_15828_ _16087_/A _15829_/C _16084_/D _15695_/A vssd1 vssd1 vccd1 vccd1 _15832_/C
+ sky130_fd_sc_hd__a22o_1
X_19596_ _19444_/A _19847_/A _19591_/X _19593_/Y vssd1 vssd1 vccd1 vccd1 _19597_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12089__B _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18547_ _18703_/A _19181_/B vssd1 vssd1 vccd1 vccd1 _18548_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15759_ fanout9/A _21404_/B vssd1 vssd1 vccd1 vccd1 _15759_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_87_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18478_ _18478_/A _18478_/B _18478_/C vssd1 vssd1 vccd1 vccd1 _18478_/X sky130_fd_sc_hd__or3_1
XFILLER_0_51_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17429_ _17312_/X _17314_/X _17426_/X _17427_/Y vssd1 vssd1 vccd1 vccd1 _17429_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_7_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11213__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20440_ _20440_/A _20440_/B _20440_/C vssd1 vssd1 vccd1 vccd1 _20441_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_71_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17505__A2_N _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11060__A0 _11059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21211__A _21311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20371_ _20513_/A _20371_/B vssd1 vssd1 vccd1 vccd1 _20643_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16305__A _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout116_A _21839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22041_ _22049_/CLK _22041_/D vssd1 vssd1 vccd1 vccd1 hold238/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout485_A _21748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16040__A _16391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14479__B _15174_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16975__A _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19351__A _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21825_ _21829_/CLK _21825_/D vssd1 vssd1 vccd1 vccd1 _21825_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__19070__B _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11912__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21756_ _22063_/CLK _21756_/D vssd1 vssd1 vccd1 vccd1 hold320/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21350__A2 _17834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout29_A _11124_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20707_ _20707_/A _20707_/B _20707_/C vssd1 vssd1 vccd1 vccd1 _20708_/C sky130_fd_sc_hd__and3_1
XFILLER_0_148_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21687_ _22069_/CLK _21687_/D vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20944__B _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11440_ _11439_/X _21256_/B _11470_/S vssd1 vssd1 vccd1 vccd1 _21818_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_135_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20638_ _20638_/A _20638_/B vssd1 vssd1 vccd1 vccd1 _20903_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16860__D _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11371_ _11370_/X _17063_/C _11401_/S vssd1 vssd1 vccd1 vccd1 _21795_/D sky130_fd_sc_hd__mux2_1
X_20569_ _20569_/A _20569_/B vssd1 vssd1 vccd1 vccd1 _20571_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__16215__A _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13110_ _13111_/A _13111_/B vssd1 vssd1 vccd1 vccd1 _13110_/Y sky130_fd_sc_hd__nor2_1
X_14090_ _14090_/A _14090_/B _14090_/C vssd1 vssd1 vccd1 vccd1 _14093_/A sky130_fd_sc_hd__or3_1
X_13041_ _13040_/B _13040_/C _13040_/A vssd1 vssd1 vccd1 vccd1 _13042_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__18787__D _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16800_ _16800_/A _16800_/B _16800_/C vssd1 vssd1 vccd1 vccd1 _16806_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_79_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17780_ _20583_/A _18789_/A _17913_/A _17780_/D vssd1 vssd1 vccd1 vccd1 _17913_/B
+ sky130_fd_sc_hd__nand4_2
X_14992_ _15632_/B _16268_/B _16266_/C _14993_/A vssd1 vssd1 vccd1 vccd1 _14994_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout270 _19664_/B vssd1 vssd1 vccd1 vccd1 _19051_/A sky130_fd_sc_hd__buf_4
XANTENNA__14389__B _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout281 _18008_/B vssd1 vssd1 vccd1 vccd1 _19644_/A sky130_fd_sc_hd__buf_4
X_16731_ _16730_/A _16730_/C _16730_/B vssd1 vssd1 vccd1 vccd1 _16738_/B sky130_fd_sc_hd__a21o_1
Xfanout292 _21797_/Q vssd1 vssd1 vccd1 vccd1 _17874_/A sky130_fd_sc_hd__buf_8
X_13943_ _13943_/A _13943_/B _13941_/X _13942_/Y vssd1 vssd1 vccd1 vccd1 _13943_/X
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_89_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18034__A2 _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11657__A2 _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19450_ _19296_/A _19296_/B _19294_/Y vssd1 vssd1 vccd1 vccd1 _19452_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_88_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16662_ _16662_/A _16662_/B _16662_/C vssd1 vssd1 vccd1 vccd1 _16694_/A sky130_fd_sc_hd__nand3_1
X_13874_ _21741_/Q _14516_/A _14365_/C _13875_/B vssd1 vssd1 vccd1 vccd1 _13877_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17793__A1 _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18401_ _18420_/B vssd1 vssd1 vccd1 vccd1 _18550_/A sky130_fd_sc_hd__inv_2
XFILLER_0_9_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15613_ _15612_/A _15612_/B _15612_/C _15612_/D vssd1 vssd1 vccd1 vccd1 _15613_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__20838__C _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19381_ _19382_/A _20419_/A _19382_/C _19382_/D vssd1 vssd1 vccd1 vccd1 _19381_/X
+ sky130_fd_sc_hd__and4_1
X_12825_ _12825_/A _12825_/B _12825_/C vssd1 vssd1 vccd1 vccd1 _12825_/X sky130_fd_sc_hd__or3_1
XANTENNA__21087__A_N _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16593_ _17526_/B _16813_/A _16743_/B _17525_/A vssd1 vssd1 vccd1 vccd1 _16594_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18332_ _18332_/A _18332_/B vssd1 vssd1 vccd1 vccd1 _18343_/A sky130_fd_sc_hd__or2_1
XFILLER_0_57_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15544_ _15545_/A _15545_/B vssd1 vssd1 vccd1 vccd1 _15727_/B sky130_fd_sc_hd__or2_1
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12756_ _14024_/B _13013_/A _13155_/D vssd1 vssd1 vccd1 vccd1 _12756_/X sky130_fd_sc_hd__and3_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17545__A1 _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21341__A2 _17484_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12637__B _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18263_ _18263_/A _18263_/B vssd1 vssd1 vccd1 vccd1 _18265_/B sky130_fd_sc_hd__xnor2_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11707_ _12267_/A _13017_/A _12444_/B _12094_/B vssd1 vssd1 vccd1 vccd1 _11707_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_72_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15475_ _15475_/A _15475_/B _15475_/C _15475_/D vssd1 vssd1 vccd1 vccd1 _15475_/Y
+ sky130_fd_sc_hd__nand4_4
XANTENNA__18850__A2_N _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12687_ _12687_/A _12687_/B _12687_/C vssd1 vssd1 vccd1 vccd1 _12687_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_155_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17214_ _17215_/A _17215_/B vssd1 vssd1 vccd1 vccd1 _17214_/X sky130_fd_sc_hd__and2_1
XFILLER_0_126_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14426_ _14426_/A _14426_/B vssd1 vssd1 vccd1 vccd1 _14427_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_115_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18194_ _18195_/A _18195_/B vssd1 vssd1 vccd1 vccd1 _18328_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11638_ _12528_/B _12020_/A _13155_/D _12619_/A vssd1 vssd1 vccd1 vccd1 _11640_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17145_ _17145_/A _17145_/B vssd1 vssd1 vccd1 vccd1 _17145_/X sky130_fd_sc_hd__or2_1
XFILLER_0_123_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14357_ _14813_/A _16369_/A _14357_/C _14357_/D vssd1 vssd1 vccd1 vccd1 _14357_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_107_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11569_ _12109_/C _13556_/A vssd1 vssd1 vccd1 vccd1 _11865_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13308_ _13308_/A _13308_/B vssd1 vssd1 vccd1 vccd1 _13318_/A sky130_fd_sc_hd__or2_2
XANTENNA__13468__B _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17076_ _17073_/A _17073_/B _17073_/C vssd1 vssd1 vccd1 vccd1 _17078_/C sky130_fd_sc_hd__a21oi_1
X_14288_ _14288_/A _14288_/B vssd1 vssd1 vccd1 vccd1 _14601_/C sky130_fd_sc_hd__and2_2
XANTENNA_clkbuf_leaf_40_clk_i_A _21822_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16027_ _16027_/A _16027_/B vssd1 vssd1 vccd1 vccd1 _16028_/B sky130_fd_sc_hd__nand2_1
X_13239_ _13237_/Y _13239_/B vssd1 vssd1 vccd1 vccd1 _13240_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_62_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11345__B2 _11089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20604__A1 _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20604__B2 _21261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17978_ _17978_/A _18117_/A vssd1 vssd1 vccd1 vccd1 _17980_/C sky130_fd_sc_hd__nor2_1
XANTENNA__13098__B2 _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16929_ _16923_/A _16923_/C _16923_/B vssd1 vssd1 vccd1 vccd1 _16930_/C sky130_fd_sc_hd__a21o_1
XANTENNA__19222__A1 _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19717_ _19580_/X _19585_/A _19715_/Y _19716_/X vssd1 vssd1 vccd1 vccd1 _19719_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__16795__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17233__B1 _17443_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19648_ _20838_/C _19487_/X _19490_/A _19490_/B vssd1 vssd1 vccd1 vccd1 _19649_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19579_ _19578_/B _19578_/C _19578_/A vssd1 vssd1 vccd1 vccd1 _19581_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12828__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21610_ _21906_/CLK _21610_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[73] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_133_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13270__A1 _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13270__B2 _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21332__A2 _17173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21541_ mstream_o[4] hold4/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22068_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_29_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout233_A _17924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21472_ hold184/X sstream_i[49] _21481_/S vssd1 vssd1 vccd1 vccd1 _21999_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_117_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20423_ _20423_/A _20423_/B vssd1 vssd1 vccd1 vccd1 _20425_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_114_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout400_A _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11584__A1 _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20354_ _20354_/A _20354_/B vssd1 vssd1 vccd1 vccd1 _20354_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20285_ _20689_/A _20562_/B _21153_/B _21264_/B vssd1 vssd1 vccd1 vccd1 _20427_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__11336__A1 _11335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17792__C _18789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22024_ _22038_/CLK _22024_/D vssd1 vssd1 vccd1 vccd1 hold316/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__16689__B _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15593__B _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15078__A2 _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13394__A _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13711__A2_N _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18400__D _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20004__B _20562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 hold67/A vssd1 vssd1 vccd1 vccd1 hold67/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 hold78/A vssd1 vssd1 vccd1 vccd1 hold78/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 hold89/A vssd1 vssd1 vccd1 vccd1 hold89/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10940_ _10940_/A _10940_/B _10938_/Y vssd1 vssd1 vccd1 vccd1 _10941_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_39_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10871_ _10871_/A _10880_/A vssd1 vssd1 vccd1 vccd1 _10873_/C sky130_fd_sc_hd__or2_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ _13983_/B _14018_/C _12610_/C _12610_/D vssd1 vssd1 vccd1 vccd1 _12728_/B
+ sky130_fd_sc_hd__and4_1
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21808_ _21809_/CLK _21808_/D vssd1 vssd1 vccd1 vccd1 _21808_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13590_ _13875_/B _14537_/A _13591_/C _13591_/D vssd1 vssd1 vccd1 vccd1 _13592_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13261__A1 _13554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17527__A1 _21802_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17527__B2 _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11272__A0 _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12457__B _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12541_ _12542_/A _12542_/B vssd1 vssd1 vccd1 vccd1 _12541_/X sky130_fd_sc_hd__and2_2
XFILLER_0_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21739_ _21803_/CLK _21739_/D vssd1 vssd1 vccd1 vccd1 _21739_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20674__B _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15260_ _16371_/A _16305_/B _16399_/A _15791_/A vssd1 vssd1 vccd1 vccd1 _15264_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12472_ _12471_/B _12471_/C _12471_/A vssd1 vssd1 vccd1 vccd1 _12472_/Y sky130_fd_sc_hd__a21oi_2
X_14211_ _14212_/B _14212_/C _14212_/D _14384_/A vssd1 vssd1 vccd1 vccd1 _14213_/A
+ sky130_fd_sc_hd__a22o_1
X_11423_ _21718_/D hold291/A fanout47/X hold164/A vssd1 vssd1 vccd1 vccd1 _11423_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15191_ _15346_/B _15191_/B vssd1 vssd1 vccd1 vccd1 _15192_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_105_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14761__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_9 _11331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12772__B1 _21765_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14142_ _14142_/A _14142_/B vssd1 vssd1 vccd1 vccd1 _14144_/B sky130_fd_sc_hd__or2_1
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11354_ _11124_/A hold225/A _11126_/B hold160/X vssd1 vssd1 vccd1 vccd1 _11354_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11089__A _11089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14073_ _14073_/A _14073_/B vssd1 vssd1 vccd1 vccd1 _14081_/A sky130_fd_sc_hd__nand2_1
X_11285_ _11325_/A1 t2y[15] t0y[15] _11498_/A1 vssd1 vssd1 vccd1 vccd1 _11285_/X sky130_fd_sc_hd__a22o_1
X_18950_ _19951_/B _19866_/C _18951_/C _19106_/A vssd1 vssd1 vccd1 vccd1 _18950_/X
+ sky130_fd_sc_hd__a22o_1
X_13024_ _13023_/A _13023_/B _13023_/C vssd1 vssd1 vccd1 vccd1 _13025_/C sky130_fd_sc_hd__a21o_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17901_ _17901_/A _17901_/B _17901_/C vssd1 vssd1 vccd1 vccd1 _17904_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_30_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18255__A2 _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18881_ _18881_/A vssd1 vssd1 vccd1 vccd1 _18881_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_20_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17832_ _17832_/A _17832_/B vssd1 vssd1 vccd1 vccd1 _21349_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__18007__A2 _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17763_ _19892_/A _19823_/A _18319_/B _18622_/B vssd1 vssd1 vccd1 vccd1 _17765_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_156_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14975_ _15085_/A _15502_/A vssd1 vssd1 vccd1 vccd1 _15363_/A sky130_fd_sc_hd__nor2_2
XANTENNA__19703__B _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16714_ _16708_/Y _16711_/X _16713_/Y _16682_/X vssd1 vssd1 vccd1 vccd1 _16718_/A
+ sky130_fd_sc_hd__o211ai_4
X_19502_ _19502_/A _19502_/B vssd1 vssd1 vccd1 vccd1 _19522_/A sky130_fd_sc_hd__or2_1
X_13926_ _14087_/A _15234_/C _14250_/B _14248_/A vssd1 vssd1 vccd1 vccd1 _13928_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17694_ _17718_/B _17694_/B _17693_/C _17693_/D vssd1 vssd1 vccd1 vccd1 _17694_/X
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_16_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18319__B _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19433_ _19433_/A _19433_/B _19598_/B vssd1 vssd1 vccd1 vccd1 _19433_/X sky130_fd_sc_hd__and3_1
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16645_ _16645_/A _16645_/B _16645_/C vssd1 vssd1 vccd1 vccd1 _16672_/A sky130_fd_sc_hd__nand3_2
X_13857_ _13858_/A _13858_/C _16414_/A _13858_/B vssd1 vssd1 vccd1 vccd1 _13859_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_16_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17223__B _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13236__A1_N _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19364_ _19365_/A _19365_/B vssd1 vssd1 vccd1 vccd1 _19364_/Y sky130_fd_sc_hd__nor2_1
X_12808_ _12837_/B _12808_/B _12807_/C _12807_/D vssd1 vssd1 vccd1 vccd1 _12808_/X
+ sky130_fd_sc_hd__or4bb_2
X_16576_ _17206_/B _17619_/B _17211_/A _16575_/D vssd1 vssd1 vccd1 vccd1 _16578_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13788_ _13787_/A _13787_/B _13787_/C vssd1 vssd1 vccd1 vccd1 _13790_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_96_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18315_ _19529_/B _18769_/B _18314_/C _18314_/D vssd1 vssd1 vccd1 vccd1 _18316_/B
+ sky130_fd_sc_hd__a22o_1
X_15527_ _15365_/A _15364_/Y _15386_/X vssd1 vssd1 vccd1 vccd1 _15529_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11263__B1 _11262_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19295_ _19295_/A _19295_/B vssd1 vssd1 vccd1 vccd1 _19296_/B sky130_fd_sc_hd__xor2_2
X_12739_ _12868_/A _12739_/B vssd1 vssd1 vccd1 vccd1 _12741_/B sky130_fd_sc_hd__and2_1
XFILLER_0_155_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18335__A _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18246_ hold190/A fanout8/X _13369_/B _21142_/A vssd1 vssd1 vccd1 vccd1 _18246_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_155_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15458_ _15459_/B _15459_/A vssd1 vssd1 vccd1 vccd1 _15458_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_964 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14409_ _14409_/A _14409_/B _14554_/B vssd1 vssd1 vccd1 vccd1 _14409_/X sky130_fd_sc_hd__and3_1
XANTENNA__13555__A2 _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18177_ _18177_/A _18177_/B vssd1 vssd1 vccd1 vccd1 _18179_/B sky130_fd_sc_hd__xnor2_1
X_15389_ _16196_/B _15911_/A _15911_/C _15717_/B vssd1 vssd1 vccd1 vccd1 _15392_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17128_ _17144_/A _17146_/C _17146_/D _17129_/B vssd1 vssd1 vccd1 vccd1 _17130_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__17893__B _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18494__A2 _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17059_ _17074_/A _17074_/B vssd1 vssd1 vccd1 vccd1 _17081_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_110_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11318__A1 _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20070_ _20070_/A _20070_/B vssd1 vssd1 vccd1 vccd1 _20072_/C sky130_fd_sc_hd__xnor2_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21250__A1 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19994__A2 _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout183_A _17666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20972_ _20973_/B _20972_/B vssd1 vssd1 vccd1 vccd1 _20974_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_36_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20478__C _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout350_A _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21524_ hold247/X sstream_i[101] _21536_/S vssd1 vssd1 vccd1 vccd1 _22051_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_35_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21455_ hold160/X sstream_i[32] _21489_/S vssd1 vssd1 vccd1 vccd1 _21982_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_105_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11401__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20406_ _20407_/A _20407_/B vssd1 vssd1 vccd1 vccd1 _20408_/A sky130_fd_sc_hd__or2_1
XANTENNA__20286__A2_N _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21386_ hold169/X _21381_/B _21384_/X _21385_/Y vssd1 vssd1 vccd1 vccd1 _21936_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18485__A2 _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15299__A2 _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20337_ _20338_/B _20338_/A vssd1 vssd1 vccd1 vccd1 _20337_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__11309__B2 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19507__C _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout96_A _21843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ _10867_/X hold99/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21665_/D sky130_fd_sc_hd__mux2_1
X_20268_ _20268_/A _20473_/B vssd1 vssd1 vccd1 vccd1 _20279_/A sky130_fd_sc_hd__nand2_1
X_22007_ _22013_/CLK _22007_/D vssd1 vssd1 vccd1 vccd1 hold207/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__19226__D _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11637__A _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20199_ _20200_/A _20200_/B vssd1 vssd1 vccd1 vccd1 _20199_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__19198__B1 _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20669__B _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17324__A _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14760_ fanout9/X _19636_/B vssd1 vssd1 vccd1 vccd1 _14760_/Y sky130_fd_sc_hd__nor2_1
X_11972_ _11901_/A _11901_/B _11901_/C vssd1 vssd1 vccd1 vccd1 _11972_/Y sky130_fd_sc_hd__a21oi_1
X_13711_ _13858_/A _16273_/A _13709_/Y _13710_/X vssd1 vssd1 vccd1 vccd1 _13713_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__20388__C _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13571__B _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10923_ _10923_/A _10923_/B vssd1 vssd1 vccd1 vccd1 _10926_/A sky130_fd_sc_hd__nand2_2
X_14691_ _14563_/A _14562_/B _14560_/X vssd1 vssd1 vccd1 vccd1 _14707_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_6_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16430_ _16430_/A _16430_/B vssd1 vssd1 vccd1 vccd1 _16431_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_116_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13642_ _13643_/A _13643_/B _13643_/C _13643_/D vssd1 vssd1 vccd1 vccd1 _13642_/Y
+ sky130_fd_sc_hd__nor4_2
X_10854_ hold29/A hold22/A vssd1 vssd1 vccd1 vccd1 _10857_/A sky130_fd_sc_hd__or2_1
XFILLER_0_39_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16882__B _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15779__A _16036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16361_ _16366_/B _16361_/B vssd1 vssd1 vccd1 vccd1 _16362_/B sky130_fd_sc_hd__nor2_1
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ _13570_/Y _13720_/A _13864_/B _13573_/D vssd1 vssd1 vccd1 vccd1 _13720_/B
+ sky130_fd_sc_hd__and4bb_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18100_ _18100_/A _18100_/B vssd1 vssd1 vccd1 vccd1 _18243_/B sky130_fd_sc_hd__xnor2_2
X_15312_ _15156_/X _15162_/A _15162_/B _15158_/B vssd1 vssd1 vccd1 vccd1 _15314_/B
+ sky130_fd_sc_hd__o31ai_2
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19080_ _18944_/B _18946_/A _19078_/X _19079_/Y vssd1 vssd1 vccd1 vccd1 _19082_/A
+ sky130_fd_sc_hd__a211o_1
X_12524_ _12436_/X _12439_/Y _12522_/Y _12523_/X vssd1 vssd1 vccd1 vccd1 _12604_/A
+ sky130_fd_sc_hd__a211oi_2
X_16292_ _16293_/A _16293_/B vssd1 vssd1 vccd1 vccd1 _16294_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_137_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18031_ _18031_/A _18031_/B vssd1 vssd1 vccd1 vccd1 _18032_/B sky130_fd_sc_hd__nand2_1
X_15243_ _15244_/A _15244_/B vssd1 vssd1 vccd1 vccd1 _15243_/X sky130_fd_sc_hd__and2_2
XANTENNA__17994__A _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12455_ _12455_/A _12455_/B vssd1 vssd1 vccd1 vccd1 _12456_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_35_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11406_ hold311/A fanout28/X _11405_/X vssd1 vssd1 vccd1 vccd1 _11406_/X sky130_fd_sc_hd__a21o_1
X_15174_ _15171_/Y _15316_/A _15702_/D _15174_/D vssd1 vssd1 vccd1 vccd1 _15316_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_105_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12386_ _12383_/Y _12384_/X _11840_/A _11839_/Y vssd1 vssd1 vccd1 vccd1 _12387_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14125_ _14291_/B _14291_/C vssd1 vssd1 vccd1 vccd1 _14126_/B sky130_fd_sc_hd__or2_2
XANTENNA__12353__D _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20283__A2 _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11337_ _11349_/A1 t2y[28] t0y[28] _21723_/D vssd1 vssd1 vccd1 vccd1 _11337_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19982_ _20126_/A _19980_/Y _19877_/B _19879_/B vssd1 vssd1 vccd1 vccd1 _19984_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14498__B1 _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14056_ _14212_/C _14055_/X _14054_/X vssd1 vssd1 vccd1 vccd1 _14057_/B sky130_fd_sc_hd__a21bo_1
X_18933_ _19092_/A _19092_/C _19262_/C _20088_/A vssd1 vssd1 vccd1 vccd1 _18936_/B
+ sky130_fd_sc_hd__a22o_1
X_11268_ _12326_/D _11267_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21768_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_120_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13007_ _12866_/Y _12869_/X _13097_/A _13006_/Y vssd1 vssd1 vccd1 vccd1 _13097_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__11547__A _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11199_ hold296/X fanout51/X fanout48/X hold271/A vssd1 vssd1 vccd1 vccd1 _11199_/X
+ sky130_fd_sc_hd__a22o_1
X_18864_ _19024_/B _18864_/B vssd1 vssd1 vccd1 vccd1 _18866_/C sky130_fd_sc_hd__nand2_1
XANTENNA__11720__A1 _13018_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11720__B2 _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17815_ _17852_/B _17815_/B _17815_/C _17815_/D vssd1 vssd1 vccd1 vccd1 _17815_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_0_20_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18795_ _19587_/A _19587_/B _19751_/C _20242_/C vssd1 vssd1 vccd1 vccd1 _18795_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_118_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_89_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17746_ _17746_/A _17746_/B vssd1 vssd1 vccd1 vccd1 _17749_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__17234__A _17334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14958_ _14793_/B _14795_/B _14956_/X _14957_/Y vssd1 vssd1 vccd1 vccd1 _14958_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_27_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13909_ _13906_/X _13907_/Y _13753_/Y _13755_/X vssd1 vssd1 vccd1 vccd1 _13943_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17677_ _17676_/A _17676_/B _17676_/C vssd1 vssd1 vccd1 vccd1 _17678_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_49_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14889_ _14889_/A _14889_/B vssd1 vssd1 vccd1 vccd1 _14892_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_134_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16628_ _16628_/A _16628_/B vssd1 vssd1 vccd1 vccd1 _16629_/C sky130_fd_sc_hd__nor2_1
X_19416_ _20650_/A _19868_/B _19417_/C _19417_/D vssd1 vssd1 vccd1 vccd1 _19416_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_147_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12097__B _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11236__A0 _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16559_ _16813_/A _17223_/A _16860_/C _16743_/B vssd1 vssd1 vccd1 vccd1 _16561_/C
+ sky130_fd_sc_hd__a22o_1
X_19347_ _19234_/A _19233_/B _19231_/X vssd1 vssd1 vccd1 vccd1 _19347_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19278_ _19951_/B _19751_/C _20242_/C _19430_/A vssd1 vssd1 vccd1 vccd1 _19281_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11251__A3 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13528__A2 _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18229_ _18230_/A _18230_/B _18230_/C vssd1 vssd1 vccd1 vccd1 _18229_/X sky130_fd_sc_hd__and3_1
XFILLER_0_4_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11539__A1 _19181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21240_ _21240_/A _21240_/B vssd1 vssd1 vccd1 vccd1 _21241_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold301 hold301/A vssd1 vssd1 vccd1 vccd1 hold301/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold312 hold312/A vssd1 vssd1 vccd1 vccd1 hold312/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold323 hold323/A vssd1 vssd1 vccd1 vccd1 hold323/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21171_ _21171_/A _21171_/B _21171_/C _21171_/D vssd1 vssd1 vccd1 vccd1 _21172_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_141_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20122_ _19984_/A _20122_/B vssd1 vssd1 vccd1 vccd1 _20124_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__19416__A1 _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12560__B _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20053_ _20053_/A _20186_/B _20053_/C vssd1 vssd1 vccd1 vccd1 _20053_/X sky130_fd_sc_hd__and3_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14768__A _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17144__A _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_207 hold270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_218 hold277/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_229 hold290/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20955_ _20784_/A _20785_/Y _20953_/A _20954_/Y vssd1 vssd1 vccd1 vccd1 _20955_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_36_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13822__D _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20886_ _20755_/A _20755_/Y _21016_/B _20885_/Y vssd1 vssd1 vccd1 vccd1 _20886_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_36_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11227__B1 _11226_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12975__B1 _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18406__C _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout11_A _11446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21507_ hold235/X sstream_i[84] _21507_/S vssd1 vssd1 vccd1 vccd1 _22034_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18703__A _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12454__C _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12240_ _12234_/A _12234_/C _12234_/B vssd1 vssd1 vccd1 vccd1 _12241_/B sky130_fd_sc_hd__o21a_1
XANTENNA__14192__A2 _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21438_ hold265/X sstream_i[15] _21442_/S vssd1 vssd1 vccd1 vccd1 _21965_/D sky130_fd_sc_hd__mux2_1
XANTENNA__16469__A1 _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16469__B2 _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12171_ _12169_/X _12172_/B vssd1 vssd1 vccd1 vccd1 _12175_/B sky130_fd_sc_hd__nand2b_1
X_21369_ hold150/X fanout40/X _21367_/X _21368_/Y vssd1 vssd1 vccd1 vccd1 _21930_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12751__A _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11122_ _11122_/A _21724_/D vssd1 vssd1 vccd1 vccd1 _11122_/X sky130_fd_sc_hd__or2_2
XFILLER_0_120_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15930_ _15933_/D vssd1 vssd1 vccd1 vccd1 _15930_/Y sky130_fd_sc_hd__inv_2
X_11053_ _11053_/A _11053_/B vssd1 vssd1 vccd1 vccd1 _11053_/X sky130_fd_sc_hd__xor2_4
XANTENNA__19534__A _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15861_ _15862_/A _15862_/B _15862_/C vssd1 vssd1 vccd1 vccd1 _15861_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__18795__D _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17600_ _18859_/A _21151_/A _17500_/A _17497_/X vssd1 vssd1 vccd1 vccd1 _17602_/C
+ sky130_fd_sc_hd__a31oi_2
X_14812_ _15653_/C _14811_/X _14810_/X vssd1 vssd1 vccd1 vccd1 _14814_/A sky130_fd_sc_hd__a21bo_1
X_18580_ _18873_/A _19223_/B _18581_/C _18581_/D vssd1 vssd1 vccd1 vccd1 _18582_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15792_ _15921_/A vssd1 vssd1 vccd1 vccd1 _15794_/D sky130_fd_sc_hd__inv_2
XFILLER_0_99_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17531_ _17532_/A _17532_/B vssd1 vssd1 vccd1 vccd1 _17531_/X sky130_fd_sc_hd__and2_2
XFILLER_0_19_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14743_ _14743_/A _14743_/B vssd1 vssd1 vccd1 vccd1 _14746_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14828__D _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11955_ _12319_/C _12312_/A vssd1 vssd1 vccd1 vccd1 _12015_/A sky130_fd_sc_hd__nand2_1
XTAP_3785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10906_ hold102/A hold126/A vssd1 vssd1 vccd1 vccd1 _10908_/B sky130_fd_sc_hd__nand2_1
X_17462_ _17461_/B _17461_/C _17461_/A vssd1 vssd1 vccd1 vccd1 _17462_/Y sky130_fd_sc_hd__a21oi_2
X_14674_ _16173_/A _14828_/B _16404_/A _16409_/A vssd1 vssd1 vccd1 vccd1 _14825_/A
+ sky130_fd_sc_hd__nand4_2
X_11886_ _11958_/A _11958_/B vssd1 vssd1 vccd1 vccd1 _11886_/X sky130_fd_sc_hd__and2_1
X_16413_ _16413_/A _16413_/B vssd1 vssd1 vccd1 vccd1 _16423_/A sky130_fd_sc_hd__xnor2_1
X_19201_ _19810_/D _19201_/B _19201_/C _19348_/A vssd1 vssd1 vccd1 vccd1 _19348_/B
+ sky130_fd_sc_hd__nand4_2
X_13625_ _14089_/A _14087_/A _15098_/B _14557_/D vssd1 vssd1 vccd1 vccd1 _13627_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_73_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10837_ _11053_/A _11053_/B _11055_/B vssd1 vssd1 vccd1 vccd1 _10837_/X sky130_fd_sc_hd__or3b_1
X_17393_ _17393_/A _17393_/B vssd1 vssd1 vccd1 vccd1 _17400_/A sky130_fd_sc_hd__or2_1
XFILLER_0_39_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19132_ _18969_/A _18969_/C _18969_/B vssd1 vssd1 vccd1 vccd1 _19133_/C sky130_fd_sc_hd__a21bo_1
X_16344_ _16344_/A _16344_/B vssd1 vssd1 vccd1 vccd1 _16345_/B sky130_fd_sc_hd__xor2_1
X_13556_ _13556_/A _13997_/C _13556_/C _13556_/D vssd1 vssd1 vccd1 vccd1 _13557_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__21150__B1 _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19894__A1 _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19894__B2 _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19063_ _19061_/X _19063_/B vssd1 vssd1 vccd1 vccd1 _19064_/B sky130_fd_sc_hd__nand2b_1
X_12507_ _12605_/A _12605_/B vssd1 vssd1 vccd1 vccd1 _12508_/B sky130_fd_sc_hd__and2_1
X_16275_ _16275_/A _16275_/B vssd1 vssd1 vccd1 vccd1 _16277_/B sky130_fd_sc_hd__or2_1
XFILLER_0_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13487_ _13486_/B _13486_/C _13486_/A vssd1 vssd1 vccd1 vccd1 _13487_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_54_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18014_ _18014_/A _18014_/B _18014_/C vssd1 vssd1 vccd1 vccd1 _18018_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12718__B1 _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15226_ _15226_/A _15226_/B vssd1 vssd1 vccd1 vccd1 _15247_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_35_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12438_ _12331_/X _12333_/X _12436_/X _12437_/Y vssd1 vssd1 vccd1 vccd1 _12475_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15157_ _14930_/D _14934_/B _15154_/X _15305_/B vssd1 vssd1 vccd1 vccd1 _15158_/B
+ sky130_fd_sc_hd__a211o_1
X_12369_ _12370_/A _12370_/B _12370_/C vssd1 vssd1 vccd1 vccd1 _12369_/X sky130_fd_sc_hd__and3_1
XANTENNA__15675__C _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14108_ _14105_/Y _14106_/X _13941_/X _13943_/X vssd1 vssd1 vccd1 vccd1 _14108_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__18051__C _19692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15088_ _15087_/A _15223_/B _15087_/C vssd1 vssd1 vccd1 vccd1 _15108_/B sky130_fd_sc_hd__a21oi_1
X_19965_ _19857_/A _19857_/C _19857_/B vssd1 vssd1 vccd1 vccd1 _19979_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14039_ _14038_/B _14190_/B _14038_/A vssd1 vssd1 vccd1 vccd1 _14040_/C sky130_fd_sc_hd__a21o_1
X_18916_ _18755_/A _18754_/B _18752_/X vssd1 vssd1 vccd1 vccd1 _18917_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11708__C _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19896_ _21199_/A _20419_/A vssd1 vssd1 vccd1 vccd1 _19898_/C sky130_fd_sc_hd__and2_1
XANTENNA__21625__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18847_ _18847_/A _18847_/B vssd1 vssd1 vccd1 vccd1 _18889_/A sky130_fd_sc_hd__or2_1
XANTENNA__18621__A2 _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18778_ _18778_/A _18925_/A _18778_/C vssd1 vssd1 vccd1 vccd1 _18925_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_59_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17729_ _17865_/A _17729_/B _18851_/C _19060_/B vssd1 vssd1 vccd1 vccd1 _17865_/B
+ sky130_fd_sc_hd__and4b_1
XANTENNA__17899__A _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11724__B _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11216__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20740_ _20740_/A _20740_/B vssd1 vssd1 vccd1 vccd1 _20742_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13749__A2 _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20671_ _21296_/A _20671_/B _20671_/C _20858_/A vssd1 vssd1 vccd1 vccd1 _20858_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__17411__B _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout146_A _21832_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout313_A _17141_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19637__B2 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14770__B _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21223_ _21109_/Y _21111_/Y _21275_/B _21222_/Y vssd1 vssd1 vccd1 vccd1 _21225_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold120 hold120/A vssd1 vssd1 vccd1 vccd1 hold120/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 hold131/A vssd1 vssd1 vccd1 vccd1 hold131/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold142 hold142/A vssd1 vssd1 vccd1 vccd1 hold142/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__A1 _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold153 hold153/A vssd1 vssd1 vccd1 vccd1 hold153/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11932__B2 _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21154_ _21154_/A _21154_/B vssd1 vssd1 vccd1 vccd1 _21163_/A sky130_fd_sc_hd__xnor2_1
Xhold164 hold164/A vssd1 vssd1 vccd1 vccd1 hold164/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold175 hold175/A vssd1 vssd1 vccd1 vccd1 hold175/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 hold186/A vssd1 vssd1 vccd1 vccd1 hold186/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12290__B _17173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout600 _21720_/Q vssd1 vssd1 vccd1 vccd1 _16363_/A sky130_fd_sc_hd__clkbuf_8
Xhold197 hold197/A vssd1 vssd1 vccd1 vccd1 hold197/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout611 _21718_/Q vssd1 vssd1 vccd1 vccd1 _11089_/B sky130_fd_sc_hd__clkbuf_4
X_20105_ _21832_/Q _20249_/B _20247_/C _21831_/Q vssd1 vssd1 vccd1 vccd1 _20105_/Y
+ sky130_fd_sc_hd__a22oi_1
Xfanout622 _21822_/Q vssd1 vssd1 vccd1 vccd1 _17146_/A sky130_fd_sc_hd__buf_4
Xfanout633 _21776_/Q vssd1 vssd1 vccd1 vccd1 _14817_/C sky130_fd_sc_hd__buf_2
X_21085_ _21085_/A _21085_/B vssd1 vssd1 vccd1 vccd1 _21086_/B sky130_fd_sc_hd__nor2_2
Xfanout644 _21329_/B1 vssd1 vssd1 vccd1 vccd1 fanout644/X sky130_fd_sc_hd__clkbuf_8
X_20036_ _20036_/A _20036_/B vssd1 vssd1 vccd1 vccd1 _20039_/A sky130_fd_sc_hd__xnor2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14634__B1 _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout59_A _10791_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17179__A2 _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21987_ _22020_/CLK _21987_/D vssd1 vssd1 vccd1 vccd1 hold139/A sky130_fd_sc_hd__dfxtp_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _12261_/A _13155_/B _13157_/A _12269_/B vssd1 vssd1 vccd1 vccd1 _11741_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20938_ _20938_/A _20938_/B vssd1 vssd1 vccd1 vccd1 _20949_/A sky130_fd_sc_hd__or2_1
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ _11672_/A _11672_/B vssd1 vssd1 vccd1 vccd1 _11671_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20869_ _20869_/A _20869_/B vssd1 vssd1 vccd1 vccd1 _20872_/C sky130_fd_sc_hd__nand2_1
XANTENNA__16218__A _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13410_ _13410_/A _13410_/B vssd1 vssd1 vccd1 vccd1 _13413_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_14_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14390_ _15375_/A _14391_/B _14391_/C _14391_/D vssd1 vssd1 vccd1 vccd1 _14393_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13341_ _13337_/X _13339_/Y _13199_/B _13199_/Y vssd1 vssd1 vccd1 vccd1 _13343_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19529__A _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16060_ _16171_/A vssd1 vssd1 vccd1 vccd1 _16060_/Y sky130_fd_sc_hd__inv_2
X_13272_ _13858_/A _13573_/D _13416_/A _13270_/Y vssd1 vssd1 vccd1 vccd1 _13273_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_32_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15011_ _15012_/A _15012_/B _15012_/C _15012_/D vssd1 vssd1 vccd1 vccd1 _15011_/Y
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_20_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12223_ _12223_/A _12269_/D vssd1 vssd1 vccd1 vccd1 _12224_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13912__A2 _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17103__A2 _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17991__B _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12154_ _12154_/A _12154_/B vssd1 vssd1 vccd1 vccd1 _12157_/A sky130_fd_sc_hd__xnor2_1
X_11105_ _10881_/X hold106/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21699_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19264__A _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19750_ _20394_/B _19874_/B _19872_/C _19972_/A vssd1 vssd1 vccd1 vccd1 _19753_/C
+ sky130_fd_sc_hd__a22o_1
X_16962_ _16961_/B _16961_/Y _16916_/Y vssd1 vssd1 vccd1 vccd1 _16962_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_21_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12085_ _12066_/A _12066_/C _12066_/B vssd1 vssd1 vccd1 vccd1 _12085_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18701_ _18701_/A _18853_/B _18702_/B vssd1 vssd1 vccd1 vccd1 _18866_/A sky130_fd_sc_hd__or3b_1
X_15913_ _16399_/A _15913_/B _15913_/C _16102_/A vssd1 vssd1 vccd1 vccd1 _16102_/B
+ sky130_fd_sc_hd__nand4_1
X_11036_ mstream_o[110] hold306/X _11039_/S vssd1 vssd1 vccd1 vccd1 hold307/A sky130_fd_sc_hd__mux2_1
X_16893_ _16888_/A _16887_/Y _16880_/X vssd1 vssd1 vccd1 vccd1 _16896_/A sky130_fd_sc_hd__a21oi_1
X_19681_ _19681_/A _19681_/B vssd1 vssd1 vccd1 vccd1 _19683_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__19414__D _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13516__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15844_ _15844_/A _15844_/B vssd1 vssd1 vccd1 vccd1 _15846_/B sky130_fd_sc_hd__xnor2_1
X_18632_ _18632_/A _18632_/B _18632_/C vssd1 vssd1 vccd1 vccd1 _18632_/Y sky130_fd_sc_hd__nor3_2
XANTENNA__20410__A2 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15775_ _16031_/A _15775_/B vssd1 vssd1 vccd1 vccd1 _15776_/B sky130_fd_sc_hd__or2_1
X_18563_ _18563_/A vssd1 vssd1 vccd1 vccd1 _18563_/Y sky130_fd_sc_hd__inv_2
XTAP_3560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12987_ _12988_/A _12988_/B vssd1 vssd1 vccd1 vccd1 _13104_/B sky130_fd_sc_hd__nand2b_1
XTAP_3571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14726_ _15076_/B _15368_/D _15234_/C _14557_/A vssd1 vssd1 vccd1 vccd1 _14729_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17514_ _17514_/A vssd1 vssd1 vccd1 vccd1 _17514_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_115_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18494_ _19438_/B _19414_/C _19866_/D _19438_/A vssd1 vssd1 vccd1 vccd1 _18495_/B
+ sky130_fd_sc_hd__a22o_1
X_11938_ _11938_/A _11938_/B vssd1 vssd1 vccd1 vccd1 _11940_/B sky130_fd_sc_hd__xnor2_1
XTAP_2870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19430__C _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17445_ _17445_/A _17445_/B vssd1 vssd1 vccd1 vccd1 _17446_/B sky130_fd_sc_hd__nor2_1
X_14657_ _15961_/D _15838_/D _15112_/D vssd1 vssd1 vccd1 vccd1 _14657_/X sky130_fd_sc_hd__and3_1
X_11869_ _11869_/A _11869_/B vssd1 vssd1 vccd1 vccd1 _11870_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_131_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15032__A _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13608_ _13608_/A _13608_/B vssd1 vssd1 vccd1 vccd1 _13618_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17376_ hold193/A fanout7/X _17375_/X vssd1 vssd1 vccd1 vccd1 _17376_/X sky130_fd_sc_hd__a21bo_1
X_14588_ _14588_/A _14588_/B vssd1 vssd1 vccd1 vccd1 _14591_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_144_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16327_ _16327_/A _16327_/B vssd1 vssd1 vccd1 vccd1 _16329_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_43_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19115_ _19115_/A _19115_/B vssd1 vssd1 vccd1 vccd1 _19135_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_55_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13539_ _13539_/A _13539_/B _13539_/C vssd1 vssd1 vccd1 vccd1 _13539_/X sky130_fd_sc_hd__and3_1
XFILLER_0_70_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12094__C _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19046_ _19046_/A _19046_/B vssd1 vssd1 vccd1 vccd1 _19048_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14156__A2 _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16258_ _16363_/A hold189/A _10978_/Y fanout5/X _16257_/Y vssd1 vssd1 vccd1 vccd1
+ _16258_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_2_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15209_ _15492_/A _15209_/B vssd1 vssd1 vccd1 vccd1 _15210_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16189_ _16303_/A _16187_/X _16070_/B _16071_/Y vssd1 vssd1 vccd1 vccd1 _16191_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11719__B _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19948_ _19816_/A _19816_/B _19817_/Y vssd1 vssd1 vccd1 vccd1 _20075_/A sky130_fd_sc_hd__a21o_1
XANTENNA__11678__B1 _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19879_ _19879_/A _19879_/B _19879_/C vssd1 vssd1 vccd1 vccd1 _19879_/X sky130_fd_sc_hd__and3_2
XANTENNA__15852__D _16418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21910_ _21945_/CLK _21910_/D vssd1 vssd1 vccd1 vccd1 hold273/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21841_ _21845_/CLK _21841_/D vssd1 vssd1 vccd1 vccd1 _21841_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA_fanout263_A _21802_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12269__C _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_35_clk_i_A clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21772_ _21789_/CLK _21772_/D vssd1 vssd1 vccd1 vccd1 _21772_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__21362__B1 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20723_ _20855_/A _20723_/B vssd1 vssd1 vccd1 vccd1 _20724_/B sky130_fd_sc_hd__nor2_1
XANTENNA__14919__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout430_A _12242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout528_A _14659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20654_ _20654_/A _20654_/B vssd1 vssd1 vccd1 vccd1 _20656_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_110_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20585_ _20721_/D _21291_/B _20586_/C _20586_/D vssd1 vssd1 vccd1 vccd1 _20587_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_2_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17333__A2 _17666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21206_ _21206_/A _21206_/B vssd1 vssd1 vccd1 vccd1 _21226_/A sky130_fd_sc_hd__xor2_2
XANTENNA__18294__B1 _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__B _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17019__D _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21137_ _21137_/A _21137_/B vssd1 vssd1 vccd1 vccd1 _21137_/Y sky130_fd_sc_hd__xnor2_1
Xfanout430 _12242_/B vssd1 vssd1 vccd1 vccd1 _12094_/B sky130_fd_sc_hd__buf_4
XFILLER_0_100_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout441 _14572_/A vssd1 vssd1 vccd1 vccd1 _12784_/A sky130_fd_sc_hd__buf_2
Xfanout452 _21758_/Q vssd1 vssd1 vccd1 vccd1 _14248_/A sky130_fd_sc_hd__clkbuf_8
Xfanout463 _21753_/Q vssd1 vssd1 vccd1 vccd1 _15098_/B sky130_fd_sc_hd__clkbuf_8
X_21068_ _21069_/A _21069_/B vssd1 vssd1 vccd1 vccd1 _21068_/X sky130_fd_sc_hd__and2_1
Xfanout474 _15093_/B vssd1 vssd1 vccd1 vccd1 _14077_/B sky130_fd_sc_hd__buf_4
XANTENNA__18597__A1 _19531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout485 _21748_/Q vssd1 vssd1 vccd1 vccd1 _16424_/A sky130_fd_sc_hd__clkbuf_4
Xfanout496 _16404_/A vssd1 vssd1 vccd1 vccd1 _16196_/B sky130_fd_sc_hd__buf_4
XANTENNA__19794__B1 _14918_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12910_ _14572_/A _14384_/D vssd1 vssd1 vccd1 vccd1 _12913_/A sky130_fd_sc_hd__and2_1
XANTENNA__11645__A _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20019_ _20168_/A _20017_/X _19915_/Y _19917_/X vssd1 vssd1 vccd1 vccd1 _20020_/D
+ sky130_fd_sc_hd__a211o_1
X_13890_ _13886_/Y _13887_/X _13730_/Y _13733_/X vssd1 vssd1 vccd1 vccd1 _13948_/B
+ sky130_fd_sc_hd__a211oi_2
X_12841_ _12842_/B vssd1 vssd1 vccd1 vccd1 _12841_/Y sky130_fd_sc_hd__inv_2
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19531__B _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14083__A1 _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14083__B2 _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20677__B _21040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13860__A _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15560_ _15560_/A _15560_/B _15560_/C vssd1 vssd1 vccd1 vccd1 _15561_/C sky130_fd_sc_hd__nand3_2
XANTENNA__17332__A _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ _13155_/A _12771_/C _21765_/Q _14195_/A vssd1 vssd1 vccd1 vccd1 _12773_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21353__B1 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14511_ _14509_/X _14511_/B vssd1 vssd1 vccd1 vccd1 _14512_/B sky130_fd_sc_hd__nand2b_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _11723_/A _11723_/B vssd1 vssd1 vccd1 vccd1 _11736_/A sky130_fd_sc_hd__xnor2_2
X_15491_ _15625_/A _15491_/B vssd1 vssd1 vccd1 vccd1 _15496_/A sky130_fd_sc_hd__or2_1
XFILLER_0_90_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17230_ _17231_/A _17231_/B vssd1 vssd1 vccd1 vccd1 _17317_/B sky130_fd_sc_hd__nand2_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14442_ _14442_/A _14442_/B vssd1 vssd1 vccd1 vccd1 _14443_/B sky130_fd_sc_hd__xor2_2
XANTENNA__12907__C _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11654_ _11652_/B _11652_/C _11652_/A vssd1 vssd1 vccd1 vccd1 _11655_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout70 _19179_/C vssd1 vssd1 vccd1 vccd1 _20838_/D sky130_fd_sc_hd__buf_4
XFILLER_0_65_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout81 _19030_/C vssd1 vssd1 vccd1 vccd1 _19199_/C sky130_fd_sc_hd__buf_4
X_17161_ _17005_/Y _17008_/X _17049_/B _17117_/A vssd1 vssd1 vccd1 vccd1 _17161_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_36_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout92 _21844_/Q vssd1 vssd1 vccd1 vccd1 _20265_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14373_ _14373_/A _14373_/B _14373_/C vssd1 vssd1 vccd1 vccd1 _14375_/B sky130_fd_sc_hd__nand3_1
XANTENNA__19259__A _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11585_ _11585_/A _11585_/B vssd1 vssd1 vccd1 vccd1 _11593_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_80_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16112_ _16112_/A _16112_/B vssd1 vssd1 vccd1 vccd1 _16114_/C sky130_fd_sc_hd__xnor2_1
X_13324_ _14572_/A _14077_/B vssd1 vssd1 vccd1 vccd1 _13327_/A sky130_fd_sc_hd__and2_1
XANTENNA__21301__B _21816_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17092_ _17144_/A _17145_/B _17146_/C _17129_/B vssd1 vssd1 vccd1 vccd1 _17094_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_49_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16043_ _16043_/A _16213_/B vssd1 vssd1 vccd1 vccd1 _16054_/A sky130_fd_sc_hd__nand2_1
X_13255_ _13858_/C _13254_/X _13253_/X vssd1 vssd1 vccd1 vccd1 _13257_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__18313__D _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13897__A1 _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13897__B2 _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17088__A1 _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12206_ _12207_/A _12207_/B _12207_/C vssd1 vssd1 vccd1 vccd1 _12206_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__17088__B2 _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13186_ _14089_/A _14087_/A _14077_/B _14234_/C vssd1 vssd1 vccd1 vccd1 _13188_/B
+ sky130_fd_sc_hd__nand4_1
X_19802_ _20026_/B _20178_/D _20838_/C _20838_/D vssd1 vssd1 vccd1 vccd1 _19804_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_23_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12137_ _12268_/A _12214_/C vssd1 vssd1 vccd1 vccd1 _12139_/B sky130_fd_sc_hd__and2_1
X_17994_ _19008_/D _19223_/B vssd1 vssd1 vccd1 vccd1 _17995_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19733_ _20088_/A _20242_/D _19734_/C _19849_/A vssd1 vssd1 vccd1 vccd1 _19735_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16768__D _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16945_ _16946_/A _16946_/B _16946_/C vssd1 vssd1 vccd1 vccd1 _16945_/Y sky130_fd_sc_hd__nor3_2
X_12068_ _12066_/A _12065_/Y _12067_/X _12011_/Y vssd1 vssd1 vccd1 vccd1 _12076_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__12321__A1 _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12321__B2 _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ mstream_o[93] hold41/X _11027_/S vssd1 vssd1 vccd1 vccd1 _21630_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13473__C _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19664_ _20590_/D _19664_/B _20733_/C _20606_/D vssd1 vssd1 vccd1 vccd1 _19820_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__20395__A1 _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16876_ _16876_/A _16876_/B _16876_/C vssd1 vssd1 vccd1 vccd1 _16890_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_95_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18615_ _19535_/A _18929_/B _19087_/B _19695_/A vssd1 vssd1 vccd1 vccd1 _18618_/A
+ sky130_fd_sc_hd__a22o_1
X_15827_ _15823_/X _15824_/Y _15650_/B _15689_/Y vssd1 vssd1 vccd1 vccd1 _15874_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_126_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14074__A1 _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19595_ _19591_/X _19593_/Y _19444_/A _19847_/A vssd1 vssd1 vccd1 vccd1 _19595_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14074__B2 _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18338__A _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15758_ _16016_/A _15758_/B vssd1 vssd1 vccd1 vccd1 _21404_/B sky130_fd_sc_hd__xnor2_2
X_18546_ _19013_/C _18545_/X _18544_/X vssd1 vssd1 vccd1 vccd1 _18548_/A sky130_fd_sc_hd__a21bo_1
XTAP_3390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21344__B1 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14709_ _14709_/A _14709_/B vssd1 vssd1 vccd1 vccd1 _14711_/B sky130_fd_sc_hd__or2_2
X_15689_ _15689_/A _15689_/B _15689_/C vssd1 vssd1 vccd1 vccd1 _15689_/Y sky130_fd_sc_hd__nor3_4
X_18477_ _18478_/A _18478_/B _18478_/C vssd1 vssd1 vccd1 vccd1 _18477_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15574__A1 _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17428_ _17312_/X _17314_/X _17426_/X _17427_/Y vssd1 vssd1 vccd1 vccd1 _17466_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11721__C _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17359_ _17356_/X _17357_/Y _17256_/C _17255_/Y vssd1 vssd1 vccd1 vccd1 _17360_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_126_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21211__B _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20370_ _20370_/A _20370_/B vssd1 vssd1 vccd1 vccd1 _20371_/B sky130_fd_sc_hd__and2_1
XFILLER_0_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19029_ _20032_/D _19199_/C _19199_/D _19810_/D vssd1 vssd1 vccd1 vccd1 _19032_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout109_A _19692_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22040_ _22049_/CLK _22040_/D vssd1 vssd1 vccd1 vccd1 hold272/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12736__A1_N _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17417__A _17417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16040__B _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout478_A _14217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16975__B _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19351__B _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout645_A _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19528__B1 _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13680__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21824_ _21829_/CLK _21824_/D vssd1 vssd1 vccd1 vccd1 _21824_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_78_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21335__B1 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11912__B _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21755_ _22063_/CLK _21755_/D vssd1 vssd1 vccd1 vccd1 _21755_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_109_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11404__S _11446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20706_ _20707_/A _20707_/B _20707_/C vssd1 vssd1 vccd1 vccd1 _20836_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21686_ _22069_/CLK _21686_/D vssd1 vssd1 vccd1 vccd1 hold85/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20637_ _20634_/Y _20635_/X _20468_/B _20471_/A vssd1 vssd1 vccd1 vccd1 _20638_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13839__B _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11370_ hold186/X fanout29/X _11369_/X vssd1 vssd1 vccd1 vccd1 _11370_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20568_ _20569_/A _20569_/B vssd1 vssd1 vccd1 vccd1 _20698_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16215__B _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18711__A _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20499_ _20499_/A _20499_/B _20499_/C _20499_/D vssd1 vssd1 vccd1 vccd1 _20499_/Y
+ sky130_fd_sc_hd__nor4_4
XFILLER_0_104_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13040_ _13040_/A _13040_/B _13040_/C vssd1 vssd1 vccd1 vccd1 _13042_/A sky130_fd_sc_hd__and3_1
XFILLER_0_30_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16817__A1 _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14991_ _14862_/A _14862_/C _14862_/B vssd1 vssd1 vccd1 vccd1 _15006_/A sky130_fd_sc_hd__a21bo_1
Xfanout260 _19823_/A vssd1 vssd1 vccd1 vccd1 _19230_/A sky130_fd_sc_hd__clkbuf_4
Xfanout271 _17417_/A vssd1 vssd1 vccd1 vccd1 _19664_/B sky130_fd_sc_hd__buf_4
XANTENNA__12303__A1 _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14389__C _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout282 _21799_/Q vssd1 vssd1 vccd1 vccd1 _18008_/B sky130_fd_sc_hd__buf_4
X_13942_ _13938_/X _13940_/Y _13790_/B _13790_/Y vssd1 vssd1 vccd1 vccd1 _13942_/Y
+ sky130_fd_sc_hd__o211ai_1
X_16730_ _16730_/A _16730_/B _16730_/C vssd1 vssd1 vccd1 vccd1 _16738_/A sky130_fd_sc_hd__nand3_1
Xfanout293 _16743_/C vssd1 vssd1 vccd1 vccd1 _17013_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16661_ _17141_/A _17434_/B _17433_/A _17141_/B vssd1 vssd1 vccd1 vccd1 _16662_/C
+ sky130_fd_sc_hd__a22o_1
X_13873_ _14195_/A _14537_/A _13744_/A _13743_/A vssd1 vssd1 vccd1 vccd1 _13878_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14056__A1 _14212_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15612_ _15612_/A _15612_/B _15612_/C _15612_/D vssd1 vssd1 vccd1 vccd1 _15612_/Y
+ sky130_fd_sc_hd__nor4_4
X_18400_ _21791_/Q _18703_/A _19013_/C _19179_/C vssd1 vssd1 vccd1 vccd1 _18420_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__17793__A2 _18789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12824_ _12824_/A _12824_/B vssd1 vssd1 vccd1 vccd1 _12827_/A sky130_fd_sc_hd__nor2_2
XANTENNA__20838__D _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16592_ _17526_/B _16813_/A _16743_/B _17525_/A vssd1 vssd1 vccd1 vccd1 _16592_/X
+ sky130_fd_sc_hd__and4_1
X_19380_ _19382_/A _19382_/B _19382_/C _19382_/D vssd1 vssd1 vccd1 vccd1 _19380_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20129__A1 _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15543_ _15543_/A _15543_/B vssd1 vssd1 vccd1 vccd1 _15545_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_97_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18331_ _18327_/X _18328_/Y _18176_/X _18178_/X vssd1 vssd1 vccd1 vccd1 _18368_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_57_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17997__A _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12755_ _12877_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _12759_/A sky130_fd_sc_hd__nand2_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18262_ _18263_/A _18263_/B vssd1 vssd1 vccd1 vccd1 _18262_/Y sky130_fd_sc_hd__nand2_1
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ _12267_/A _12094_/B _13017_/A _12444_/B vssd1 vssd1 vccd1 vccd1 _11709_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__12637__C _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15474_ _15473_/B _15473_/C _15473_/A vssd1 vssd1 vccd1 vccd1 _15475_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_126_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ _12687_/A _12687_/B _12687_/C vssd1 vssd1 vccd1 vccd1 _12686_/X sky130_fd_sc_hd__and3_1
XFILLER_0_84_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14425_ _14426_/A _14426_/B vssd1 vssd1 vccd1 vccd1 _14425_/X sky130_fd_sc_hd__and2b_1
X_17213_ _17213_/A _17213_/B vssd1 vssd1 vccd1 vccd1 _17215_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18193_ _18193_/A _18193_/B vssd1 vssd1 vccd1 vccd1 _18195_/B sky130_fd_sc_hd__xnor2_2
X_11637_ _12426_/B _12512_/A vssd1 vssd1 vccd1 vccd1 _11640_/A sky130_fd_sc_hd__and2_1
XFILLER_0_155_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17144_ _17144_/A _17146_/D vssd1 vssd1 vccd1 vccd1 _17150_/A sky130_fd_sc_hd__nand2_1
X_14356_ _14813_/A _15022_/B _14357_/C _14357_/D vssd1 vssd1 vccd1 vccd1 _14356_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_107_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11568_ _12229_/A _12155_/B _12528_/B _12619_/A vssd1 vssd1 vccd1 vccd1 _11568_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_141_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13307_ _13306_/B _13306_/C _13306_/A vssd1 vssd1 vccd1 vccd1 _13343_/B sky130_fd_sc_hd__a21oi_2
X_17075_ _17081_/A _17075_/B vssd1 vssd1 vccd1 vccd1 _17078_/B sky130_fd_sc_hd__nand2_1
X_14287_ _14289_/A _14289_/B vssd1 vssd1 vccd1 vccd1 _14288_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13468__C _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11499_ _11502_/A1 t2x[16] v1z[16] fanout20/X _11498_/X vssd1 vssd1 vccd1 vccd1 _11499_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16026_ hold36/X _16025_/X fanout1/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__mux2_1
XFILLER_0_0_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13238_ _13376_/B _13237_/C _13237_/A vssd1 vssd1 vccd1 vccd1 _13239_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17237__A _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20604__A2 _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13169_ _13169_/A _13169_/B vssd1 vssd1 vccd1 vccd1 _13179_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13098__A2 _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17977_ _21791_/Q _18703_/A _19030_/C _19199_/D vssd1 vssd1 vccd1 vccd1 _18117_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19716_ _19715_/B _19715_/C _19715_/A vssd1 vssd1 vccd1 vccd1 _19716_/X sky130_fd_sc_hd__a21o_1
X_16928_ _16928_/A _16928_/B vssd1 vssd1 vccd1 vccd1 _16930_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_137_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16795__B _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17233__A1 _17334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17233__B2 _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19647_ _19647_/A _19647_/B vssd1 vssd1 vccd1 vccd1 _19649_/A sky130_fd_sc_hd__xnor2_2
X_16859_ _16859_/A _16859_/B vssd1 vssd1 vccd1 vccd1 _17167_/A sky130_fd_sc_hd__and2_1
XFILLER_0_149_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19578_ _19578_/A _19578_/B _19578_/C vssd1 vssd1 vccd1 vccd1 _19581_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_133_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12828__B _17599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18529_ _18529_/A _18529_/B _18529_/C vssd1 vssd1 vccd1 vccd1 _18684_/B sky130_fd_sc_hd__or3_2
XFILLER_0_87_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13270__A2 _13269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11281__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21540_ mstream_o[3] hold21/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22067_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_34_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13558__B1 _14663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21471_ hold154/X sstream_i[48] _21494_/S vssd1 vssd1 vccd1 vccd1 _21998_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13419__A1_N _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout226_A _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11033__A1 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20422_ _20423_/A _20423_/B vssd1 vssd1 vccd1 vccd1 _20616_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_132_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11584__A2 _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20353_ _20354_/A _20354_/B vssd1 vssd1 vccd1 vccd1 _20353_/X sky130_fd_sc_hd__or2_1
XFILLER_0_144_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16976__A1_N _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20284_ _20287_/D vssd1 vssd1 vccd1 vccd1 _20284_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_144_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17792__D _21040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout595_A _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22023_ _22038_/CLK _22023_/D vssd1 vssd1 vccd1 vccd1 hold308/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13394__B _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20004__C _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 hold68/A vssd1 vssd1 vccd1 vccd1 hold68/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 hold79/A vssd1 vssd1 vccd1 vccd1 hold79/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10870_ hold140/A hold97/A vssd1 vssd1 vccd1 vccd1 _10880_/A sky130_fd_sc_hd__and2_1
XFILLER_0_78_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21807_ _21809_/CLK _21807_/D vssd1 vssd1 vccd1 vccd1 _21807_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13261__A2 _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15538__A1 _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12540_ _12540_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _12542_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_137_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21738_ _21803_/CLK _21738_/D vssd1 vssd1 vccd1 vccd1 _21738_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__16735__B1 _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20674__C _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12471_ _12471_/A _12471_/B _12471_/C vssd1 vssd1 vccd1 vccd1 _12471_/Y sky130_fd_sc_hd__nand3_2
X_21669_ _21906_/CLK _21669_/D vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14210_ _14081_/A _14080_/B _14078_/X vssd1 vssd1 vccd1 vccd1 _14226_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_124_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15130__A _16173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11024__A1 hold239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11422_ _11421_/X _21311_/A _11446_/S vssd1 vssd1 vccd1 vccd1 _21812_/D sky130_fd_sc_hd__mux2_1
X_15190_ _15346_/A _15188_/X _14962_/Y _14965_/X vssd1 vssd1 vccd1 vccd1 _15191_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12772__A1 _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14141_ _14141_/A _14141_/B vssd1 vssd1 vccd1 vccd1 _14144_/A sky130_fd_sc_hd__xnor2_1
X_11353_ _21718_/D _21724_/D _11126_/B _21422_/A vssd1 vssd1 vccd1 vccd1 wire16/A
+ sky130_fd_sc_hd__o31ai_2
XANTENNA__19537__A _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12772__B2 _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_4_clk_i_A _21806_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14072_ _14072_/A _14072_/B vssd1 vssd1 vccd1 vccd1 _14105_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11089__B _11089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11284_ _13012_/B _11283_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21772_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_67_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13721__B1 _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13023_ _13023_/A _13023_/B _13023_/C vssd1 vssd1 vccd1 vccd1 _13148_/A sky130_fd_sc_hd__nand3_2
X_17900_ _20583_/A _18319_/B _18622_/B _19892_/A vssd1 vssd1 vccd1 vccd1 _17901_/C
+ sky130_fd_sc_hd__a22o_1
X_18880_ _18716_/A _18717_/Y _18878_/X _18879_/Y vssd1 vssd1 vccd1 vccd1 _18881_/A
+ sky130_fd_sc_hd__a211oi_2
X_17831_ _17831_/A _17831_/B vssd1 vssd1 vccd1 vccd1 _17832_/B sky130_fd_sc_hd__nand2_2
X_17762_ _18030_/B _18624_/A vssd1 vssd1 vccd1 vccd1 _17765_/A sky130_fd_sc_hd__and2_1
X_14974_ _14974_/A _14974_/B vssd1 vssd1 vccd1 vccd1 _14974_/X sky130_fd_sc_hd__or2_1
XFILLER_0_89_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19703__C _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19501_ _19501_/A _19501_/B vssd1 vssd1 vccd1 vccd1 _19502_/B sky130_fd_sc_hd__and2_1
XFILLER_0_117_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16713_ _16682_/A _16682_/B _16682_/C vssd1 vssd1 vccd1 vccd1 _16713_/Y sky130_fd_sc_hd__o21ai_2
X_13925_ _14572_/A _14557_/D vssd1 vssd1 vccd1 vccd1 _13928_/A sky130_fd_sc_hd__and2_1
XFILLER_0_57_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17693_ _17718_/B _17694_/B _17693_/C _17693_/D vssd1 vssd1 vccd1 vccd1 _17693_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_88_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19432_ _19432_/A _19751_/C _19432_/C _19598_/A vssd1 vssd1 vccd1 vccd1 _19598_/B
+ sky130_fd_sc_hd__nand4_2
X_13856_ _13972_/A _13854_/X _13695_/Y _13698_/X vssd1 vssd1 vccd1 vccd1 _13952_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18319__C _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16644_ _16644_/A _16644_/B vssd1 vssd1 vccd1 vccd1 _16645_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__16974__B1 _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12807_ _12837_/B _12808_/B _12807_/C _12807_/D vssd1 vssd1 vccd1 vccd1 _12807_/X
+ sky130_fd_sc_hd__and4bb_2
XFILLER_0_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19363_ _19363_/A _19363_/B vssd1 vssd1 vccd1 vccd1 _19365_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_57_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13787_ _13787_/A _13787_/B _13787_/C vssd1 vssd1 vccd1 vccd1 _13790_/B sky130_fd_sc_hd__nand3_2
X_16575_ _17206_/B _17619_/B _17211_/A _16575_/D vssd1 vssd1 vccd1 vccd1 _17211_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__14134__A1_N _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10999_ mstream_o[73] hold25/X _11005_/S vssd1 vssd1 vccd1 vccd1 _21610_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_128_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18616__A _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11044__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17520__A _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18314_ _19529_/B _18769_/B _18314_/C _18314_/D vssd1 vssd1 vccd1 vccd1 _18316_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15526_ _15526_/A _15648_/B vssd1 vssd1 vccd1 vccd1 _15529_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12738_ _12856_/B _12736_/X _12639_/C _12641_/A vssd1 vssd1 vccd1 vccd1 _12739_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_127_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16726__B1 _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19294_ _19295_/A _19295_/B vssd1 vssd1 vccd1 vccd1 _19294_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_72_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20522__A1 _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18335__B _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15457_ _15457_/A _15587_/B vssd1 vssd1 vccd1 vccd1 _15459_/B sky130_fd_sc_hd__or2_1
X_18245_ _18394_/A _18245_/B vssd1 vssd1 vccd1 vccd1 _21358_/B sky130_fd_sc_hd__xnor2_4
X_12669_ _13173_/C _12780_/A _12780_/B _13034_/D vssd1 vssd1 vccd1 vccd1 _12669_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_127_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14408_ _14859_/A _15091_/C _14408_/C _14554_/A vssd1 vssd1 vccd1 vccd1 _14554_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_115_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15388_ _15224_/Y _15248_/Y _15385_/Y _15386_/X vssd1 vssd1 vccd1 vccd1 _15426_/B
+ sky130_fd_sc_hd__a211oi_4
X_18176_ _18177_/B _18177_/A vssd1 vssd1 vccd1 vccd1 _18176_/X sky130_fd_sc_hd__and2b_2
XFILLER_0_128_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14339_ _14340_/A _14340_/B vssd1 vssd1 vccd1 vccd1 _14339_/Y sky130_fd_sc_hd__nor2_1
X_17127_ _17123_/X _17140_/A _17089_/X _17122_/Y vssd1 vssd1 vccd1 vccd1 _17133_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_111_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17058_ _17058_/A _17058_/B vssd1 vssd1 vccd1 vccd1 _17074_/B sky130_fd_sc_hd__and2_1
X_16009_ _16010_/A _16010_/B vssd1 vssd1 vccd1 vccd1 _16009_/X sky130_fd_sc_hd__or2_1
XFILLER_0_111_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18651__B1 _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11219__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18403__B1 _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20971_ _20971_/A _20971_/B vssd1 vssd1 vccd1 vccd1 _20973_/B sky130_fd_sc_hd__or2_1
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout176_A _16734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11254__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11254__B2 _11459_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21523_ hold290/X sstream_i[100] _21536_/S vssd1 vssd1 vccd1 vccd1 _22050_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_29_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout510_A _21742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout608_A _21718_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21454_ hold148/X sstream_i[31] _21507_/S vssd1 vssd1 vccd1 vccd1 _21981_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_90_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20405_ _20239_/A _20238_/Y _20260_/X vssd1 vssd1 vccd1 vccd1 _20407_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_16_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21385_ _21720_/D _19636_/B fanout40/X vssd1 vssd1 vccd1 vccd1 _21385_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__17142__B1 _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18296__A2_N _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20336_ _20336_/A _20472_/B vssd1 vssd1 vccd1 vccd1 _20338_/B sky130_fd_sc_hd__or2_1
XFILLER_0_12_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19507__D _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold290_A hold290/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20267_ _21199_/A _21264_/A _20267_/C _20473_/A vssd1 vssd1 vccd1 vccd1 _20473_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_101_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22006_ _22013_/CLK _22006_/D vssd1 vssd1 vccd1 vccd1 hold130/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout89_A _18894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11637__B _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20198_ _20198_/A _20198_/B vssd1 vssd1 vccd1 vccd1 _20200_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__19804__B _20841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11129__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19092__A _19092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21529__A0 hold299/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19198__A1 _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20669__C _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17324__B _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11971_ _11971_/A _11971_/B _11971_/C vssd1 vssd1 vccd1 vccd1 _11982_/A sky130_fd_sc_hd__nand3_2
X_13710_ _13864_/B _13867_/A _14354_/C _14663_/D vssd1 vssd1 vccd1 vccd1 _13710_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_98_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10922_ hold20/A hold50/A vssd1 vssd1 vccd1 vccd1 _10923_/B sky130_fd_sc_hd__nand2_1
X_14690_ _14690_/A _14690_/B vssd1 vssd1 vccd1 vccd1 _14711_/A sky130_fd_sc_hd__nand2_2
XANTENNA__13571__C _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20388__D _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11493__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20966__A _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13641_ _13637_/X _13639_/Y _13486_/B _13486_/Y vssd1 vssd1 vccd1 vccd1 _13643_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10853_ mstream_o[43] _10852_/X _21579_/S vssd1 vssd1 vccd1 vccd1 _21580_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_116_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13234__A2 _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16360_ _16360_/A _16360_/B vssd1 vssd1 vccd1 vccd1 _16362_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11245__A1 _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16882__C _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13572_ _13864_/B _16286_/A _13570_/Y _13720_/A vssd1 vssd1 vccd1 vccd1 _13572_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_94_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11245__B2 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15311_ _15311_/A _15311_/B vssd1 vssd1 vccd1 vccd1 _15314_/A sky130_fd_sc_hd__xnor2_1
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12523_ _12522_/B _12522_/C _12522_/A vssd1 vssd1 vccd1 vccd1 _12523_/X sky130_fd_sc_hd__o21a_1
X_16291_ _16291_/A _16291_/B vssd1 vssd1 vccd1 vccd1 _16293_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15242_ _15242_/A _15242_/B vssd1 vssd1 vccd1 vccd1 _15244_/B sky130_fd_sc_hd__xor2_2
X_18030_ _19823_/A _18030_/B _18767_/B _18616_/D vssd1 vssd1 vccd1 vccd1 _18031_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_23_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12454_ _13155_/A _13155_/B _12780_/A _12780_/B vssd1 vssd1 vccd1 vccd1 _12455_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_81_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17994__B _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11405_ _11447_/A1 hold279/A fanout49/X hold184/A vssd1 vssd1 vccd1 vccd1 _11405_/X
+ sky130_fd_sc_hd__a22o_1
X_15173_ _15702_/D _15174_/D _15171_/Y _15316_/A vssd1 vssd1 vccd1 vccd1 _15175_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_105_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12385_ _11840_/A _11839_/Y _12383_/Y _12384_/X vssd1 vssd1 vccd1 vccd1 _12708_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__18171__A _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14124_ _14285_/B _14123_/C _14290_/A vssd1 vssd1 vccd1 vccd1 _14291_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11336_ _15829_/C _11335_/X _11348_/S vssd1 vssd1 vccd1 vccd1 _21785_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_50_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19981_ _19877_/B _19879_/B _20126_/A _19980_/Y vssd1 vssd1 vccd1 vccd1 _20126_/B
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__14498__A1 _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14498__B2 _14659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14055_ _15763_/A _14384_/A _14212_/D vssd1 vssd1 vccd1 vccd1 _14055_/X sky130_fd_sc_hd__and3_1
X_18932_ _19092_/B _19906_/C vssd1 vssd1 vccd1 vccd1 _18936_/A sky130_fd_sc_hd__and2_1
X_11267_ fanout58/X v0z[10] fanout17/X _11266_/X vssd1 vssd1 vccd1 vccd1 _11267_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13006_ _13003_/A _13004_/Y _12891_/Y _12895_/A vssd1 vssd1 vccd1 vccd1 _13006_/Y
+ sky130_fd_sc_hd__o211ai_1
X_18863_ _18863_/A _18863_/B vssd1 vssd1 vccd1 vccd1 _18864_/B sky130_fd_sc_hd__or2_1
XANTENNA__11547__B _11555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11198_ _13913_/C _11197_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21749_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11720__A2 _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17814_ _17810_/X _17811_/Y _17689_/C _17688_/Y vssd1 vssd1 vccd1 vccd1 _17815_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_59_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15961__C hold319/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18794_ _19587_/B _19751_/C _20242_/C _19587_/A vssd1 vssd1 vccd1 vccd1 _18794_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_59_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21037__A _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17745_ _17743_/X _17745_/B vssd1 vssd1 vccd1 vccd1 _17746_/B sky130_fd_sc_hd__and2b_1
XANTENNA__17234__B _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14957_ _14956_/B _14956_/C _14956_/A vssd1 vssd1 vccd1 vccd1 _14957_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__12659__A _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13908_ _13753_/Y _13755_/X _13906_/X _13907_/Y vssd1 vssd1 vccd1 vccd1 _13943_/A
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__11484__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17676_ _17676_/A _17676_/B _17676_/C vssd1 vssd1 vccd1 vccd1 _17678_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_134_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14888_ _14887_/A _14887_/B _14887_/C _14887_/D vssd1 vssd1 vccd1 vccd1 _14889_/B
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19415_ _19417_/D vssd1 vssd1 vccd1 vccd1 _19415_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_58_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16627_ _16870_/A _17526_/B _16590_/A _16588_/Y vssd1 vssd1 vccd1 vccd1 _16628_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_13839_ _13975_/B _16328_/B _13839_/C _13839_/D vssd1 vssd1 vccd1 vccd1 _13839_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_43_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20976__A2_N _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19346_ _19346_/A _19346_/B vssd1 vssd1 vccd1 vccd1 _19366_/A sky130_fd_sc_hd__or2_1
X_16558_ _16870_/A _17223_/A _16557_/B _16554_/X vssd1 vssd1 vccd1 vccd1 _16563_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_73_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15509_ _16027_/A _16391_/B _15510_/C _15670_/A vssd1 vssd1 vccd1 vccd1 _15511_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19277_ _19439_/A _20242_/C _19116_/X _19117_/X _20242_/D vssd1 vssd1 vccd1 vccd1
+ _19282_/A sky130_fd_sc_hd__a32o_1
X_16489_ _17636_/B _17387_/A _16489_/C _16489_/D vssd1 vssd1 vccd1 vccd1 _16495_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_116_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18228_ _18225_/X _18226_/Y _18087_/C _18086_/Y vssd1 vssd1 vccd1 vccd1 _18230_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18159_ _18044_/B _18046_/A _18157_/Y _18158_/X vssd1 vssd1 vccd1 vccd1 _18250_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold302 hold302/A vssd1 vssd1 vccd1 vccd1 hold302/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold313 hold313/A vssd1 vssd1 vccd1 vccd1 hold313/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 hold324/A vssd1 vssd1 vccd1 vccd1 hold324/X sky130_fd_sc_hd__dlygate4sd3_1
X_21170_ _21171_/A _21171_/B _21171_/C _21171_/D vssd1 vssd1 vccd1 vccd1 _21172_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20121_ _20121_/A _20121_/B vssd1 vssd1 vccd1 vccd1 _20124_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19416__A2 _19868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12560__C _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20052_ _20186_/A _20051_/C _20051_/A vssd1 vssd1 vccd1 vccd1 _20053_/C sky130_fd_sc_hd__a21o_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout293_A _16743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14768__B _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout460_A _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17144__B _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14661__A1 _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16667__A2_N _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout558_A _21731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14661__B2 _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_208 hold270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11475__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_219 hold277/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20954_ _20952_/B _20952_/C _20952_/A vssd1 vssd1 vccd1 vccd1 _20954_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11475__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16402__A2 _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14413__A1 _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20885_ _20885_/A _20885_/B vssd1 vssd1 vccd1 vccd1 _20885_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__14413__B2 _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18256__A _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11227__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12975__A1 _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18406__D _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20317__A_N _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21506_ hold246/X sstream_i[83] _21507_/S vssd1 vssd1 vccd1 vccd1 _22033_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_8_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12735__C _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18703__B _19185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12454__D _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21437_ hold266/X sstream_i[14] _21442_/S vssd1 vssd1 vccd1 vccd1 _21964_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19087__A _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16469__A2 _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ _12124_/X _12132_/Y _12168_/A _12167_/Y vssd1 vssd1 vccd1 vccd1 _12172_/B
+ sky130_fd_sc_hd__a211o_1
X_21368_ _21412_/A _18689_/B fanout40/X vssd1 vssd1 vccd1 vccd1 _21368_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__20026__A _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12751__B _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11121_ _10988_/Y hold67/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21715_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_43_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20319_ _20317_/D _20178_/B _21261_/B _19644_/A vssd1 vssd1 vccd1 vccd1 _20321_/C
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14024__A _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21299_ _21299_/A _21299_/B vssd1 vssd1 vccd1 vccd1 _21300_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17418__A1 _17417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11052_ _11051_/Y hold11/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21655_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17418__B2 _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18615__B1 _19087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19534__B _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13863__A _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15860_ _15860_/A _15860_/B vssd1 vssd1 vccd1 vccd1 _15862_/C sky130_fd_sc_hd__nand2_1
XANTENNA__18173__A2_N _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14811_ _16092_/D _15961_/D _15112_/D vssd1 vssd1 vccd1 vccd1 _14811_/X sky130_fd_sc_hd__and3_1
XTAP_3720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15791_ _15791_/A _15916_/B _16396_/A _16377_/B vssd1 vssd1 vccd1 vccd1 _15921_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_98_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17530_ _17520_/A _17206_/B _17419_/B _17417_/X vssd1 vssd1 vccd1 vccd1 _17532_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11466__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14742_ _14742_/A _14742_/B vssd1 vssd1 vccd1 vccd1 _14743_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_87_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11954_ _11956_/A _11956_/B vssd1 vssd1 vccd1 vccd1 _11954_/Y sky130_fd_sc_hd__nand2_1
XTAP_3764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10905_ hold102/A hold126/A vssd1 vssd1 vccd1 vccd1 _10908_/A sky130_fd_sc_hd__or2_1
XFILLER_0_86_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14673_ _14828_/B _16404_/A _16409_/A _16173_/A vssd1 vssd1 vccd1 vccd1 _14676_/C
+ sky130_fd_sc_hd__a22o_1
X_17461_ _17461_/A _17461_/B _17461_/C vssd1 vssd1 vccd1 vccd1 _17461_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__14404__A1 _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11885_ _11885_/A _11969_/A vssd1 vssd1 vccd1 vccd1 _11958_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18166__A _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14404__B2 _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19200_ _19810_/D _19201_/B _19201_/C _19348_/A vssd1 vssd1 vccd1 vccd1 _19202_/B
+ sky130_fd_sc_hd__a22o_1
X_16412_ _16412_/A _16412_/B vssd1 vssd1 vccd1 vccd1 _16413_/B sky130_fd_sc_hd__xnor2_1
X_13624_ _14572_/A _15370_/B vssd1 vssd1 vccd1 vccd1 _13627_/A sky130_fd_sc_hd__and2_1
X_10836_ _10836_/A _10836_/B vssd1 vssd1 vccd1 vccd1 _11055_/B sky130_fd_sc_hd__nor2_2
X_17392_ _17282_/A _17741_/B _17285_/B _17283_/X vssd1 vssd1 vccd1 vccd1 _17402_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_67_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19131_ _19130_/B _19130_/C _19130_/A vssd1 vssd1 vccd1 vccd1 _19133_/B sky130_fd_sc_hd__a21o_1
X_16343_ _16343_/A _16343_/B vssd1 vssd1 vccd1 vccd1 _16344_/B sky130_fd_sc_hd__xnor2_1
X_13555_ _13556_/A _13997_/C _13556_/C _13556_/D vssd1 vssd1 vccd1 vccd1 _13557_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21150__A1 _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19894__A2 _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21150__B2 _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12506_ _12605_/A _12605_/B vssd1 vssd1 vccd1 vccd1 _12606_/A sky130_fd_sc_hd__nor2_1
X_16274_ _16274_/A _16274_/B vssd1 vssd1 vccd1 vccd1 _16277_/A sky130_fd_sc_hd__xnor2_1
X_19062_ _19058_/X _19060_/Y _18897_/X _18900_/X vssd1 vssd1 vccd1 vccd1 _19063_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13486_ _13486_/A _13486_/B _13486_/C vssd1 vssd1 vccd1 vccd1 _13486_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12718__A1 _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15225_ _15225_/A _15225_/B vssd1 vssd1 vccd1 vccd1 _15249_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12718__B2 _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18013_ _18144_/B _18012_/C _18012_/A vssd1 vssd1 vccd1 vccd1 _18014_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_23_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12437_ _12437_/A _12437_/B _12437_/C vssd1 vssd1 vccd1 vccd1 _12437_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_129_1264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16414__A _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15156_ _15154_/X _15305_/B _14930_/D _14934_/B vssd1 vssd1 vccd1 vccd1 _15156_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_105_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12368_ _12367_/A _12367_/B _12367_/C vssd1 vssd1 vccd1 vccd1 _12370_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_121_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14107_ _13941_/X _13943_/X _14105_/Y _14106_/X vssd1 vssd1 vccd1 vccd1 _14107_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11319_ fanout59/X v0z[23] fanout18/X _11318_/X vssd1 vssd1 vccd1 vccd1 _11319_/X
+ sky130_fd_sc_hd__a31o_2
XANTENNA__18051__D _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11558__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15087_ _15087_/A _15223_/B _15087_/C vssd1 vssd1 vccd1 vccd1 _15108_/A sky130_fd_sc_hd__and3_1
X_19964_ _19963_/A _20095_/B _19963_/C vssd1 vssd1 vccd1 vccd1 _19984_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12299_ _13012_/B _12511_/A _11690_/B _11688_/X vssd1 vssd1 vccd1 vccd1 _12306_/A
+ sky130_fd_sc_hd__a31oi_2
X_14038_ _14038_/A _14038_/B _14190_/B vssd1 vssd1 vccd1 vccd1 _14040_/B sky130_fd_sc_hd__nand3_1
X_18915_ _18914_/B _18914_/C _18914_/A vssd1 vssd1 vccd1 vccd1 _18917_/B sky130_fd_sc_hd__a21o_1
X_19895_ _20863_/C _20416_/A _21291_/A _20416_/B vssd1 vssd1 vccd1 vccd1 _19898_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_129_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13773__A _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18846_ _18846_/A _18846_/B vssd1 vssd1 vccd1 vccd1 _18991_/A sky130_fd_sc_hd__nor2_1
XANTENNA__16093__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18777_ _18774_/Y _18775_/X _18624_/D _18625_/B vssd1 vssd1 vccd1 vccd1 _18778_/C
+ sky130_fd_sc_hd__o211ai_1
X_15989_ _15861_/Y _15863_/Y _15987_/X _15988_/Y vssd1 vssd1 vccd1 vccd1 _15991_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17728_ _17729_/B vssd1 vssd1 vccd1 vccd1 _17728_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11457__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20716__A1 _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17899__B _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17659_ _19892_/A _19432_/A _17777_/A _17659_/D vssd1 vssd1 vccd1 vccd1 _17777_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_148_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20670_ _21296_/A _21264_/A _20671_/C _20858_/A vssd1 vssd1 vccd1 vccd1 _20672_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17411__C _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19329_ _19252_/A _19252_/C _19252_/B vssd1 vssd1 vccd1 vccd1 _19368_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__16148__A1 _16036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11232__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout139_A _18929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17896__A1 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19637__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout306_A _19337_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold110 hold110/A vssd1 vssd1 vccd1 vccd1 hold110/X sky130_fd_sc_hd__dlygate4sd3_1
X_21222_ _21222_/A _21222_/B _21222_/C vssd1 vssd1 vccd1 vccd1 _21222_/Y sky130_fd_sc_hd__nand3_1
Xhold121 hold121/A vssd1 vssd1 vccd1 vccd1 hold121/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold132 hold132/A vssd1 vssd1 vccd1 vccd1 hold132/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_31_clk_i_A clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 hold143/A vssd1 vssd1 vccd1 vccd1 hold143/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11932__A2 _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold154 hold154/A vssd1 vssd1 vccd1 vccd1 hold154/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20652__B1 _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21153_ _21264_/A _21153_/B vssd1 vssd1 vccd1 vccd1 _21154_/B sky130_fd_sc_hd__nand2_1
Xhold165 hold165/A vssd1 vssd1 vccd1 vccd1 hold165/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold176 hold176/A vssd1 vssd1 vccd1 vccd1 hold176/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 hold187/A vssd1 vssd1 vccd1 vccd1 hold187/X sky130_fd_sc_hd__dlygate4sd3_1
Xfanout601 _11459_/B2 vssd1 vssd1 vccd1 vccd1 _21724_/D sky130_fd_sc_hd__clkbuf_8
XANTENNA__21376__S _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout612 _21568_/S vssd1 vssd1 vccd1 vccd1 _21554_/S sky130_fd_sc_hd__clkbuf_8
Xhold198 hold198/A vssd1 vssd1 vccd1 vccd1 hold198/X sky130_fd_sc_hd__dlygate4sd3_1
X_20104_ _20104_/A _20282_/B vssd1 vssd1 vccd1 vccd1 _20114_/A sky130_fd_sc_hd__nand2_1
X_21084_ _21084_/A _21194_/B vssd1 vssd1 vccd1 vccd1 _21086_/A sky130_fd_sc_hd__or2_2
Xfanout623 _17557_/A vssd1 vssd1 vccd1 vccd1 _19123_/A sky130_fd_sc_hd__buf_4
Xfanout634 _16380_/A vssd1 vssd1 vccd1 vccd1 _15791_/A sky130_fd_sc_hd__buf_4
Xfanout645 _21422_/A vssd1 vssd1 vccd1 vccd1 _21329_/B1 sky130_fd_sc_hd__buf_4
XFILLER_0_42_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20035_ _20035_/A _20035_/B vssd1 vssd1 vccd1 vccd1 _20036_/B sky130_fd_sc_hd__nor2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14634__B2 _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11407__S _11446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21986_ _22020_/CLK _21986_/D vssd1 vssd1 vccd1 vccd1 hold177/A sky130_fd_sc_hd__dfxtp_1
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19573__A1 _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20937_ _21110_/B _20937_/B vssd1 vssd1 vccd1 vccd1 _20952_/A sky130_fd_sc_hd__and2_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21380__A1 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11931__A _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11670_ _11670_/A _11670_/B vssd1 vssd1 vccd1 vccd1 _11672_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_55_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20868_ _20868_/A _20868_/B vssd1 vssd1 vccd1 vccd1 _20869_/B sky130_fd_sc_hd__or2_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16218__B _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20799_ _21256_/A _21153_/B _20800_/C _20800_/D vssd1 vssd1 vccd1 vccd1 _20802_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_9_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13340_ _13199_/B _13199_/Y _13337_/X _13339_/Y vssd1 vssd1 vccd1 vccd1 _13343_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_91_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19529__B _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13858__A _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13271_ _13416_/A _13270_/Y _13858_/A _13573_/D vssd1 vssd1 vccd1 vccd1 _13416_/B
+ sky130_fd_sc_hd__and4bb_1
X_15010_ _15012_/A _15012_/B _15012_/C _15012_/D vssd1 vssd1 vccd1 vccd1 _15010_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_121_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17639__A1 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12222_ _12222_/A _12222_/B vssd1 vssd1 vccd1 vccd1 _12224_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13174__A1_N _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12153_ _12153_/A _12153_/B vssd1 vssd1 vccd1 vccd1 _12154_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_130_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15114__A2 _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17991__C _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11104_ _10874_/Y hold8/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21698_/D sky130_fd_sc_hd__mux2_1
X_16961_ _16961_/A _16961_/B _16961_/C vssd1 vssd1 vccd1 vccd1 _16961_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__16862__A2 _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12084_ _12076_/A _12075_/C _12075_/B vssd1 vssd1 vccd1 vccd1 _12084_/X sky130_fd_sc_hd__a21o_1
X_18700_ _18703_/A _19181_/B _18544_/X _18545_/X _19013_/C vssd1 vssd1 vccd1 vccd1
+ _18702_/B sky130_fd_sc_hd__a32o_1
XFILLER_0_21_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15912_ _16328_/A _15788_/B _15913_/C _16102_/A vssd1 vssd1 vccd1 vccd1 _15914_/A
+ sky130_fd_sc_hd__a22o_1
X_11035_ mstream_o[109] hold262/X _11039_/S vssd1 vssd1 vccd1 vccd1 _21646_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19261__B1 _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19680_ _19681_/B _19681_/A vssd1 vssd1 vccd1 vccd1 _19798_/A sky130_fd_sc_hd__and2b_1
X_16892_ _16890_/A _16890_/Y _16891_/Y _16823_/X vssd1 vssd1 vccd1 vccd1 _16903_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18631_ _18632_/A _18632_/B _18632_/C vssd1 vssd1 vccd1 vccd1 _18631_/X sky130_fd_sc_hd__o21a_2
X_15843_ _15706_/A _15705_/A _15705_/B _15701_/B _15701_/A vssd1 vssd1 vccd1 vccd1
+ _15844_/B sky130_fd_sc_hd__o32ai_4
XFILLER_0_99_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18562_ _18564_/A _18564_/B _18564_/C vssd1 vssd1 vccd1 vccd1 _18563_/A sky130_fd_sc_hd__a21oi_2
X_15774_ _16031_/A _15775_/B vssd1 vssd1 vccd1 vccd1 _15776_/A sky130_fd_sc_hd__nand2_2
XTAP_3550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12986_ _12986_/A _12986_/B vssd1 vssd1 vccd1 vccd1 _12988_/B sky130_fd_sc_hd__xnor2_1
XTAP_3561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17513_ _17513_/A _17513_/B _17513_/C vssd1 vssd1 vccd1 vccd1 _17514_/A sky130_fd_sc_hd__and3_2
XTAP_3583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14725_ _14568_/A _14568_/C _14568_/B vssd1 vssd1 vccd1 vccd1 _14730_/A sky130_fd_sc_hd__a21bo_1
XTAP_3594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18493_ _19438_/A _19438_/B _19414_/C _19866_/D vssd1 vssd1 vccd1 vccd1 _18493_/X
+ sky130_fd_sc_hd__and4_1
X_11937_ _11938_/A _11938_/B vssd1 vssd1 vccd1 vccd1 _11960_/A sky130_fd_sc_hd__nand2b_1
XTAP_2860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21371__A1 _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16409__A _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17444_ _17915_/A _19587_/A _17443_/D _17657_/A vssd1 vssd1 vccd1 vccd1 _17445_/B
+ sky130_fd_sc_hd__a22oi_1
X_14656_ _15961_/D _15653_/C _15112_/D _15838_/D vssd1 vssd1 vccd1 vccd1 _14656_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11868_ _11869_/A _11869_/B vssd1 vssd1 vccd1 vccd1 _11889_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15032__B _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13607_ _13604_/Y _13605_/X _13446_/X _13448_/X vssd1 vssd1 vccd1 vccd1 _13643_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_83_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10819_ hold203/A hold215/A vssd1 vssd1 vccd1 vccd1 _10821_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17375_ _21142_/A _12493_/B _21337_/B _20770_/B vssd1 vssd1 vccd1 vccd1 _17375_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_138_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14587_ _14587_/A _14587_/B vssd1 vssd1 vccd1 vccd1 _14588_/B sky130_fd_sc_hd__xor2_4
X_11799_ _11799_/A _11799_/B vssd1 vssd1 vccd1 vccd1 _11801_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__11052__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18624__A _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19114_ _19112_/X _19114_/B vssd1 vssd1 vccd1 vccd1 _19115_/B sky130_fd_sc_hd__and2b_1
X_16326_ _16326_/A _16418_/A _16396_/B _16418_/B vssd1 vssd1 vccd1 vccd1 _16327_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_83_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13538_ _13538_/A vssd1 vssd1 vccd1 vccd1 _13538_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19439__B _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14871__B _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15889__B1 _10959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19045_ _19176_/B _19045_/B vssd1 vssd1 vccd1 vccd1 _19046_/B sky130_fd_sc_hd__nor2_1
XANTENNA__12094__D _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13469_ _14713_/B _13913_/C _14077_/B _14713_/A vssd1 vssd1 vccd1 vccd1 _13470_/B
+ sky130_fd_sc_hd__a22o_1
X_16257_ fanout9/A _21142_/B vssd1 vssd1 vccd1 vccd1 _16257_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15208_ _14918_/B _15207_/Y _15205_/X vssd1 vssd1 vccd1 vccd1 _15209_/B sky130_fd_sc_hd__o21ba_2
XFILLER_0_51_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16188_ _16070_/B _16071_/Y _16303_/A _16187_/X vssd1 vssd1 vccd1 vccd1 _16303_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_112_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15139_ _15282_/B _15138_/B _15138_/C vssd1 vssd1 vccd1 vccd1 _15140_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19947_ hold89/X _19946_/Y fanout4/X vssd1 vssd1 vccd1 vccd1 _21906_/D sky130_fd_sc_hd__mux2_1
Xclkbuf_2_3__f_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3__f_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__19185__A_N _17854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11678__A1 _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11678__B2 _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19878_ _19877_/B _19877_/C _19877_/A vssd1 vssd1 vccd1 vccd1 _19879_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_65_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18829_ _18826_/Y _18827_/X _18676_/Y _18678_/X vssd1 vssd1 vccd1 vccd1 _18830_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14616__A1 _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21840_ _21845_/CLK _21840_/D vssd1 vssd1 vccd1 vccd1 _21840_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12269__D _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21771_ _21789_/CLK _21771_/D vssd1 vssd1 vccd1 vccd1 _21771_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__21362__A1 _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout256_A _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20722_ _20721_/D _21293_/B _21261_/B _20590_/D vssd1 vssd1 vccd1 vccd1 _20723_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_148_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17141__C _17141_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20653_ _20774_/A _20774_/B hold294/A _21056_/B vssd1 vssd1 vccd1 vccd1 _20654_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA_fanout423_A _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20584_ _20719_/A vssd1 vssd1 vccd1 vccd1 _20586_/D sky130_fd_sc_hd__inv_2
XANTENNA__18190__A1_N _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19068__C _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21417__A2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21205_ _21206_/B vssd1 vssd1 vccd1 vccd1 _21205_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18294__A1 _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18294__B2 _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11629__C _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21136_ _21137_/A _21137_/B vssd1 vssd1 vccd1 vccd1 _21253_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11118__A0 _10972_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout420 _21765_/Q vssd1 vssd1 vccd1 vccd1 _15076_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__14855__A1 _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout431 _12780_/B vssd1 vssd1 vccd1 vccd1 _12242_/B sky130_fd_sc_hd__clkbuf_4
Xfanout442 _21760_/Q vssd1 vssd1 vccd1 vccd1 _14572_/A sky130_fd_sc_hd__clkbuf_8
Xfanout453 hold313/A vssd1 vssd1 vccd1 vccd1 _16173_/B sky130_fd_sc_hd__clkbuf_8
X_21067_ _21067_/A _21067_/B vssd1 vssd1 vccd1 vccd1 _21069_/B sky130_fd_sc_hd__xor2_1
Xfanout464 _21753_/Q vssd1 vssd1 vccd1 vccd1 _15510_/B sky130_fd_sc_hd__clkbuf_4
Xfanout475 _15093_/B vssd1 vssd1 vccd1 vccd1 _16268_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__18597__A2 _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout486 _21747_/Q vssd1 vssd1 vccd1 vccd1 _14384_/D sky130_fd_sc_hd__clkbuf_8
XANTENNA__19794__B2 _11550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20018_ _19915_/Y _19917_/X _20168_/A _20017_/X vssd1 vssd1 vccd1 vccd1 _20168_/B
+ sky130_fd_sc_hd__o211ai_2
Xfanout497 _21745_/Q vssd1 vssd1 vccd1 vccd1 _16404_/A sky130_fd_sc_hd__buf_4
XANTENNA__11645__B _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15804__B1 _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12840_ _13822_/B _14176_/C _13402_/D _13983_/B vssd1 vssd1 vccd1 vccd1 _12842_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14083__A2 _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13860__B _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ _13155_/A _14195_/A _12771_/C _21765_/Q vssd1 vssd1 vccd1 vccd1 _12896_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__17332__B _18058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21353__A1 _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21969_ _21974_/CLK _21969_/D vssd1 vssd1 vccd1 vccd1 hold301/A sky130_fd_sc_hd__dfxtp_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14510_ _14506_/X _14508_/Y _14353_/X _14356_/X vssd1 vssd1 vccd1 vccd1 _14511_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ _11722_/A _11722_/B vssd1 vssd1 vccd1 vccd1 _11723_/B sky130_fd_sc_hd__nor2_1
X_15490_ _15490_/A _15490_/B vssd1 vssd1 vccd1 vccd1 _15491_/B sky130_fd_sc_hd__and2_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14441_ _14442_/A _14442_/B vssd1 vssd1 vccd1 vccd1 _14441_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_83_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11653_ _11585_/A _11585_/B _11592_/X vssd1 vssd1 vccd1 vccd1 _11799_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout60 _21407_/S vssd1 vssd1 vccd1 vccd1 _21420_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__18444__A _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout71 hold329/X vssd1 vssd1 vccd1 vccd1 _19179_/C sky130_fd_sc_hd__buf_4
XFILLER_0_153_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14372_ _14198_/A _14198_/C _14198_/B vssd1 vssd1 vccd1 vccd1 _14373_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_92_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17160_ _17117_/A _17117_/B _17117_/C vssd1 vssd1 vccd1 vccd1 _17160_/Y sky130_fd_sc_hd__a21oi_1
Xfanout82 _21846_/Q vssd1 vssd1 vccd1 vccd1 _19030_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout93 _19051_/C vssd1 vssd1 vccd1 vccd1 _18732_/C sky130_fd_sc_hd__clkbuf_8
X_11584_ _12426_/B _12511_/A _11583_/B _11580_/X vssd1 vssd1 vccd1 vccd1 _11585_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16111_ _16112_/A _16112_/B vssd1 vssd1 vccd1 vccd1 _16111_/Y sky130_fd_sc_hd__nand2_1
X_13323_ _13323_/A _13323_/B vssd1 vssd1 vccd1 vccd1 _13332_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17091_ _17091_/A _17091_/B _17091_/C vssd1 vssd1 vccd1 vccd1 _17099_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_51_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16042_ _16424_/A _16377_/A _16042_/C _16213_/A vssd1 vssd1 vccd1 vccd1 _16213_/B
+ sky130_fd_sc_hd__nand4_1
X_13254_ _14138_/A _14463_/D _13402_/D vssd1 vssd1 vccd1 vccd1 _13254_/X sky130_fd_sc_hd__and3_1
XFILLER_0_0_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13897__A2 _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12205_ _12160_/X _12177_/Y _12203_/A _12202_/Y vssd1 vssd1 vccd1 vccd1 _12207_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_60_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17088__A2 _17086_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13185_ _14572_/A _13913_/C vssd1 vssd1 vccd1 vccd1 _13188_/A sky130_fd_sc_hd__and2_1
XFILLER_0_103_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19801_ _20026_/B _20838_/C _20838_/D _20178_/D vssd1 vssd1 vccd1 vccd1 _19804_/C
+ sky130_fd_sc_hd__a22o_1
X_12136_ _12269_/A _12245_/B _12530_/A _12512_/A vssd1 vssd1 vccd1 vccd1 _12139_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11109__A0 _10912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17993_ _17991_/X _17993_/B vssd1 vssd1 vccd1 vccd1 _17995_/A sky130_fd_sc_hd__nand2b_1
X_19732_ _19732_/A _19732_/B _20249_/B _20247_/C vssd1 vssd1 vccd1 vccd1 _19849_/A
+ sky130_fd_sc_hd__nand4_2
X_16944_ _16933_/A _16933_/C _16933_/B vssd1 vssd1 vccd1 vccd1 _16946_/C sky130_fd_sc_hd__a21oi_1
X_12067_ _12011_/A _12011_/C _12011_/B vssd1 vssd1 vccd1 vccd1 _12067_/X sky130_fd_sc_hd__a21o_1
XANTENNA__14212__A _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11018_ mstream_o[92] hold44/X _11027_/S vssd1 vssd1 vccd1 vccd1 _21629_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12321__A2 _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11555__B _11555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19663_ _20590_/D _20733_/C _20606_/D _19664_/B vssd1 vssd1 vccd1 vccd1 _19666_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16875_ _16806_/A _16806_/B _16806_/C vssd1 vssd1 vccd1 vccd1 _16876_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13473__D _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20395__A2 _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18619__A _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18614_ _18610_/Y _18611_/X _18454_/A _18454_/Y vssd1 vssd1 vccd1 vccd1 _18674_/B
+ sky130_fd_sc_hd__a211oi_2
X_15826_ _15650_/B _15689_/Y _15823_/X _15824_/Y vssd1 vssd1 vccd1 vccd1 _15826_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__12609__B1 _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13681__A1_N _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19594_ _19591_/X _19593_/Y _19444_/A _19847_/A vssd1 vssd1 vccd1 vccd1 _19597_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_56_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14074__A2 _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18338__B _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18545_ _19008_/D _18857_/B _19179_/C vssd1 vssd1 vccd1 vccd1 _18545_/X sky130_fd_sc_hd__and3_1
XTAP_3380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15757_ _15622_/Y _15626_/B _15624_/B vssd1 vssd1 vccd1 vccd1 _15758_/B sky130_fd_sc_hd__o21ai_2
XTAP_3391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12969_ _12969_/A _12969_/B vssd1 vssd1 vccd1 vccd1 _12971_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__21344__A1 _21349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14708_ _14707_/B _14707_/C _14707_/A vssd1 vssd1 vccd1 vccd1 _14709_/B sky130_fd_sc_hd__a21oi_1
X_18476_ _18478_/A _18478_/B _18478_/C vssd1 vssd1 vccd1 vccd1 _18476_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_47_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15688_ _15687_/B _15687_/C _15687_/A vssd1 vssd1 vccd1 vccd1 _15689_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_129_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17427_ _17427_/A _17427_/B _17427_/C vssd1 vssd1 vccd1 vccd1 _17427_/Y sky130_fd_sc_hd__nand3_4
X_14639_ _14638_/B _14785_/B _14638_/A vssd1 vssd1 vccd1 vccd1 _14640_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_7_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15574__A2 _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11721__D _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17358_ _17256_/C _17255_/Y _17356_/X _17357_/Y vssd1 vssd1 vccd1 vccd1 _17360_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19169__B _19169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16309_ _16309_/A _16309_/B vssd1 vssd1 vccd1 vccd1 _16311_/B sky130_fd_sc_hd__or2_1
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21211__C _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17289_ _17290_/A _17290_/B vssd1 vssd1 vccd1 vccd1 _17404_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_71_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16305__C _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14534__B1 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19028_ _19028_/A _19028_/B vssd1 vssd1 vccd1 vccd1 _19035_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11348__A0 _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18801__B _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16602__A _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17417__B _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19225__B1 _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17787__B1 _17670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout373_A _21775_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16975__C _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17433__A _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19351__C _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19528__A1 _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19528__B2 _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21823_ _21829_/CLK _21823_/D vssd1 vssd1 vccd1 vccd1 _21823_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_149_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout540_A _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21335__A1 _21349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout638_A fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21754_ _22049_/CLK _21754_/D vssd1 vssd1 vccd1 vccd1 _21754_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_78_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20794__A _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20705_ _20705_/A _20705_/B vssd1 vssd1 vccd1 vccd1 _20707_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_93_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21685_ _22069_/CLK _21685_/D vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20636_ _20468_/B _20471_/A _20634_/Y _20635_/X vssd1 vssd1 vccd1 vccd1 _20638_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15317__A2 _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20567_ _20567_/A _20567_/B vssd1 vssd1 vccd1 vccd1 _20569_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__17711__B1 _21346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16215__C _16396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11339__B1 _11338_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20498_ _20498_/A _20498_/B _20498_/C vssd1 vssd1 vccd1 vccd1 _20499_/D sky130_fd_sc_hd__nor3_2
XANTENNA__12843__A1_N _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18711__B _19493_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17608__A _19337_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16512__A _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16817__A2 _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21119_ _21188_/B _21117_/X _20955_/X _20958_/Y vssd1 vssd1 vccd1 vccd1 _21119_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19823__A _19823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14990_ _14990_/A _14990_/B _14990_/C vssd1 vssd1 vccd1 vccd1 _15012_/B sky130_fd_sc_hd__and3_2
XFILLER_0_121_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22099_ _22105_/CLK _22099_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[35] sky130_fd_sc_hd__dfrtp_4
Xfanout250 _20583_/A vssd1 vssd1 vccd1 vccd1 _20975_/D sky130_fd_sc_hd__buf_4
XANTENNA__20969__A _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12303__A2 _12402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout261 _19823_/A vssd1 vssd1 vccd1 vccd1 _20721_/D sky130_fd_sc_hd__buf_4
Xfanout272 _21801_/Q vssd1 vssd1 vccd1 vccd1 _17417_/A sky130_fd_sc_hd__buf_4
X_13941_ _13790_/B _13790_/Y _13938_/X _13940_/Y vssd1 vssd1 vccd1 vccd1 _13941_/X
+ sky130_fd_sc_hd__a211o_1
Xfanout283 _17520_/B vssd1 vssd1 vccd1 vccd1 _16917_/C sky130_fd_sc_hd__buf_4
Xfanout294 _17619_/B vssd1 vssd1 vccd1 vccd1 _16743_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__21574__A1 _11055_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16660_ _17145_/A _17526_/B vssd1 vssd1 vccd1 vccd1 _16662_/B sky130_fd_sc_hd__and2_1
X_13872_ _13875_/B _14024_/B _14516_/A _14365_/C _13724_/X vssd1 vssd1 vccd1 vccd1
+ _13881_/A sky130_fd_sc_hd__a41o_1
XFILLER_0_69_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15611_ _15608_/Y _15609_/X _15469_/B _15469_/Y vssd1 vssd1 vccd1 vccd1 _15612_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_0_clk_i_A _21822_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12823_ _12947_/B _12947_/C _12822_/C vssd1 vssd1 vccd1 vccd1 _12824_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__21326__A1 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16591_ _16989_/C _17520_/A vssd1 vssd1 vccd1 vccd1 _16595_/A sky130_fd_sc_hd__nand2_1
XANTENNA__20129__A2 _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18330_ _18176_/X _18178_/X _18327_/X _18328_/Y vssd1 vssd1 vccd1 vccd1 _18330_/Y
+ sky130_fd_sc_hd__o211ai_4
X_15542_ _15543_/A _15543_/B vssd1 vssd1 vccd1 vccd1 _15727_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_139_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12754_ _12754_/A _12754_/B vssd1 vssd1 vccd1 vccd1 _12764_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_16_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17997__B _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18261_ _18261_/A _18261_/B vssd1 vssd1 vccd1 vccd1 _18263_/B sky130_fd_sc_hd__xor2_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11705_ _11705_/A _11705_/B vssd1 vssd1 vccd1 vccd1 _11718_/A sky130_fd_sc_hd__nand2_1
X_15473_ _15473_/A _15473_/B _15473_/C vssd1 vssd1 vccd1 vccd1 _15475_/C sky130_fd_sc_hd__nand3_4
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12685_ _12684_/A _12684_/B _12684_/C vssd1 vssd1 vccd1 vccd1 _12687_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_38_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17212_ _17213_/B _17213_/A vssd1 vssd1 vccd1 vccd1 _17212_/X sky130_fd_sc_hd__and2b_1
X_14424_ _14260_/A _14260_/C _14260_/B vssd1 vssd1 vccd1 vccd1 _14426_/B sky130_fd_sc_hd__a21bo_2
XFILLER_0_126_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11636_ _11793_/A _11635_/B _11632_/X vssd1 vssd1 vccd1 vccd1 _11652_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_65_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18192_ _18193_/A _18332_/B _18192_/C vssd1 vssd1 vccd1 vccd1 _18328_/A sky130_fd_sc_hd__or3_1
XFILLER_0_53_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16406__B _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17143_ _17145_/A _17146_/D _17142_/X _17141_/X vssd1 vssd1 vccd1 vccd1 _17149_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_64_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14355_ _14813_/A _15022_/B _14357_/C _14357_/D vssd1 vssd1 vccd1 vccd1 _14355_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11567_ _11573_/A _11573_/B vssd1 vssd1 vccd1 vccd1 _11610_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_52_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13306_ _13306_/A _13306_/B _13306_/C vssd1 vssd1 vccd1 vccd1 _13306_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_123_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14286_ _14289_/A _14289_/B vssd1 vssd1 vccd1 vccd1 _14288_/A sky130_fd_sc_hd__or2_2
X_17074_ _17074_/A _17074_/B vssd1 vssd1 vccd1 vccd1 _17075_/B sky130_fd_sc_hd__or2_1
X_11498_ _11498_/A1 t1y[16] t0x[16] _11507_/B2 vssd1 vssd1 vccd1 vccd1 _11498_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_40_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13468__D _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16025_ _16363_/A hold117/A _10965_/Y fanout5/X _16024_/Y vssd1 vssd1 vccd1 vccd1
+ _16025_/X sky130_fd_sc_hd__a221o_1
X_13237_ _13237_/A _13376_/B _13237_/C vssd1 vssd1 vccd1 vccd1 _13237_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_122_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13168_ _13168_/A _13168_/B vssd1 vssd1 vccd1 vccd1 _13204_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17237__B _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _12120_/A _12120_/B _12120_/C vssd1 vssd1 vccd1 vccd1 _12127_/A sky130_fd_sc_hd__o21ai_1
X_13099_ _13381_/C _13394_/A _14155_/C _14155_/D vssd1 vssd1 vccd1 vccd1 _13240_/A
+ sky130_fd_sc_hd__and4_2
X_17976_ _18857_/B _19030_/C _21847_/Q _18703_/A vssd1 vssd1 vccd1 vccd1 _17978_/A
+ sky130_fd_sc_hd__a22oi_1
X_19715_ _19715_/A _19715_/B _19715_/C vssd1 vssd1 vccd1 vccd1 _19715_/Y sky130_fd_sc_hd__nand3_1
X_16927_ _17096_/A _17019_/C vssd1 vssd1 vccd1 vccd1 _16928_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18349__A _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17233__A2 _17666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19646_ _19810_/D _20841_/B vssd1 vssd1 vccd1 vccd1 _19647_/B sky130_fd_sc_hd__nand2_1
X_16858_ _16851_/A _16851_/B _16851_/C vssd1 vssd1 vccd1 vccd1 _16859_/B sky130_fd_sc_hd__a21o_1
X_15809_ _15809_/A _15927_/B vssd1 vssd1 vccd1 vccd1 _15811_/B sky130_fd_sc_hd__or2_1
XFILLER_0_149_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19577_ _19573_/X _19575_/Y _19415_/Y _19417_/X vssd1 vssd1 vccd1 vccd1 _19578_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16789_ _16789_/A _16790_/A _16789_/C vssd1 vssd1 vccd1 vccd1 _17165_/A sky130_fd_sc_hd__nand3_4
XANTENNA__12397__A _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18528_ _18525_/Y _18526_/X _18377_/C _18378_/X vssd1 vssd1 vccd1 vccd1 _18529_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18459_ _18305_/A _18305_/Y _18456_/X _18457_/Y vssd1 vssd1 vccd1 vccd1 _18459_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_75_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13558__A1 _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13558__B2 _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21470_ hold153/X sstream_i[47] _21494_/S vssd1 vssd1 vccd1 vccd1 _21997_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20421_ _20421_/A _20421_/B vssd1 vssd1 vccd1 vccd1 _20423_/B sky130_fd_sc_hd__or2_1
XFILLER_0_132_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19908__A _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11240__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout219_A _18789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20352_ _20352_/A _20352_/B vssd1 vssd1 vccd1 vccd1 _20354_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12860__A _13554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20283_ _20562_/B _21153_/B _21264_/B _20689_/A vssd1 vssd1 vccd1 vccd1 _20287_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22022_ _22038_/CLK _22022_/D vssd1 vssd1 vccd1 vccd1 hold298/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout490_A _21746_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout588_A _11549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20147__A1_N _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20004__D _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold69 hold69/A vssd1 vssd1 vccd1 vccd1 hold69/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21806_ _21806_/CLK _21806_/D vssd1 vssd1 vccd1 vccd1 _21806_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout34_A _21490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21737_ _21803_/CLK _21737_/D vssd1 vssd1 vccd1 vccd1 _21737_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16735__B2 _16734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16507__A _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20674__D _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12470_ _12471_/A _12471_/B _12471_/C vssd1 vssd1 vccd1 vccd1 _12470_/X sky130_fd_sc_hd__and3_1
XFILLER_0_152_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21668_ _21906_/CLK _21668_/D vssd1 vssd1 vccd1 vccd1 hold68/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11421_ hold305/A fanout28/X _11420_/X vssd1 vssd1 vccd1 vccd1 _11421_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15130__B _16284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12152__A1_N _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20619_ _20485_/Y _20487_/Y _20617_/X _20618_/Y vssd1 vssd1 vccd1 vccd1 _20621_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_152_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19685__B1 _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14027__A _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21599_ _21934_/CLK _21599_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[62] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11150__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14140_ _14312_/D _16404_/B vssd1 vssd1 vccd1 vccd1 _14141_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12782__A1_N _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11352_ hold319/X _11351_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21789_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12772__A2 _12771_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19537__B _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15171__B1 _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14071_ _14070_/B _14070_/C _14070_/A vssd1 vssd1 vccd1 vccd1 _14072_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13866__A _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11283_ fanout58/X v0z[14] fanout17/X _11282_/X vssd1 vssd1 vccd1 vccd1 _11283_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17338__A _17557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19437__B1 _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13022_ _12884_/A _12884_/C _12884_/B vssd1 vssd1 vccd1 vccd1 _13023_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__13721__A1 _13875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13721__B2 _13877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17830_ _17830_/A _17830_/B _17837_/B vssd1 vssd1 vccd1 vccd1 _17831_/B sky130_fd_sc_hd__or3_1
X_17761_ _17761_/A _17761_/B vssd1 vssd1 vccd1 vccd1 _17770_/A sky130_fd_sc_hd__xor2_1
X_14973_ _14974_/A _14974_/B vssd1 vssd1 vccd1 vccd1 _15502_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_22_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19500_ _19501_/A _19501_/B vssd1 vssd1 vccd1 vccd1 _19502_/A sky130_fd_sc_hd__nor2_1
XANTENNA__19703__D _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16712_ _16715_/B _16712_/B _16712_/C _16712_/D vssd1 vssd1 vccd1 vccd1 _16712_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_57_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13924_ _13924_/A _13924_/B vssd1 vssd1 vccd1 vccd1 _13933_/A sky130_fd_sc_hd__nor2_1
X_17692_ _17689_/X _17690_/Y _17575_/C _17574_/Y vssd1 vssd1 vccd1 vccd1 _17693_/D
+ sky130_fd_sc_hd__a211o_1
XANTENNA__17504__C _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19431_ _19432_/A _19751_/C _19432_/C _19598_/A vssd1 vssd1 vccd1 vccd1 _19433_/B
+ sky130_fd_sc_hd__a22o_1
X_16643_ _16642_/A _16642_/C _16642_/B vssd1 vssd1 vccd1 vccd1 _16645_/B sky130_fd_sc_hd__a21o_1
X_13855_ _13695_/Y _13698_/X _13972_/A _13854_/X vssd1 vssd1 vccd1 vccd1 _13972_/B
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__18319__D _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16974__A1 _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16974__B2 _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19362_ _19519_/B _19362_/B vssd1 vssd1 vccd1 vccd1 _19365_/A sky130_fd_sc_hd__nand2b_1
X_12806_ _12803_/X _12804_/Y _12692_/C _12691_/Y vssd1 vssd1 vccd1 vccd1 _12807_/D
+ sky130_fd_sc_hd__a211o_1
X_16574_ _17520_/B _17417_/C _16899_/B _17874_/A vssd1 vssd1 vccd1 vccd1 _16575_/D
+ sky130_fd_sc_hd__a22o_1
X_13786_ _13632_/A _13632_/C _13632_/B vssd1 vssd1 vccd1 vccd1 _13787_/C sky130_fd_sc_hd__a21bo_1
X_10998_ mstream_o[72] hold40/X _11005_/S vssd1 vssd1 vccd1 vccd1 _21609_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_146_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18313_ _19686_/A _19686_/B _18929_/B _18616_/D vssd1 vssd1 vccd1 vccd1 _18314_/D
+ sky130_fd_sc_hd__nand4_2
XANTENNA__18616__B _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15525_ _16036_/A _15525_/B vssd1 vssd1 vccd1 vccd1 _15648_/B sky130_fd_sc_hd__nor2_1
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16726__A1 _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17520__B _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19293_ _19130_/A _19130_/C _19130_/B vssd1 vssd1 vccd1 vccd1 _19295_/B sky130_fd_sc_hd__a21bo_1
X_12737_ _12639_/C _12641_/A _12856_/B _12736_/X vssd1 vssd1 vccd1 vccd1 _12868_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_57_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20522__A2 _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16726__B2 _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18244_ _18100_/B _18242_/Y _18394_/B _17969_/A vssd1 vssd1 vccd1 vccd1 _18245_/B
+ sky130_fd_sc_hd__o22a_2
XFILLER_0_38_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15456_ _15587_/A _15978_/B _15961_/D _15456_/D vssd1 vssd1 vccd1 vccd1 _15587_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_128_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12668_ _13173_/C _12780_/B _13034_/D _12780_/A vssd1 vssd1 vccd1 vccd1 _12668_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_154_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14407_ _14859_/A _15091_/C _14408_/C _14554_/A vssd1 vssd1 vccd1 vccd1 _14409_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18175_ _18175_/A _18175_/B vssd1 vssd1 vccd1 vccd1 _18177_/B sky130_fd_sc_hd__and2_1
X_11619_ _11588_/A _11591_/A _11615_/X _11617_/Y vssd1 vssd1 vccd1 vccd1 _12316_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_53_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15387_ _15385_/Y _15386_/X _15224_/Y _15248_/Y vssd1 vssd1 vccd1 vccd1 _15426_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11060__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12599_ _12957_/A vssd1 vssd1 vccd1 vccd1 _12600_/B sky130_fd_sc_hd__inv_2
XFILLER_0_142_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17126_ _17145_/A _17493_/A _17126_/C _17126_/D vssd1 vssd1 vccd1 vccd1 _17140_/A
+ sky130_fd_sc_hd__and4_1
X_14338_ _14162_/X _14338_/B vssd1 vssd1 vccd1 vccd1 _14340_/B sky130_fd_sc_hd__and2b_2
XFILLER_0_123_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21619__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13776__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17057_ _17029_/A _17146_/C _17146_/D _17029_/B vssd1 vssd1 vccd1 vccd1 _17058_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14269_ _14268_/B _14268_/C _14268_/A vssd1 vssd1 vccd1 vccd1 _14269_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_64_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16008_ _15844_/A _15844_/B _15847_/A vssd1 vssd1 vccd1 vccd1 _16010_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18651__A1 _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17959_ _17958_/B _17958_/C _17958_/A vssd1 vssd1 vccd1 vccd1 _17959_/Y sky130_fd_sc_hd__a21oi_2
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18403__A1 _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20970_ _20970_/A _21085_/B vssd1 vssd1 vccd1 vccd1 _20972_/B sky130_fd_sc_hd__or2_1
XANTENNA__18403__B2 _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19600__B1 _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12839__B _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19629_ _19629_/A _19629_/B vssd1 vssd1 vccd1 vccd1 _19630_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout169_A _19732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_671 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15231__A _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21522_ hold256/X sstream_i[99] _21528_/S vssd1 vssd1 vccd1 vccd1 _22049_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_134_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21453_ hold120/X sstream_i[30] _21507_/S vssd1 vssd1 vccd1 vccd1 _21980_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_17_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout503_A _21743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21379__S _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20404_ _21034_/A _20404_/B vssd1 vssd1 vccd1 vccd1 _20407_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21384_ _21720_/D _21384_/B vssd1 vssd1 vccd1 vccd1 _21384_/X sky130_fd_sc_hd__or2_1
XFILLER_0_71_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20335_ _20472_/A _21311_/B _20845_/D _20335_/D vssd1 vssd1 vccd1 vccd1 _20472_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_98_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20266_ _21261_/A _21264_/A _20267_/C _20473_/A vssd1 vssd1 vccd1 vccd1 _20268_/A
+ sky130_fd_sc_hd__a22o_1
X_22005_ _22005_/CLK _22005_/D vssd1 vssd1 vccd1 vccd1 hold164/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__19373__A _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold283_A hold283/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20197_ _20198_/A _20198_/B vssd1 vssd1 vccd1 vccd1 _20197_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__19092__B _19092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20312__A _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19198__A2 _19030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20669__D _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11970_ _11979_/A _11970_/B vssd1 vssd1 vccd1 vccd1 _11971_/C sky130_fd_sc_hd__and2_1
XANTENNA__17324__C _19430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10921_ hold20/A hold50/A vssd1 vssd1 vccd1 vccd1 _10923_/A sky130_fd_sc_hd__or2_1
XANTENNA__13571__D _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20966__B _21293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13640_ _13486_/B _13486_/Y _13637_/X _13639_/Y vssd1 vssd1 vccd1 vccd1 _13643_/C
+ sky130_fd_sc_hd__a211oi_4
X_10852_ _10859_/B _10852_/B vssd1 vssd1 vccd1 vccd1 _10852_/X sky130_fd_sc_hd__and2_2
XANTENNA_clkbuf_leaf_26_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ _13877_/A _14027_/A _14516_/A _14365_/C vssd1 vssd1 vccd1 vccd1 _13720_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_39_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15310_ _15449_/A _15310_/B vssd1 vssd1 vccd1 vccd1 _15311_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_82_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12522_ _12522_/A _12522_/B _12522_/C vssd1 vssd1 vccd1 vccd1 _12522_/Y sky130_fd_sc_hd__nor3_2
X_16290_ _16383_/S _16290_/B vssd1 vssd1 vccd1 vccd1 _16291_/B sky130_fd_sc_hd__xor2_1
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15241_ _15242_/A _15242_/B vssd1 vssd1 vccd1 vccd1 _15384_/B sky130_fd_sc_hd__or2_1
XANTENNA__19548__A _21839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12453_ _13155_/A _12780_/A _12780_/B _13155_/B vssd1 vssd1 vccd1 vccd1 _12455_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_87_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11404_ _11403_/X _17657_/A _11446_/S vssd1 vssd1 vccd1 vccd1 _21806_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_151_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15172_ _15961_/D _15838_/D _15717_/C _15976_/D vssd1 vssd1 vccd1 vccd1 _15316_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_90_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12384_ _12381_/Y _12382_/X _11669_/X _11671_/Y vssd1 vssd1 vccd1 vccd1 _12384_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__18171__B _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14123_ _14290_/A _14285_/B _14123_/C vssd1 vssd1 vccd1 vccd1 _14291_/B sky130_fd_sc_hd__and3_1
X_11335_ _21407_/S v0z[27] fanout20/X _11334_/X vssd1 vssd1 vccd1 vccd1 _11335_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_123_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19980_ _20098_/B _19979_/C _19979_/A vssd1 vssd1 vccd1 vccd1 _19980_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18931_ _18931_/A _18931_/B vssd1 vssd1 vccd1 vccd1 _18940_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_123_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14054_ _14384_/A _14212_/C _14212_/D _15763_/A vssd1 vssd1 vccd1 vccd1 _14054_/X
+ sky130_fd_sc_hd__a22o_1
X_11266_ _11502_/A1 t1x[10] v2z[10] _11501_/B2 _11265_/X vssd1 vssd1 vccd1 vccd1 _11266_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_24_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13005_ _12891_/Y _12895_/A _13003_/A _13004_/Y vssd1 vssd1 vccd1 vccd1 _13097_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_123_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18862_ _18863_/A _18863_/B vssd1 vssd1 vccd1 vccd1 _19024_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12005__A _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11197_ hold164/X fanout22/X _11196_/X vssd1 vssd1 vccd1 vccd1 _11197_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17813_ _17689_/C _17688_/Y _17810_/X _17811_/Y vssd1 vssd1 vccd1 vccd1 _17815_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_118_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18793_ _18793_/A _18793_/B vssd1 vssd1 vccd1 vccd1 _18813_/A sky130_fd_sc_hd__xor2_2
X_17744_ _17870_/B _17743_/C _17743_/A vssd1 vssd1 vccd1 vccd1 _17745_/B sky130_fd_sc_hd__a21o_1
X_14956_ _14956_/A _14956_/B _14956_/C vssd1 vssd1 vccd1 vccd1 _14956_/X sky130_fd_sc_hd__and3_2
XANTENNA__21037__B _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17234__C _17666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12659__B _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20607__A1_N _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13907_ _14051_/B _13906_/C _13906_/A vssd1 vssd1 vccd1 vccd1 _13907_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17675_ _17559_/A _17559_/C _17559_/B vssd1 vssd1 vccd1 vccd1 _17676_/C sky130_fd_sc_hd__a21bo_1
X_14887_ _14887_/A _14887_/B _14887_/C _14887_/D vssd1 vssd1 vccd1 vccd1 _14889_/A
+ sky130_fd_sc_hd__nor4_2
X_19414_ _19972_/A _20394_/B _19414_/C _19866_/D vssd1 vssd1 vccd1 vccd1 _19417_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_134_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16626_ _16625_/A _16625_/C _16625_/B vssd1 vssd1 vccd1 vccd1 _16629_/B sky130_fd_sc_hd__a21o_1
X_13838_ _13975_/B _16328_/B _13839_/C _13839_/D vssd1 vssd1 vccd1 vccd1 _13838_/Y
+ sky130_fd_sc_hd__a22oi_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19345_ _19345_/A _19345_/B vssd1 vssd1 vccd1 vccd1 _19346_/B sky130_fd_sc_hd__and2_1
XFILLER_0_18_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16557_ _16554_/X _16557_/B vssd1 vssd1 vccd1 vccd1 _16644_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_31_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13769_ _13767_/X _13769_/B vssd1 vssd1 vccd1 vccd1 _13770_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_130_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15508_ _15892_/A _15632_/B _16369_/B _16177_/B vssd1 vssd1 vccd1 vccd1 _15670_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_70_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19276_ _19276_/A _19276_/B vssd1 vssd1 vccd1 vccd1 _19285_/A sky130_fd_sc_hd__nand2_1
X_16488_ _16495_/A vssd1 vssd1 vccd1 vccd1 _16489_/D sky130_fd_sc_hd__inv_2
XFILLER_0_45_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18227_ _18087_/C _18086_/Y _18225_/X _18226_/Y vssd1 vssd1 vccd1 vccd1 _18230_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_155_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15439_ _21735_/Q _15838_/B _16314_/D _15439_/D vssd1 vssd1 vccd1 vccd1 _15442_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_26_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18158_ _18157_/A _18157_/B _18143_/Y vssd1 vssd1 vccd1 vccd1 _18158_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_29_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold303 hold303/A vssd1 vssd1 vccd1 vccd1 hold303/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17109_ _17078_/X _17083_/Y _17106_/A _17120_/A vssd1 vssd1 vccd1 vccd1 _17110_/C
+ sky130_fd_sc_hd__a211o_1
Xhold314 hold314/A vssd1 vssd1 vccd1 vccd1 hold314/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold325 hold325/A vssd1 vssd1 vccd1 vccd1 hold325/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18089_ _17953_/B _17952_/Y _18087_/X _18088_/Y vssd1 vssd1 vccd1 vccd1 _18091_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_29_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18872__A1 _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20120_ _20121_/A _20121_/B vssd1 vssd1 vccd1 vccd1 _20120_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_106_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14623__A2_N _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20051_ _20051_/A _20186_/A _20051_/C vssd1 vssd1 vccd1 vccd1 _20186_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12560__D _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16610__A _21822_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout286_A _18010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14768__C _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_209 hold275/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20953_ _20953_/A vssd1 vssd1 vccd1 vccd1 _20953_/Y sky130_fd_sc_hd__inv_2
XANTENNA_fanout453_A hold313/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20884_ _20885_/A _20885_/B vssd1 vssd1 vccd1 vccd1 _21016_/B sky130_fd_sc_hd__and2_2
XFILLER_0_49_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14413__A2 _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18256__B _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12424__A1 _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout620_A _21717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13621__B1 _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19352__A2 _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12975__A2 _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14177__A1 _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21505_ hold281/X sstream_i[82] _21507_/S vssd1 vssd1 vccd1 vccd1 _22032_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_17_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12735__D _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21436_ hold254/X sstream_i[13] _21442_/S vssd1 vssd1 vccd1 vccd1 _21963_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_72_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19087__B _19087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18312__B1 _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21367_ _21720_/D _21367_/B vssd1 vssd1 vccd1 vccd1 _21367_/X sky130_fd_sc_hd__or2_1
XFILLER_0_32_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11120_ _10984_/Y hold53/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21714_/D sky130_fd_sc_hd__mux2_1
XANTENNA__20026__B _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20670__A1 _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20318_ _20321_/B vssd1 vssd1 vccd1 vccd1 _20470_/A sky130_fd_sc_hd__inv_2
X_21298_ _21298_/A _21298_/B vssd1 vssd1 vccd1 vccd1 _21299_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__14024__B _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11051_ _11051_/A _11051_/B vssd1 vssd1 vccd1 vccd1 _11051_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_101_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18615__A1 _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20249_ _20249_/A _20249_/B vssd1 vssd1 vccd1 vccd1 _20250_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18615__B2 _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19812__B1 _10798_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19534__C _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13863__B _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14810_ _16092_/D _15653_/C _15112_/D _15961_/D vssd1 vssd1 vccd1 vccd1 _14810_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15790_ _15916_/B _16396_/A _16377_/B _15791_/A vssd1 vssd1 vccd1 vccd1 _15794_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_3721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14741_ _14742_/B _14742_/A vssd1 vssd1 vccd1 vccd1 _14741_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_93_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11953_ _11953_/A _12019_/A vssd1 vssd1 vccd1 vccd1 _11956_/B sky130_fd_sc_hd__or2_1
XTAP_3765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17460_ _17461_/A _17461_/B _17461_/C vssd1 vssd1 vccd1 vccd1 _17460_/X sky130_fd_sc_hd__and3_1
X_10904_ mstream_o[50] _10903_/Y _10992_/S vssd1 vssd1 vccd1 vccd1 _21587_/D sky130_fd_sc_hd__mux2_1
XTAP_3798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14672_ _15768_/A _16409_/A _14534_/X _14535_/X _16326_/A vssd1 vssd1 vccd1 vccd1
+ _14677_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_15_1108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11884_ _12319_/C _12420_/D _12302_/A _12312_/A vssd1 vssd1 vccd1 vccd1 _11969_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__14404__A2 _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16411_ _16411_/A _16411_/B vssd1 vssd1 vccd1 vccd1 _16412_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__18166__B _19230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13623_ _13623_/A _13623_/B vssd1 vssd1 vccd1 vccd1 _13632_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10835_ _10836_/B hold215/A hold203/A vssd1 vssd1 vccd1 vccd1 _10835_/Y sky130_fd_sc_hd__nand3b_1
X_17391_ _17489_/A _17391_/B vssd1 vssd1 vccd1 vccd1 _17405_/A sky130_fd_sc_hd__or2_1
XFILLER_0_156_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19130_ _19130_/A _19130_/B _19130_/C vssd1 vssd1 vccd1 vccd1 _19133_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_67_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16342_ _16343_/A _16343_/B vssd1 vssd1 vccd1 vccd1 _16342_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_39_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13554_ _13860_/A _13554_/B _13858_/C _16414_/A vssd1 vssd1 vccd1 vccd1 _13556_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21150__A2 _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19061_ _18897_/X _18900_/X _19058_/X _19060_/Y vssd1 vssd1 vccd1 vccd1 _19061_/X
+ sky130_fd_sc_hd__o211a_1
X_12505_ _12505_/A _12505_/B vssd1 vssd1 vccd1 vccd1 _12605_/B sky130_fd_sc_hd__xnor2_1
X_16273_ _16273_/A _16391_/B vssd1 vssd1 vccd1 vccd1 _16274_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_70_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13485_ _13486_/A _13486_/B _13486_/C vssd1 vssd1 vccd1 vccd1 _13485_/X sky130_fd_sc_hd__and3_1
XANTENNA__15021__D _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18012_ _18012_/A _18144_/B _18012_/C vssd1 vssd1 vccd1 vccd1 _18014_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_152_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15224_ _15225_/A _15225_/B vssd1 vssd1 vccd1 vccd1 _15224_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__12718__A2 _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12436_ _12437_/A _12437_/B _12437_/C vssd1 vssd1 vccd1 vccd1 _12436_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_63_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16414__B _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15155_ _15152_/Y _15305_/A _15155_/C _15698_/B vssd1 vssd1 vccd1 vccd1 _15305_/B
+ sky130_fd_sc_hd__and4bb_1
X_12367_ _12367_/A _12367_/B _12367_/C vssd1 vssd1 vccd1 vccd1 _12370_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14106_ _14105_/B _14105_/C _14105_/A vssd1 vssd1 vccd1 vccd1 _14106_/X sky130_fd_sc_hd__o21a_1
X_11318_ _11224_/A t1x[23] v2z[23] _11223_/A _11317_/X vssd1 vssd1 vccd1 vccd1 _11318_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_26_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11558__B _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15086_ _14974_/X _14984_/Y _14985_/X _15085_/A vssd1 vssd1 vccd1 vccd1 _15087_/C
+ sky130_fd_sc_hd__a31o_1
X_12298_ _12402_/B _12312_/A _11661_/B _11659_/X vssd1 vssd1 vccd1 vccd1 _12307_/A
+ sky130_fd_sc_hd__a31o_1
X_19963_ _19963_/A _20095_/B _19963_/C vssd1 vssd1 vccd1 vccd1 _19984_/A sky130_fd_sc_hd__and3_1
X_14037_ _21741_/Q _14365_/C _14037_/C _14190_/A vssd1 vssd1 vccd1 vccd1 _14190_/B
+ sky130_fd_sc_hd__nand4_2
X_11249_ _11122_/A t2y[6] t0y[6] _11123_/A vssd1 vssd1 vccd1 vccd1 _11249_/X sky130_fd_sc_hd__a22o_1
XANTENNA__17526__A _21802_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18914_ _18914_/A _18914_/B _18914_/C vssd1 vssd1 vccd1 vccd1 _18917_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19894_ _20416_/A _18773_/B _20416_/B _20863_/C vssd1 vssd1 vccd1 vccd1 _19898_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13773__B _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18845_ _18841_/A _18841_/B _18835_/Y vssd1 vssd1 vccd1 vccd1 _19001_/A sky130_fd_sc_hd__o21a_1
XANTENNA__16093__B2 _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18776_ _18624_/D _18625_/B _18774_/Y _18775_/X vssd1 vssd1 vccd1 vccd1 _18925_/A
+ sky130_fd_sc_hd__a211o_1
X_15988_ _15984_/Y _15986_/X _15856_/Y _15860_/A vssd1 vssd1 vccd1 vccd1 _15988_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_136_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17727_ _21795_/Q _19692_/C _19691_/D _19337_/D vssd1 vssd1 vccd1 vccd1 _17729_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19031__A1 _19650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14939_ _14939_/A _14939_/B vssd1 vssd1 vccd1 vccd1 _14940_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17899__C _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17658_ _17657_/A _19951_/A _19951_/B _20583_/A vssd1 vssd1 vccd1 vccd1 _17659_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16609_ _16608_/B _16608_/C _16608_/A vssd1 vssd1 vccd1 vccd1 _16615_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_148_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17589_ _17589_/A _17589_/B vssd1 vssd1 vccd1 vccd1 _17705_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_92_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17411__D _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19328_ _19214_/A _19214_/B _19212_/Y vssd1 vssd1 vccd1 vccd1 _19370_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21634__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11090__A0 _11043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13013__B _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19259_ _20103_/A _19705_/B vssd1 vssd1 vccd1 vccd1 _19260_/B sky130_fd_sc_hd__and2_1
XFILLER_0_143_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16605__A _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold100 hold100/A vssd1 vssd1 vccd1 vccd1 hold100/X sky130_fd_sc_hd__dlygate4sd3_1
X_21221_ _21222_/A _21222_/B _21222_/C vssd1 vssd1 vccd1 vccd1 _21275_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_41_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold111 hold111/A vssd1 vssd1 vccd1 vccd1 hold111/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold122 hold122/A vssd1 vssd1 vccd1 vccd1 hold122/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 hold133/A vssd1 vssd1 vccd1 vccd1 hold133/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold144 hold144/A vssd1 vssd1 vccd1 vccd1 hold144/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20652__A1 _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21152_ _21046_/B _21151_/X _21150_/X vssd1 vssd1 vccd1 vccd1 _21154_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__20652__B2 _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold155 hold155/A vssd1 vssd1 vccd1 vccd1 hold155/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 hold166/A vssd1 vssd1 vccd1 vccd1 hold166/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 hold177/A vssd1 vssd1 vccd1 vccd1 hold177/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 hold188/A vssd1 vssd1 vccd1 vccd1 hold188/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20103_ _20103_/A _21815_/Q _20103_/C _20282_/A vssd1 vssd1 vccd1 vccd1 _20282_/B
+ sky130_fd_sc_hd__nand4_1
Xfanout602 _11459_/B2 vssd1 vssd1 vccd1 vccd1 _11501_/B2 sky130_fd_sc_hd__buf_4
Xhold199 hold199/A vssd1 vssd1 vccd1 vccd1 hold199/X sky130_fd_sc_hd__dlygate4sd3_1
X_21083_ _21199_/A _21291_/B _21083_/C _21083_/D vssd1 vssd1 vccd1 vccd1 _21194_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_10_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout613 _21568_/S vssd1 vssd1 vccd1 vccd1 _21562_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout624 _17557_/A vssd1 vssd1 vccd1 vccd1 _18652_/A sky130_fd_sc_hd__clkbuf_4
Xfanout635 _21776_/Q vssd1 vssd1 vccd1 vccd1 _16380_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout646 nrst_i vssd1 vssd1 vccd1 vccd1 _21422_/A sky130_fd_sc_hd__buf_12
X_20034_ _20032_/D _20178_/B _21261_/B _19487_/B vssd1 vssd1 vccd1 vccd1 _20035_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20797__A _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_917 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11448__A2 _11124_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21985_ _22020_/CLK _21985_/D vssd1 vssd1 vccd1 vccd1 hold196/A sky130_fd_sc_hd__dfxtp_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19573__A2 _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20936_ _20936_/A _20936_/B vssd1 vssd1 vccd1 vccd1 _20937_/B sky130_fd_sc_hd__nand2_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11931__B _12403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20867_ _20868_/A _20868_/B vssd1 vssd1 vccd1 vccd1 _20869_/A sky130_fd_sc_hd__nand2_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20798_ _20931_/A vssd1 vssd1 vccd1 vccd1 _20800_/D sky130_fd_sc_hd__inv_2
XFILLER_0_9_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11081__A0 _10946_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19529__C _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13858__B _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13270_ _13864_/B _13269_/C _13269_/D _13867_/A vssd1 vssd1 vccd1 vccd1 _13270_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_51_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12221_ _12267_/A _12242_/B _12246_/D _12269_/C vssd1 vssd1 vccd1 vccd1 _12222_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__11659__A _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21419_ hold195/X _21418_/X _21421_/S vssd1 vssd1 vccd1 vccd1 _21948_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14035__A _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12152_ _12109_/C _12269_/D _12110_/A _12108_/Y vssd1 vssd1 vccd1 vccd1 _12153_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__17991__D _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11103_ _10867_/X hold31/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21697_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16960_ _16956_/B _16956_/C _16958_/X _16949_/Y vssd1 vssd1 vccd1 vccd1 _16961_/C
+ sky130_fd_sc_hd__a211o_1
X_12083_ _12083_/A _12083_/B vssd1 vssd1 vccd1 vccd1 _12130_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_120_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15911_ _15911_/A _16424_/A _15911_/C _16040_/C vssd1 vssd1 vccd1 vccd1 _16102_/A
+ sky130_fd_sc_hd__nand4_1
X_11034_ mstream_o[108] hold274/X _11039_/S vssd1 vssd1 vccd1 vccd1 _21645_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19261__A1 _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16891_ _16823_/A _16823_/B _16823_/C vssd1 vssd1 vccd1 vccd1 _16891_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_21_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19261__B2 _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18630_ _18630_/A _18630_/B vssd1 vssd1 vccd1 vccd1 _18632_/C sky130_fd_sc_hd__xor2_1
XANTENNA__17272__B1 _21334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15842_ _15842_/A _15966_/B vssd1 vssd1 vccd1 vccd1 _15844_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_21_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18561_ _18561_/A _18561_/B vssd1 vssd1 vccd1 vccd1 _18564_/C sky130_fd_sc_hd__xnor2_1
X_15773_ _15904_/B _15773_/B vssd1 vssd1 vccd1 vccd1 _15775_/B sky130_fd_sc_hd__nor2_1
XTAP_3540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12985_ _12986_/B _12986_/A vssd1 vssd1 vccd1 vccd1 _13104_/A sky130_fd_sc_hd__nand2b_1
XTAP_3551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15016__D _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17512_ _17512_/A _17512_/B _17512_/C vssd1 vssd1 vccd1 vccd1 _17513_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_58_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14724_ _14724_/A _14724_/B vssd1 vssd1 vccd1 vccd1 _14732_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18492_ _19723_/A _19262_/C vssd1 vssd1 vccd1 vccd1 _18496_/A sky130_fd_sc_hd__nand2_1
X_11936_ _11936_/A _11936_/B vssd1 vssd1 vccd1 vccd1 _11938_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21371__A2 _18842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16409__B _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17443_ _17915_/A _17657_/A _17666_/A _17443_/D vssd1 vssd1 vccd1 vccd1 _17445_/A
+ sky130_fd_sc_hd__and4_1
X_14655_ _14524_/A _14524_/B _14524_/C _14526_/X vssd1 vssd1 vccd1 vccd1 _14689_/A
+ sky130_fd_sc_hd__a31o_2
XTAP_2883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11867_ _11867_/A _11867_/B vssd1 vssd1 vccd1 vccd1 _11869_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13606_ _13446_/X _13448_/X _13604_/Y _13605_/X vssd1 vssd1 vccd1 vccd1 _13643_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_55_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10818_ hold227/A hold229/A vssd1 vssd1 vccd1 vccd1 _10836_/B sky130_fd_sc_hd__nor2_2
X_17374_ _17381_/C _17374_/B vssd1 vssd1 vccd1 vccd1 _21337_/B sky130_fd_sc_hd__xor2_4
XANTENNA__15032__C _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14586_ _14587_/A _14587_/B vssd1 vssd1 vccd1 vccd1 _14586_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_83_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11798_ _11771_/X _11796_/Y _11795_/Y _11795_/A vssd1 vssd1 vccd1 vccd1 _11801_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11072__A0 _10881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18624__B _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19113_ _19112_/B _19276_/B _19112_/A vssd1 vssd1 vccd1 vccd1 _19114_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_138_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16325_ _16418_/A _16396_/B _16418_/B _16326_/A vssd1 vssd1 vccd1 vccd1 _16327_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_40_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21331__A _21349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13537_ _13539_/A _13539_/B _13539_/C vssd1 vssd1 vccd1 vccd1 _13538_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12953__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20331__B1 _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15889__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14871__C _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15889__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19044_ _19174_/B _19043_/B _19176_/A _19043_/D vssd1 vssd1 vccd1 vccd1 _19045_/B
+ sky130_fd_sc_hd__o22a_1
X_16256_ _16256_/A _16256_/B vssd1 vssd1 vccd1 vccd1 _21142_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_140_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13468_ _14713_/A _14713_/B _13913_/C _14077_/B vssd1 vssd1 vccd1 vccd1 _13468_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_152_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15207_ _15207_/A vssd1 vssd1 vccd1 vccd1 _15207_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11569__A _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ _12415_/X _12416_/Y _12309_/Y _12312_/X vssd1 vssd1 vccd1 vccd1 _12479_/B
+ sky130_fd_sc_hd__a211oi_2
X_16187_ _16184_/X _16185_/Y _16032_/A _16035_/A vssd1 vssd1 vccd1 vccd1 _16187_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_140_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13399_ _13400_/A _13400_/B vssd1 vssd1 vccd1 vccd1 _13523_/B sky130_fd_sc_hd__and2_1
XANTENNA__18640__A _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11375__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15138_ _15282_/B _15138_/B _15138_/C vssd1 vssd1 vccd1 vccd1 _15253_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_50_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15069_ _15069_/A _15206_/B vssd1 vssd1 vccd1 vccd1 _15070_/B sky130_fd_sc_hd__xnor2_4
X_19946_ _19636_/A _15070_/B _19944_/Y _20770_/B _19945_/Y vssd1 vssd1 vccd1 vccd1
+ _19946_/Y sky130_fd_sc_hd__o221ai_1
XFILLER_0_26_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16160__A _16380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13296__A1_N _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11678__A2 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19877_ _19877_/A _19877_/B _19877_/C vssd1 vssd1 vccd1 vccd1 _19879_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_4_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18828_ _18676_/Y _18678_/X _18826_/Y _18827_/X vssd1 vssd1 vccd1 vccd1 _18830_/B
+ sky130_fd_sc_hd__a211oi_2
X_18759_ _18758_/B _18758_/C _18758_/A vssd1 vssd1 vccd1 vccd1 _18759_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17015__B1 _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15504__A _15907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21770_ _21789_/CLK _21770_/D vssd1 vssd1 vccd1 vccd1 _21770_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_72_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21362__A2 _18390_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20721_ _20590_/D _21293_/B _20721_/C _20721_/D vssd1 vssd1 vccd1 vccd1 _20855_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_93_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout151_A _21831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17141__D _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout249_A _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20652_ _20774_/B hold294/A _21056_/B _20774_/A vssd1 vssd1 vccd1 vccd1 _20654_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20583_ _20583_/A _20845_/D _21286_/B _21296_/B vssd1 vssd1 vccd1 vccd1 _20719_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_6_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout416_A _21766_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19068__D _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21204_ _21204_/A _21204_/B vssd1 vssd1 vccd1 vccd1 _21206_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__18294__A2 _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11629__D _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21135_ _21135_/A _21135_/B vssd1 vssd1 vccd1 vccd1 _21137_/B sky130_fd_sc_hd__or2_1
XFILLER_0_44_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout410 _15514_/A vssd1 vssd1 vccd1 vccd1 _15373_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__14855__A2 _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout421 _12897_/C vssd1 vssd1 vccd1 vccd1 _12229_/A sky130_fd_sc_hd__buf_4
Xfanout432 _21762_/Q vssd1 vssd1 vccd1 vccd1 _12780_/B sky130_fd_sc_hd__buf_4
X_21066_ _20949_/A _20949_/B _20946_/X vssd1 vssd1 vccd1 vccd1 _21067_/B sky130_fd_sc_hd__a21oi_1
Xfanout443 _12357_/C vssd1 vssd1 vccd1 vccd1 _12269_/B sky130_fd_sc_hd__buf_4
Xfanout454 hold313/A vssd1 vssd1 vccd1 vccd1 _16027_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__16057__A1 _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout465 _21753_/Q vssd1 vssd1 vccd1 vccd1 _16391_/B sky130_fd_sc_hd__clkbuf_8
Xfanout476 _15093_/B vssd1 vssd1 vccd1 vccd1 _16396_/A sky130_fd_sc_hd__clkbuf_4
X_20017_ _20125_/B _20015_/X _19879_/X _19885_/C vssd1 vssd1 vccd1 vccd1 _20017_/X
+ sky130_fd_sc_hd__a211o_1
Xfanout487 _21747_/Q vssd1 vssd1 vccd1 vccd1 _14218_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__19794__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout498 _14365_/D vssd1 vssd1 vccd1 vccd1 _13034_/D sky130_fd_sc_hd__buf_4
XANTENNA__15804__A1 _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout64_A _19185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15804__B2 _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12618__A1 _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13291__A1 _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ _14024_/B _12899_/B _12661_/X _12660_/X _12771_/C vssd1 vssd1 vccd1 vccd1
+ _12778_/A sky130_fd_sc_hd__a32o_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21968_ _21974_/CLK _21968_/D vssd1 vssd1 vccd1 vccd1 hold295/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__21353__A2 _17970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11721_ _13157_/A _12094_/A _12780_/B _13017_/A vssd1 vssd1 vccd1 vccd1 _11722_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20919_ _20918_/A _20787_/B _20788_/A vssd1 vssd1 vccd1 vccd1 _20920_/B sky130_fd_sc_hd__o21ba_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21899_ _21942_/CLK _21899_/D vssd1 vssd1 vccd1 vccd1 hold115/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11153__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14440_ _14277_/A _14277_/C _14277_/B vssd1 vssd1 vccd1 vccd1 _14442_/B sky130_fd_sc_hd__a21boi_4
XFILLER_0_49_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _11652_/A _11652_/B _11652_/C vssd1 vssd1 vccd1 vccd1 _11655_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_65_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_627 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout50 _11122_/X vssd1 vssd1 vccd1 vccd1 _11126_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11054__A0 _11053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout61 _10791_/Y vssd1 vssd1 vccd1 vccd1 _21407_/S sky130_fd_sc_hd__buf_6
XANTENNA__18444__B _19531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21151__A _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout72 _20838_/C vssd1 vssd1 vccd1 vccd1 _21286_/B sky130_fd_sc_hd__buf_4
X_14371_ _14370_/B _14370_/C _14370_/A vssd1 vssd1 vccd1 vccd1 _14373_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_36_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout83 _20733_/C vssd1 vssd1 vccd1 vccd1 _21283_/B sky130_fd_sc_hd__buf_4
XFILLER_0_153_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout94 fanout96/X vssd1 vssd1 vccd1 vccd1 _19051_/C sky130_fd_sc_hd__buf_4
XFILLER_0_25_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11583_ _11580_/X _11583_/B vssd1 vssd1 vccd1 vccd1 _11595_/B sky130_fd_sc_hd__and2b_1
XANTENNA__12773__A _13018_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16110_ _16110_/A _16110_/B vssd1 vssd1 vccd1 vccd1 _16112_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13322_ _13320_/X _13322_/B vssd1 vssd1 vccd1 vccd1 _13323_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17090_ _17089_/B _17089_/C _17089_/A vssd1 vssd1 vccd1 vccd1 _17091_/C sky130_fd_sc_hd__o21bai_1
XFILLER_0_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16041_ _16424_/A _16377_/A _16042_/C _16213_/A vssd1 vssd1 vccd1 vccd1 _16043_/A
+ sky130_fd_sc_hd__a22o_1
X_13253_ _14138_/A _13858_/C _13402_/D _14463_/D vssd1 vssd1 vccd1 vccd1 _13253_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12204_ _12203_/A _12202_/Y _12160_/X _12177_/Y vssd1 vssd1 vccd1 vccd1 _12207_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_62_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13184_ _13184_/A _13184_/B vssd1 vssd1 vccd1 vccd1 _13193_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_270 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19800_ _19719_/A _19719_/C _19719_/B vssd1 vssd1 vccd1 vccd1 _19841_/A sky130_fd_sc_hd__a21bo_1
X_12135_ _12091_/A _12091_/C _12091_/B vssd1 vssd1 vccd1 vccd1 _12141_/B sky130_fd_sc_hd__a21o_1
X_17992_ _18849_/B _18732_/C _19221_/C _19185_/D vssd1 vssd1 vccd1 vccd1 _17993_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16943_ _16943_/A _16943_/B vssd1 vssd1 vccd1 vccd1 _16946_/B sky130_fd_sc_hd__xnor2_2
X_19731_ _19732_/B _20249_/B _21171_/B _19732_/A vssd1 vssd1 vccd1 vccd1 _19734_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15308__B _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12066_ _12066_/A _12066_/B _12066_/C vssd1 vssd1 vccd1 vccd1 _12066_/X sky130_fd_sc_hd__or3_1
XANTENNA__12857__A1 _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12857__B2 _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14212__B _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11328__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11017_ mstream_o[91] hold56/X _11027_/S vssd1 vssd1 vccd1 vccd1 _21628_/D sky130_fd_sc_hd__mux2_1
X_16874_ _16873_/B _16873_/C _16873_/A vssd1 vssd1 vccd1 vccd1 _16876_/B sky130_fd_sc_hd__a21bo_1
X_19662_ _19531_/A _20671_/B _19528_/X _19529_/X _21278_/A vssd1 vssd1 vccd1 vccd1
+ _19667_/A sky130_fd_sc_hd__a32o_1
XANTENNA__14059__B1 _14217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15825_ _15650_/B _15689_/Y _15823_/X _15824_/Y vssd1 vssd1 vccd1 vccd1 _15874_/A
+ sky130_fd_sc_hd__o211a_1
X_18613_ _18454_/A _18454_/Y _18610_/Y _18611_/X vssd1 vssd1 vccd1 vccd1 _18613_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__18619__B _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19593_ _19291_/A _19291_/B _19589_/X _19590_/Y vssd1 vssd1 vccd1 vccd1 _19593_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__12609__A1 _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15756_ _15756_/A _15756_/B vssd1 vssd1 vccd1 vccd1 _16016_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_99_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18544_ _19008_/D _19013_/C _19179_/C _18857_/B vssd1 vssd1 vccd1 vccd1 _18544_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12968_ _12969_/A _12969_/B vssd1 vssd1 vccd1 vccd1 _13112_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21344__A2 _17595_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14707_ _14707_/A _14707_/B _14707_/C vssd1 vssd1 vccd1 vccd1 _14709_/A sky130_fd_sc_hd__and3_2
XANTENNA__19009__A1_N _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18475_ _18475_/A _18475_/B vssd1 vssd1 vccd1 vccd1 _18478_/C sky130_fd_sc_hd__xor2_1
X_11919_ _12781_/D _12619_/A vssd1 vssd1 vccd1 vccd1 _11923_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15687_ _15687_/A _15687_/B _15687_/C vssd1 vssd1 vccd1 vccd1 _15689_/B sky130_fd_sc_hd__nor3_2
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12899_ _14195_/A _12899_/B _13032_/A _12899_/D vssd1 vssd1 vccd1 vccd1 _13032_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17426_ _17427_/A _17427_/B _17427_/C vssd1 vssd1 vccd1 vccd1 _17426_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14638_ _14638_/A _14638_/B _14785_/B vssd1 vssd1 vccd1 vccd1 _14640_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15978__B _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17357_ _17356_/A _17356_/B _17356_/C _17356_/D vssd1 vssd1 vccd1 vccd1 _17357_/Y
+ sky130_fd_sc_hd__o22ai_1
X_14569_ _14418_/A _14418_/B _14567_/X _14568_/Y vssd1 vssd1 vccd1 vccd1 _14571_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19170__B1 _14296_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16308_ _16308_/A _16308_/B vssd1 vssd1 vccd1 vccd1 _16310_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17288_ _17288_/A _17288_/B vssd1 vssd1 vccd1 vccd1 _17290_/B sky130_fd_sc_hd__xor2_1
XANTENNA__21211__D _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19027_ _18905_/A _18904_/B _18902_/X vssd1 vssd1 vccd1 vccd1 _19037_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_71_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16239_ _16235_/A _16237_/Y _16119_/B _16120_/Y vssd1 vssd1 vccd1 vccd1 _16240_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__14534__A1 _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20108__C _20249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16305__D _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11348__A1 _11347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18801__C _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19185__B _19185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16602__B _17666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19225__A1 _19379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19929_ _19929_/A _19929_/B vssd1 vssd1 vccd1 vccd1 _19932_/A sky130_fd_sc_hd__xor2_1
XANTENNA__16039__A1 _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16039__B2 _16391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout199_A _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11520__A1 _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11520__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16975__D _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17433__B _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20791__B1 _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12858__A _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout366_A _14663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19351__D _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15234__A _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19528__A2 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21822_ _21822_/CLK _21822_/D vssd1 vssd1 vccd1 vccd1 _21822_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__13680__C _14477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21335__A2 _12392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11284__A0 _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21753_ _22049_/CLK _21753_/D vssd1 vssd1 vccd1 vccd1 _21753_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_fanout533_A _21737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20794__B _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18545__A _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20704_ _20700_/A _20701_/Y _20530_/Y _20532_/Y vssd1 vssd1 vccd1 vccd1 _20705_/B
+ sky130_fd_sc_hd__o211ai_1
X_21684_ _22069_/CLK _21684_/D vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20635_ _20632_/Y _20633_/X _20501_/Y _20503_/Y vssd1 vssd1 vccd1 vccd1 _20635_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20566_ _20567_/B _20567_/A vssd1 vssd1 vccd1 vccd1 _20698_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_104_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17711__B2 _11547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16215__D _16418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20497_ _20498_/A _20498_/B _20498_/C vssd1 vssd1 vccd1 vccd1 _20499_/C sky130_fd_sc_hd__o21a_2
XFILLER_0_14_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11339__A1 _21407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18711__C _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17608__B _18851_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16512__B _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_886 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21118_ _20955_/X _20958_/Y _21188_/B _21117_/X vssd1 vssd1 vccd1 vccd1 _21236_/A
+ sky130_fd_sc_hd__a211oi_2
X_22098_ _22105_/CLK _22098_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[34] sky130_fd_sc_hd__dfrtp_4
XANTENNA__19823__B _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout240 _21808_/Q vssd1 vssd1 vccd1 vccd1 _17915_/D sky130_fd_sc_hd__buf_4
Xfanout251 _17334_/B vssd1 vssd1 vccd1 vccd1 _20583_/A sky130_fd_sc_hd__buf_6
Xfanout262 _21803_/Q vssd1 vssd1 vccd1 vccd1 _19823_/A sky130_fd_sc_hd__buf_4
XFILLER_0_121_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13940_ _13939_/B _13939_/C _13939_/A vssd1 vssd1 vccd1 vccd1 _13940_/Y sky130_fd_sc_hd__a21oi_1
X_21049_ _21050_/A _21050_/B vssd1 vssd1 vccd1 vccd1 _21207_/A sky130_fd_sc_hd__nand2b_1
Xfanout273 _21800_/Q vssd1 vssd1 vccd1 vccd1 _17223_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_156_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11511__A1 _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout284 _21798_/Q vssd1 vssd1 vccd1 vccd1 _17520_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_89_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout295 _21796_/Q vssd1 vssd1 vccd1 vccd1 _17619_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_92_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11511__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13871_ _13871_/A _13871_/B vssd1 vssd1 vccd1 vccd1 _13884_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_97_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15610_ _15469_/B _15469_/Y _15608_/Y _15609_/X vssd1 vssd1 vccd1 vccd1 _15612_/C
+ sky130_fd_sc_hd__o211a_2
X_12822_ _12947_/B _12947_/C _12822_/C vssd1 vssd1 vccd1 vccd1 _12824_/A sky130_fd_sc_hd__and3_1
X_16590_ _16590_/A _16628_/A vssd1 vssd1 vccd1 vccd1 _16597_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_97_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_1011 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15541_ _15541_/A _15541_/B vssd1 vssd1 vccd1 vccd1 _15543_/B sky130_fd_sc_hd__or2_1
XFILLER_0_5_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11275__B1 _11274_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12753_ _13152_/C _12751_/X _12752_/X vssd1 vssd1 vccd1 vccd1 _12754_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_9_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17997__C _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18260_ _18261_/A _18261_/B vssd1 vssd1 vccd1 vccd1 _18260_/X sky130_fd_sc_hd__or2_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ _12297_/A _11702_/Y _11650_/A _11652_/B vssd1 vssd1 vccd1 vccd1 _11776_/B
+ sky130_fd_sc_hd__o211a_1
X_15472_ _15469_/Y _15470_/X _15287_/Y _15289_/Y vssd1 vssd1 vccd1 vccd1 _15473_/C
+ sky130_fd_sc_hd__o211ai_4
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ _12684_/A _12684_/B _12684_/C vssd1 vssd1 vccd1 vccd1 _12687_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_139_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17211_ _17211_/A _17211_/B vssd1 vssd1 vccd1 vccd1 _17213_/B sky130_fd_sc_hd__and2_1
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14423_ _14423_/A _14423_/B vssd1 vssd1 vccd1 vccd1 _14426_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_126_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18191_ _18332_/B _18192_/C vssd1 vssd1 vccd1 vccd1 _18193_/B sky130_fd_sc_hd__nor2_1
X_11635_ _11632_/X _11635_/B vssd1 vssd1 vccd1 vccd1 _11793_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_154_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11578__A1 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20837__A1 _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17142_ _17141_/A _17145_/B _17146_/C _17141_/B vssd1 vssd1 vccd1 vccd1 _17142_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14354_ _15695_/A _14508_/A _14354_/C _14817_/D vssd1 vssd1 vccd1 vccd1 _14357_/D
+ sky130_fd_sc_hd__nand4_1
XANTENNA__20837__B2 _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11566_ _11566_/A _11566_/B vssd1 vssd1 vccd1 vccd1 _11573_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_53_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13305_ _13306_/A _13306_/B _13306_/C vssd1 vssd1 vccd1 vccd1 _13343_/A sky130_fd_sc_hd__and3_2
XFILLER_0_80_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17073_ _17073_/A _17073_/B _17073_/C vssd1 vssd1 vccd1 vccd1 _17078_/A sky130_fd_sc_hd__and3_1
XFILLER_0_122_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14285_ _14121_/A _14285_/B vssd1 vssd1 vccd1 vccd1 _14289_/B sky130_fd_sc_hd__and2b_1
X_11497_ _11496_/X _19068_/C _11521_/S vssd1 vssd1 vccd1 vccd1 _21837_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_123_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16024_ fanout9/A _21409_/B vssd1 vssd1 vccd1 vccd1 _16024_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_122_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13236_ _13394_/A _16328_/B _13376_/A _13234_/Y vssd1 vssd1 vccd1 vccd1 _13237_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_27_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13167_ _13166_/B _13166_/C _13166_/A vssd1 vssd1 vccd1 vccd1 _13168_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_23_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12118_ _12118_/A _12118_/B vssd1 vssd1 vccd1 vccd1 _12120_/C sky130_fd_sc_hd__nor2_1
X_13098_ _13381_/C _14155_/C _14155_/D _13394_/A vssd1 vssd1 vccd1 vccd1 _13100_/A
+ sky130_fd_sc_hd__a22oi_1
X_17975_ _17975_/A _17975_/B vssd1 vssd1 vccd1 vccd1 _17989_/A sky130_fd_sc_hd__and2_1
XFILLER_0_137_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11058__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19714_ _19715_/A _19715_/B _19715_/C vssd1 vssd1 vccd1 vccd1 _19714_/X sky130_fd_sc_hd__and3_1
X_16926_ _16926_/A _16926_/B vssd1 vssd1 vccd1 vccd1 _16928_/A sky130_fd_sc_hd__nor2_1
X_12049_ _12043_/A _12043_/C _12043_/B vssd1 vssd1 vccd1 vccd1 _12050_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11502__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11502__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21056__A _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18349__B _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19645_ _19645_/A _19645_/B vssd1 vssd1 vccd1 vccd1 _19647_/A sky130_fd_sc_hd__nand2_1
X_16857_ _17165_/C _16855_/C _16855_/A vssd1 vssd1 vccd1 vccd1 _17168_/B sky130_fd_sc_hd__o21a_1
X_15808_ _15927_/A _16414_/B _15808_/C _15808_/D vssd1 vssd1 vccd1 vccd1 _15927_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_88_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13255__A1 _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16788_ _16718_/Y _16786_/X _16785_/X _16778_/X vssd1 vssd1 vccd1 vccd1 _16789_/C
+ sky130_fd_sc_hd__a211o_1
X_19576_ _19415_/Y _19417_/X _19573_/X _19575_/Y vssd1 vssd1 vccd1 vccd1 _19578_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_62_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21490__S _21490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12397__B _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15739_ _15737_/B _15737_/C _15737_/A vssd1 vssd1 vccd1 vccd1 _15741_/D sky130_fd_sc_hd__a21oi_2
XFILLER_0_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18527_ _18377_/C _18378_/X _18525_/Y _18526_/X vssd1 vssd1 vccd1 vccd1 _18529_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18458_ _18305_/A _18305_/Y _18456_/X _18457_/Y vssd1 vssd1 vccd1 vccd1 _18521_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14204__B1 _14203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13558__A2 _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17409_ _17409_/A _17487_/A _17409_/C vssd1 vssd1 vccd1 vccd1 _17487_/B sky130_fd_sc_hd__nor3_1
X_18389_ _18389_/A _18389_/B vssd1 vssd1 vccd1 vccd1 _18394_/C sky130_fd_sc_hd__xor2_4
XFILLER_0_69_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11521__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20420_ _20420_/A _20552_/B vssd1 vssd1 vccd1 vccd1 _20423_/A sky130_fd_sc_hd__or2_1
XFILLER_0_145_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20351_ _20352_/A _20352_/B vssd1 vssd1 vccd1 vccd1 _20351_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__15704__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout114_A _21839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20282_ _20282_/A _20282_/B vssd1 vssd1 vccd1 vccd1 _20290_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12860__B _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22021_ _22021_/CLK _22021_/D vssd1 vssd1 vccd1 vccd1 hold149/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_140_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_1104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15229__A _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout483_A _21748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18957__B1 _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21805_ _22021_/CLK _21805_/D vssd1 vssd1 vccd1 vccd1 hold330/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21736_ _21803_/CLK _21736_/D vssd1 vssd1 vccd1 vccd1 _21736_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16735__A2 _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout27_A _11348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16507__B _16734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21667_ _21906_/CLK _21667_/D vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14308__A _14463_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11431__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12757__B1 _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11420_ _11447_/A1 hold297/A fanout49/X hold116/A vssd1 vssd1 vccd1 vccd1 _11420_/X
+ sky130_fd_sc_hd__a22o_1
X_20618_ _20614_/Y _20616_/X _20480_/Y _20484_/A vssd1 vssd1 vccd1 vccd1 _20618_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_149_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15130__C _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19685__A1 _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21598_ _21888_/CLK _21598_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[61] sky130_fd_sc_hd__dfrtp_4
XANTENNA__19685__B2 _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17619__A _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11351_ fanout58/X v0z[31] fanout17/X _11350_/X vssd1 vssd1 vccd1 vccd1 _11351_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20549_ _21256_/A _20924_/A _20550_/C _20550_/D vssd1 vssd1 vccd1 vccd1 _20551_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_104_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14070_ _14070_/A _14070_/B _14070_/C vssd1 vssd1 vccd1 vccd1 _14072_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_104_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13866__B _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11282_ _11502_/A1 t1x[14] v2z[14] _11501_/B2 _11281_/X vssd1 vssd1 vccd1 vccd1 _11282_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__17338__B _17557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13182__B1 _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13021_ _13020_/B _13020_/C _13020_/A vssd1 vssd1 vccd1 vccd1 _13023_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13721__A2 _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14972_ _15085_/A vssd1 vssd1 vccd1 vccd1 _15501_/A sky130_fd_sc_hd__inv_2
X_17760_ _18767_/B _17758_/X _17759_/X vssd1 vssd1 vccd1 vccd1 _17761_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__18948__B1 _19751_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13923_ _14848_/A _14234_/C _13920_/Y _13921_/X vssd1 vssd1 vccd1 vccd1 _13924_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16711_ _16715_/B _16712_/B _16712_/C _16712_/D vssd1 vssd1 vccd1 vccd1 _16711_/X
+ sky130_fd_sc_hd__and4_1
X_17691_ _17575_/C _17574_/Y _17689_/X _17690_/Y vssd1 vssd1 vccd1 vccd1 _17693_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_117_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17504__D _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17620__B1 _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16642_ _16642_/A _16642_/B _16642_/C vssd1 vssd1 vccd1 vccd1 _16645_/A sky130_fd_sc_hd__nand3_1
X_19430_ _19430_/A _19951_/B _20242_/C _20242_/D vssd1 vssd1 vccd1 vccd1 _19598_/A
+ sky130_fd_sc_hd__nand4_2
X_13854_ _13973_/B _13852_/X _13736_/Y _13739_/Y vssd1 vssd1 vccd1 vccd1 _13854_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_57_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16974__A2 _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11248__A0 _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_97_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12805_ _12692_/C _12691_/Y _12803_/X _12804_/Y vssd1 vssd1 vccd1 vccd1 _12807_/C
+ sky130_fd_sc_hd__o211ai_4
X_16573_ _17520_/B _17874_/A _17041_/A _16899_/B vssd1 vssd1 vccd1 vccd1 _17211_/A
+ sky130_fd_sc_hd__nand4_1
X_19361_ _19519_/A _19359_/Y _19204_/B _19206_/B vssd1 vssd1 vccd1 vccd1 _19362_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13785_ _13784_/B _13784_/C _13784_/A vssd1 vssd1 vccd1 vccd1 _13787_/B sky130_fd_sc_hd__a21o_1
X_10997_ mstream_o[71] hold66/X _11005_/S vssd1 vssd1 vccd1 vccd1 _21608_/D sky130_fd_sc_hd__mux2_1
X_15524_ _16036_/A _15525_/B vssd1 vssd1 vccd1 vccd1 _15526_/A sky130_fd_sc_hd__and2_1
XFILLER_0_96_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18312_ _19686_/A _18929_/B _18616_/D _19686_/B vssd1 vssd1 vccd1 vccd1 _18314_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12736_ _13556_/A _13573_/D _12856_/A _12734_/Y vssd1 vssd1 vccd1 vccd1 _12736_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_29_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18616__C _18929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19292_ _19292_/A _19292_/B vssd1 vssd1 vccd1 vccd1 _19295_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__17520__C _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16726__A2 _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11263__A3 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18243_ _18243_/A _18243_/B vssd1 vssd1 vccd1 vccd1 _18394_/B sky130_fd_sc_hd__or2_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19810__A_N _19650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15455_ _15961_/D _15978_/B _15453_/Y _15587_/A vssd1 vssd1 vccd1 vccd1 _15457_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_26_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18335__D _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12667_ _12667_/A _12667_/B vssd1 vssd1 vccd1 vccd1 _12687_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_127_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14218__A _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14406_ _14557_/A _14557_/B _15001_/B _15510_/B vssd1 vssd1 vccd1 vccd1 _14554_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_26_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18174_ _18322_/B _18174_/B vssd1 vssd1 vccd1 vccd1 _18177_/A sky130_fd_sc_hd__nor2_1
X_11618_ _11588_/A _11591_/A _11615_/X _11617_/Y vssd1 vssd1 vccd1 vccd1 _11667_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_154_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15386_ _15386_/A _15386_/B _15386_/C vssd1 vssd1 vccd1 vccd1 _15386_/X sky130_fd_sc_hd__and3_1
XFILLER_0_128_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12598_ _12825_/B _12598_/B vssd1 vssd1 vccd1 vccd1 _12957_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17125_ _17146_/A _17123_/C _17141_/C _17146_/B vssd1 vssd1 vccd1 vccd1 _17126_/D
+ sky130_fd_sc_hd__a22o_1
X_14337_ _14489_/B _14337_/B vssd1 vssd1 vccd1 vccd1 _14340_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_107_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11420__B1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11549_ _11549_/A hold2/A vssd1 vssd1 vccd1 vccd1 _11550_/B sky130_fd_sc_hd__or2_4
XFILLER_0_52_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17056_ _17096_/A _17146_/C _17054_/B _17052_/X vssd1 vssd1 vccd1 vccd1 _17074_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13776__B _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14268_ _14268_/A _14268_/B _14268_/C vssd1 vssd1 vccd1 vccd1 _14268_/X sky130_fd_sc_hd__and3_1
XFILLER_0_111_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19428__B2 _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16007_ _16007_/A _16007_/B vssd1 vssd1 vccd1 vccd1 _16010_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13219_ _13218_/B _13218_/C _13218_/A vssd1 vssd1 vccd1 vccd1 _13219_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11577__A _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14199_ _14198_/B _14198_/C _14198_/A vssd1 vssd1 vccd1 vccd1 _14201_/B sky130_fd_sc_hd__a21o_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17958_ _17958_/A _17958_/B _17958_/C vssd1 vssd1 vccd1 vccd1 _17958_/X sky130_fd_sc_hd__and3_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14673__B1 _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18403__A2 _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16909_ _16909_/A _16916_/A vssd1 vssd1 vccd1 vccd1 _17167_/B sky130_fd_sc_hd__nand2_1
XANTENNA__19600__A1 _19732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17889_ _17975_/A _17887_/Y _17747_/Y _17750_/X vssd1 vssd1 vccd1 vccd1 _17890_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__19600__B2 _19732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12839__C _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19628_ _19629_/A _19629_/B vssd1 vssd1 vccd1 vccd1 _19628_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11239__B1 _11238_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19559_ _19556_/X _19557_/Y _19424_/B _19426_/A vssd1 vssd1 vccd1 vccd1 _19560_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_87_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17914__B2 _17670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15231__B _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14728__A1 _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21521_ hold239/X sstream_i[98] _21528_/S vssd1 vssd1 vccd1 vccd1 _22048_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout231_A _17670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19116__B1 _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout329_A _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21452_ hold175/X sstream_i[29] _21507_/S vssd1 vssd1 vccd1 vccd1 _21979_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15154__A1_N _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20403_ _20403_/A _20403_/B vssd1 vssd1 vccd1 vccd1 _20404_/B sky130_fd_sc_hd__xor2_1
X_21383_ _21381_/B _21382_/X _21381_/Y vssd1 vssd1 vccd1 vccd1 _21935_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17142__A2 _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20334_ _20845_/D _21311_/B _20332_/Y _20472_/A vssd1 vssd1 vccd1 vccd1 _20336_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_141_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16062__B _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20265_ _20863_/C _21291_/A _21278_/A _20265_/D vssd1 vssd1 vccd1 vccd1 _20473_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_101_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22004_ _22005_/CLK _22004_/D vssd1 vssd1 vccd1 vccd1 hold116/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19373__B _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20196_ _20196_/A _20196_/B vssd1 vssd1 vccd1 vccd1 _20198_/B sky130_fd_sc_hd__xor2_1
XANTENNA__17324__D _17324_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10920_ mstream_o[52] _10919_/X _10992_/S vssd1 vssd1 vccd1 vccd1 _21589_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_67_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10851_ _10802_/X _10859_/A _10805_/Y _11066_/A vssd1 vssd1 vccd1 vccd1 _10852_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ _14024_/B _14516_/A _14365_/C _14027_/A vssd1 vssd1 vccd1 vccd1 _13570_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_52_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ _12521_/A _12521_/B _12521_/C vssd1 vssd1 vccd1 vccd1 _12522_/C sky130_fd_sc_hd__and3_1
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21719_ _21974_/CLK hold1/X _21422_/A vssd1 vssd1 vccd1 vccd1 _21719_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15240_ _15240_/A _15240_/B vssd1 vssd1 vccd1 vccd1 _15242_/B sky130_fd_sc_hd__xnor2_2
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12452_ _13157_/A _12781_/D vssd1 vssd1 vccd1 vccd1 _12456_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11403_ hold285/A fanout28/X _11402_/X vssd1 vssd1 vccd1 vccd1 _11403_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_152_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15171_ _15961_/D _15717_/C _15976_/D _15838_/D vssd1 vssd1 vccd1 vccd1 _15171_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__13877__A _13877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12383_ _11669_/X _11671_/Y _12381_/Y _12382_/X vssd1 vssd1 vccd1 vccd1 _12383_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_22_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14122_ _14121_/A _14121_/B _13834_/A vssd1 vssd1 vccd1 vccd1 _14123_/C sky130_fd_sc_hd__o21bai_2
XANTENNA__18171__C _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11334_ _11544_/A1 t1x[27] v2z[27] _11543_/B2 _11333_/X vssd1 vssd1 vccd1 vccd1 _11334_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_120_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14053_ _14212_/B _14365_/D vssd1 vssd1 vccd1 vccd1 _14057_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18930_ _18773_/B _18929_/X _18928_/X vssd1 vssd1 vccd1 vccd1 _18931_/B sky130_fd_sc_hd__a21bo_1
X_11265_ _11325_/A1 t2y[10] t0y[10] _11498_/A1 vssd1 vssd1 vccd1 vccd1 _11265_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_123_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13004_ _13002_/B _13002_/C _13002_/A vssd1 vssd1 vccd1 vccd1 _13004_/Y sky130_fd_sc_hd__a21oi_1
X_18861_ _18861_/A vssd1 vssd1 vccd1 vccd1 _18863_/B sky130_fd_sc_hd__inv_2
XANTENNA__20976__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11196_ hold291/X fanout51/X fanout48/X hold233/X vssd1 vssd1 vccd1 vccd1 _11196_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12005__B _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17812_ _17689_/C _17688_/Y _17810_/X _17811_/Y vssd1 vssd1 vccd1 vccd1 _17812_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14501__A _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18792_ _18790_/X _18792_/B vssd1 vssd1 vccd1 vccd1 _18793_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_118_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14955_ _14954_/B _14954_/C _14954_/A vssd1 vssd1 vccd1 vccd1 _14956_/C sky130_fd_sc_hd__a21o_1
X_17743_ _17743_/A _17870_/B _17743_/C vssd1 vssd1 vccd1 vccd1 _17743_/X sky130_fd_sc_hd__and3_1
XANTENNA__21037__C _21283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18397__A1 _17841_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11336__S _11348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17234__D _17443_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13906_ _13906_/A _14051_/B _13906_/C vssd1 vssd1 vccd1 vccd1 _13906_/X sky130_fd_sc_hd__and3_2
X_14886_ _14883_/X _14884_/Y _14705_/B _14707_/B vssd1 vssd1 vccd1 vccd1 _14887_/D
+ sky130_fd_sc_hd__o211a_1
X_17674_ _17673_/B _17673_/C _17673_/A vssd1 vssd1 vccd1 vccd1 _17676_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19413_ _20394_/B _19414_/C _19866_/D _19972_/A vssd1 vssd1 vccd1 vccd1 _19417_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21334__A _21407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13837_ _14306_/A _14138_/A _14477_/C _14155_/D vssd1 vssd1 vccd1 vccd1 _13839_/D
+ sky130_fd_sc_hd__nand4_1
X_16625_ _16625_/A _16625_/B _16625_/C vssd1 vssd1 vccd1 vccd1 _16629_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_43_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13572__A1_N _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11860__A _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16556_ _21825_/Q _17433_/A _17526_/B _16734_/B vssd1 vssd1 vccd1 vccd1 _16557_/B
+ sky130_fd_sc_hd__a22o_1
X_19344_ _19345_/A _19345_/B vssd1 vssd1 vccd1 vccd1 _19346_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_57_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13768_ _13767_/B _13910_/B _13767_/A vssd1 vssd1 vccd1 vccd1 _13769_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_73_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15507_ _15632_/B _16369_/B _16177_/B _15892_/A vssd1 vssd1 vccd1 vccd1 _15510_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12719_ _12719_/A vssd1 vssd1 vccd1 vccd1 _12721_/A sky130_fd_sc_hd__inv_2
X_16487_ _17300_/C _17520_/D _17282_/A _17277_/A vssd1 vssd1 vccd1 vccd1 _16495_/A
+ sky130_fd_sc_hd__and4_1
X_19275_ _19275_/A _19275_/B vssd1 vssd1 vccd1 vccd1 _19300_/A sky130_fd_sc_hd__and2_1
XFILLER_0_57_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13699_ _13698_/B _13698_/C _13698_/A vssd1 vssd1 vccd1 vccd1 _13699_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_116_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15438_ _15438_/A _15438_/B vssd1 vssd1 vccd1 vccd1 _15443_/A sky130_fd_sc_hd__xnor2_2
X_18226_ _18225_/B _18225_/C _18225_/A vssd1 vssd1 vccd1 vccd1 _18226_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_127_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15369_ _16027_/A _15370_/B _15370_/C _15548_/A vssd1 vssd1 vccd1 vccd1 _15371_/A
+ sky130_fd_sc_hd__a22o_1
X_18157_ _18157_/A _18157_/B _18143_/Y vssd1 vssd1 vccd1 vccd1 _18157_/Y sky130_fd_sc_hd__nor3b_4
XFILLER_0_26_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16163__A _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold304 hold304/A vssd1 vssd1 vccd1 vccd1 hold304/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17108_ _17106_/A _17120_/A _17078_/X _17083_/Y vssd1 vssd1 vccd1 vccd1 _17110_/B
+ sky130_fd_sc_hd__o211ai_1
Xhold315 hold315/A vssd1 vssd1 vccd1 vccd1 hold315/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18088_ _18107_/B _18087_/B _18087_/C _18087_/D vssd1 vssd1 vccd1 vccd1 _18088_/Y
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__18872__A2 _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold326 hold326/A vssd1 vssd1 vccd1 vccd1 hold326/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17039_ _17028_/Y _17038_/X _16994_/Y _17010_/X vssd1 vssd1 vccd1 vccd1 _17046_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_7_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11738__C _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20050_ _20049_/B _20188_/B _20049_/A vssd1 vssd1 vccd1 vccd1 _20051_/C sky130_fd_sc_hd__o21ai_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19821__A1 _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19821__B2 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20413__A _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16610__B _21823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14768__D _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout279_A _21799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20952_ _20952_/A _20952_/B _20952_/C vssd1 vssd1 vccd1 vccd1 _20953_/A sky130_fd_sc_hd__and3_1
XFILLER_0_36_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20883_ _20883_/A _20883_/B vssd1 vssd1 vccd1 vccd1 _20885_/B sky130_fd_sc_hd__xor2_1
XANTENNA__15071__B1 _10919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout446_A _21759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18256__C _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13621__A1 _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11227__A3 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12424__A2 _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13621__B2 _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21504_ hold311/X sstream_i[81] _21507_/S vssd1 vssd1 vccd1 vccd1 _22031_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21435_ hold250/X sstream_i[12] _21442_/S vssd1 vssd1 vccd1 vccd1 _21962_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18312__A1 _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18312__B2 _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21366_ hold94/X fanout40/X _21365_/X vssd1 vssd1 vccd1 vccd1 _21929_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20026__C _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20670__A2 _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20317_ _20178_/D _21293_/B _20721_/C _20317_/D vssd1 vssd1 vccd1 vccd1 _20321_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_101_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21297_ _21297_/A _21297_/B vssd1 vssd1 vccd1 vccd1 _21298_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout94_A fanout96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14024__C _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11050_ _11050_/A _11050_/B vssd1 vssd1 vccd1 vccd1 _11051_/B sky130_fd_sc_hd__nor2_2
XANTENNA__18615__A2 _18929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20248_ _20248_/A _20248_/B vssd1 vssd1 vccd1 vccd1 _20250_/A sky130_fd_sc_hd__nor2_1
XANTENNA__19812__B2 _19650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19534__D _19691_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20179_ _19644_/A _20178_/B _21261_/B _20032_/D vssd1 vssd1 vccd1 vccd1 _20180_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13863__C _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11156__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14740_ _14580_/A _14580_/B _14578_/X vssd1 vssd1 vccd1 vccd1 _14742_/B sky130_fd_sc_hd__a21oi_4
XTAP_3744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11952_ _12426_/B _12312_/A _11952_/C _11952_/D vssd1 vssd1 vccd1 vccd1 _12019_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_59_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10903_ _10911_/B _10903_/B vssd1 vssd1 vccd1 vccd1 _10903_/Y sky130_fd_sc_hd__nor2_2
XTAP_3788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14671_ _14671_/A _14671_/B vssd1 vssd1 vccd1 vccd1 _14679_/A sky130_fd_sc_hd__nand2_1
XTAP_3799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11883_ _11883_/A vssd1 vssd1 vccd1 vccd1 _11885_/A sky130_fd_sc_hd__inv_2
XFILLER_0_129_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16410_ _16410_/A _16410_/B vssd1 vssd1 vccd1 vccd1 _16411_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11680__A _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13622_ _13620_/X _13622_/B vssd1 vssd1 vccd1 vccd1 _13623_/B sky130_fd_sc_hd__and2b_1
XANTENNA__18166__C _18929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10834_ _11053_/A _11053_/B _10821_/A vssd1 vssd1 vccd1 vccd1 _11055_/A sky130_fd_sc_hd__o21a_2
X_17390_ _17488_/A _17488_/B vssd1 vssd1 vccd1 vccd1 _17391_/B sky130_fd_sc_hd__and2_1
XANTENNA__13612__A1 _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16341_ _16341_/A _16341_/B vssd1 vssd1 vccd1 vccd1 _16343_/B sky130_fd_sc_hd__xnor2_2
X_13553_ _13860_/A _13858_/C _13402_/D _13554_/B vssd1 vssd1 vccd1 vccd1 _13556_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_81_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19060_ _19373_/B _19060_/B _19060_/C _19060_/D vssd1 vssd1 vccd1 vccd1 _19060_/Y
+ sky130_fd_sc_hd__nand4_1
X_12504_ _13394_/A _14018_/C vssd1 vssd1 vccd1 vccd1 _12505_/B sky130_fd_sc_hd__nand2_1
X_16272_ _16177_/B _16271_/X _16270_/X vssd1 vssd1 vccd1 vccd1 _16274_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_152_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13484_ _13483_/A _13483_/B _13483_/C vssd1 vssd1 vccd1 vccd1 _13486_/C sky130_fd_sc_hd__a21o_1
X_15223_ _15501_/A _15223_/B vssd1 vssd1 vccd1 vccd1 _15225_/B sky130_fd_sc_hd__nand2_1
X_18011_ _18010_/A _20148_/C _18144_/A _18010_/D vssd1 vssd1 vccd1 vccd1 _18012_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12435_ _12435_/A _12435_/B vssd1 vssd1 vccd1 vccd1 _12437_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15154_ _15155_/C _15698_/B _15152_/Y _15305_/A vssd1 vssd1 vccd1 vccd1 _15154_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_12366_ _11736_/A _11736_/C _11736_/B vssd1 vssd1 vccd1 vccd1 _12367_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_23_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14105_ _14105_/A _14105_/B _14105_/C vssd1 vssd1 vccd1 vccd1 _14105_/Y sky130_fd_sc_hd__nor3_2
X_11317_ _11325_/A1 t2y[23] t0y[23] _21723_/D vssd1 vssd1 vccd1 vccd1 _11317_/X sky130_fd_sc_hd__a22o_1
X_15085_ _15085_/A _15502_/A _15085_/C _15085_/D vssd1 vssd1 vccd1 vccd1 _15223_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_10_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19962_ _19847_/X _19857_/Y _19858_/X _19961_/A vssd1 vssd1 vccd1 vccd1 _19963_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13679__A1 _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12297_ _12297_/A _12297_/B vssd1 vssd1 vccd1 vccd1 _12315_/A sky130_fd_sc_hd__nor2_1
X_14036_ _21741_/Q _14365_/C _14037_/C _14190_/A vssd1 vssd1 vccd1 vccd1 _14038_/B
+ sky130_fd_sc_hd__a22o_1
X_18913_ _18912_/B _19065_/B _18912_/A vssd1 vssd1 vccd1 vccd1 _18914_/C sky130_fd_sc_hd__a21o_1
X_11248_ _12223_/A _11247_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21763_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17526__B _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19893_ _19893_/A _19893_/B vssd1 vssd1 vccd1 vccd1 _19902_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18844_ hold115/X _18843_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _21899_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13773__C _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11179_ hold184/X fanout22/X _11178_/X vssd1 vssd1 vccd1 vccd1 _11179_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_101_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1025 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18775_ _18775_/A _18775_/B _18775_/C vssd1 vssd1 vccd1 vccd1 _18775_/X sky130_fd_sc_hd__and3_1
X_15987_ _15856_/Y _15860_/A _15984_/Y _15986_/X vssd1 vssd1 vccd1 vccd1 _15987_/X
+ sky130_fd_sc_hd__a211o_2
XANTENNA__12103__A1 _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15761__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18638__A _19732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17726_ _21795_/Q _19337_/D _19692_/C _19691_/D vssd1 vssd1 vccd1 vccd1 _17865_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__17542__A _21803_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14938_ _21733_/Q _15838_/B _16374_/B _14774_/D vssd1 vssd1 vccd1 vccd1 _14939_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__19031__A2 _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17899__D _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17657_ _17657_/A _20583_/A _19951_/A _19951_/B vssd1 vssd1 vccd1 vccd1 _17777_/A
+ sky130_fd_sc_hd__nand4_2
X_14869_ _14732_/A _14732_/C _14732_/B vssd1 vssd1 vccd1 vccd1 _14883_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16608_ _16608_/A _16608_/B _16608_/C vssd1 vssd1 vccd1 vccd1 _16615_/A sky130_fd_sc_hd__nand3_1
X_17588_ _17589_/A _17589_/B vssd1 vssd1 vccd1 vccd1 _17830_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19327_ _19327_/A _19327_/B vssd1 vssd1 vccd1 vccd1 _19465_/A sky130_fd_sc_hd__or2_1
XFILLER_0_46_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16539_ _17636_/B _17282_/A _16531_/B _16530_/B vssd1 vssd1 vccd1 vccd1 _16547_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19258_ _19258_/A _19258_/B vssd1 vssd1 vccd1 vccd1 _19260_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16605__B _17334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18209_ _18209_/A _18209_/B _18209_/C vssd1 vssd1 vccd1 vccd1 _18212_/A sky130_fd_sc_hd__nand3_2
X_19189_ _19189_/A _19189_/B vssd1 vssd1 vccd1 vccd1 _19190_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__14406__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16204__A2_N _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21220_ _21220_/A _21220_/B vssd1 vssd1 vccd1 vccd1 _21222_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold101 hold101/A vssd1 vssd1 vccd1 vccd1 hold101/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 hold112/A vssd1 vssd1 vccd1 vccd1 hold112/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold123 hold123/A vssd1 vssd1 vccd1 vccd1 hold123/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold134 hold134/A vssd1 vssd1 vccd1 vccd1 hold134/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold145 hold145/A vssd1 vssd1 vccd1 vccd1 hold145/X sky130_fd_sc_hd__dlygate4sd3_1
X_21151_ _21151_/A _21301_/A _21815_/Q vssd1 vssd1 vccd1 vccd1 _21151_/X sky130_fd_sc_hd__and3_1
Xhold156 hold156/A vssd1 vssd1 vccd1 vccd1 hold156/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 hold167/A vssd1 vssd1 vccd1 vccd1 hold167/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold178 hold178/A vssd1 vssd1 vccd1 vccd1 hold178/X sky130_fd_sc_hd__dlygate4sd3_1
X_20102_ _20103_/A _21815_/Q _20103_/C _20282_/A vssd1 vssd1 vccd1 vccd1 _20104_/A
+ sky130_fd_sc_hd__a22o_1
Xhold189 hold189/A vssd1 vssd1 vccd1 vccd1 hold189/X sky130_fd_sc_hd__dlygate4sd3_1
X_21082_ _21199_/A _21291_/B _21083_/C _21083_/D vssd1 vssd1 vccd1 vccd1 _21084_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_10_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout603 _11459_/B2 vssd1 vssd1 vccd1 vccd1 _11507_/B2 sky130_fd_sc_hd__buf_2
Xfanout614 _21568_/S vssd1 vssd1 vccd1 vccd1 _21579_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout625 _21822_/Q vssd1 vssd1 vccd1 vccd1 _17557_/A sky130_fd_sc_hd__buf_4
XANTENNA_fanout396_A _21770_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11145__A2 _11122_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout636 _11089_/A vssd1 vssd1 vccd1 vccd1 fanout636/X sky130_fd_sc_hd__clkbuf_8
X_20033_ _20035_/A vssd1 vssd1 vccd1 vccd1 _20185_/A sky130_fd_sc_hd__inv_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout563_A _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20797__B _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15831__A2 _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21365__B1 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21984_ _22016_/CLK _21984_/D vssd1 vssd1 vccd1 vccd1 hold209/A sky130_fd_sc_hd__dfxtp_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20935_ _20936_/A _20936_/B vssd1 vssd1 vccd1 vccd1 _21110_/B sky130_fd_sc_hd__or2_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20866_ _20866_/A _20866_/B vssd1 vssd1 vccd1 vccd1 _20868_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold239_A hold239/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20797_ _20797_/A _21258_/A _21815_/Q _21046_/B vssd1 vssd1 vccd1 vccd1 _20931_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__18283__A _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13858__C _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12220_ _12267_/A _12246_/D _12269_/C _12242_/B vssd1 vssd1 vccd1 vccd1 _12222_/A
+ sky130_fd_sc_hd__a22oi_2
X_21418_ _16362_/Y _21248_/Y _21420_/S vssd1 vssd1 vccd1 vccd1 _21418_/X sky130_fd_sc_hd__mux2_1
XANTENNA__11659__B _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14035__B _21742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12151_ _12223_/A _12246_/D _12146_/A _12144_/B vssd1 vssd1 vccd1 vccd1 _12154_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_102_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21349_ _21349_/A _21349_/B vssd1 vssd1 vccd1 vccd1 _21349_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_124_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18049__B1 _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11102_ _10860_/Y hold152/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21696_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12082_ _12286_/C _12036_/X _12078_/Y _12080_/X vssd1 vssd1 vccd1 vccd1 _12082_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_60_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15910_ _16326_/A _15911_/C _16040_/C _15911_/A vssd1 vssd1 vccd1 vccd1 _15913_/C
+ sky130_fd_sc_hd__a22o_1
X_11033_ mstream_o[107] hold288/X _11039_/S vssd1 vssd1 vccd1 vccd1 hold289/A sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16890_ _16890_/A _16890_/B _16890_/C vssd1 vssd1 vccd1 vccd1 _16890_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_21_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17272__A1 _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15841_ _15841_/A _15971_/A _15841_/C vssd1 vssd1 vccd1 vccd1 _15966_/B sky130_fd_sc_hd__nor3_1
XANTENNA__17272__B2 _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18560_ _18561_/A _18561_/B vssd1 vssd1 vccd1 vccd1 _18560_/Y sky130_fd_sc_hd__nand2_1
X_15772_ _15772_/A _16029_/A vssd1 vssd1 vccd1 vccd1 _15773_/B sky130_fd_sc_hd__and2_1
XTAP_3530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12984_ _12984_/A _12984_/B vssd1 vssd1 vccd1 vccd1 _12986_/B sky130_fd_sc_hd__nor2_1
XTAP_3541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17511_ _17512_/A _17512_/B _17512_/C vssd1 vssd1 vccd1 vccd1 _17513_/B sky130_fd_sc_hd__a21o_2
X_14723_ _14723_/A _14723_/B vssd1 vssd1 vccd1 vccd1 _14735_/A sky130_fd_sc_hd__nor2_2
X_11935_ _11923_/A _11922_/A _11922_/B vssd1 vssd1 vccd1 vccd1 _11938_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__11844__B1 _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18491_ _18491_/A _18491_/B vssd1 vssd1 vccd1 vccd1 _18511_/A sky130_fd_sc_hd__xnor2_2
XTAP_3585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14654_ _14654_/A _14654_/B vssd1 vssd1 vccd1 vccd1 _14747_/A sky130_fd_sc_hd__xnor2_4
X_17442_ _20583_/A _18058_/A vssd1 vssd1 vccd1 vccd1 _17446_/A sky130_fd_sc_hd__nand2_1
XTAP_2884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11866_ _11867_/A _11867_/B vssd1 vssd1 vccd1 vccd1 _11889_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_156_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13605_ _13605_/A _13605_/B _13605_/C vssd1 vssd1 vccd1 vccd1 _13605_/X sky130_fd_sc_hd__or3_2
XFILLER_0_89_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10817_ hold227/A hold229/A vssd1 vssd1 vccd1 vccd1 _10817_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14585_ _14431_/A _14431_/B _14429_/X vssd1 vssd1 vccd1 vccd1 _14587_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_89_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17373_ _17381_/A _17381_/B _17380_/B vssd1 vssd1 vccd1 vccd1 _17374_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_39_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15032__D _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11797_ _11795_/A _11795_/Y _11796_/Y _11771_/X vssd1 vssd1 vccd1 vccd1 _11801_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_131_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19112_ _19112_/A _19112_/B _19276_/B vssd1 vssd1 vccd1 vccd1 _19112_/X sky130_fd_sc_hd__and3_1
X_16324_ _16324_/A _16324_/B vssd1 vssd1 vccd1 vccd1 _16331_/A sky130_fd_sc_hd__nor2_1
X_13536_ _13536_/A _13536_/B vssd1 vssd1 vccd1 vccd1 _13539_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20331__A1 _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21331__B _21331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20331__B2 _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12953__B _17834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16255_ _16143_/A _16143_/B _16142_/A _16141_/Y _16256_/A vssd1 vssd1 vccd1 vccd1
+ _16361_/B sky130_fd_sc_hd__o311a_1
X_19043_ _19174_/B _19043_/B _19176_/A _19043_/D vssd1 vssd1 vccd1 vccd1 _19176_/B
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_70_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13467_ _14848_/A _14391_/B vssd1 vssd1 vccd1 vccd1 _13471_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_153_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15206_ _15206_/A _15206_/B vssd1 vssd1 vccd1 vccd1 _15207_/A sky130_fd_sc_hd__and2_1
XANTENNA__13130__A _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12418_ _12479_/A vssd1 vssd1 vccd1 vccd1 _12418_/Y sky130_fd_sc_hd__inv_2
X_16186_ _16032_/A _16035_/A _16184_/X _16185_/Y vssd1 vssd1 vccd1 vccd1 _16303_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11569__B _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13398_ _13398_/A _13398_/B vssd1 vssd1 vccd1 vccd1 _13400_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18640__B _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15137_ _15037_/A _15037_/C _15037_/B vssd1 vssd1 vccd1 vccd1 _15138_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12349_ _12350_/A _12350_/B vssd1 vssd1 vccd1 vccd1 _12437_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_142_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15068_ _15068_/A _15068_/B vssd1 vssd1 vccd1 vccd1 _15206_/B sky130_fd_sc_hd__nor2_2
X_19945_ hold87/X fanout8/X vssd1 vssd1 vccd1 vccd1 _19945_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__16160__B _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14019_ _15155_/C _16414_/A _14020_/C _14020_/D vssd1 vssd1 vccd1 vccd1 _14021_/A
+ sky130_fd_sc_hd__a22o_1
X_19876_ _19873_/Y _19874_/X _19753_/D _19753_/Y vssd1 vssd1 vccd1 vccd1 _19877_/C
+ sky130_fd_sc_hd__o211ai_2
X_18827_ _18846_/B _18826_/B _18826_/C _18826_/D vssd1 vssd1 vccd1 vccd1 _18827_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18758_ _18758_/A _18758_/B _18758_/C vssd1 vssd1 vccd1 vccd1 _18758_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__21347__B1 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17709_ _17594_/A _17595_/A _17708_/X vssd1 vssd1 vccd1 vccd1 _17710_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_77_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18689_ _21142_/A _18689_/B vssd1 vssd1 vccd1 vccd1 _18689_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_78_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11524__S _11545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20720_ _20720_/A _20720_/B vssd1 vssd1 vccd1 vccd1 _20724_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_77_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13588__B1 _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19199__A _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20651_ _20651_/A _20651_/B vssd1 vssd1 vccd1 vccd1 _20662_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout144_A _21833_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15520__A _16031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18433__A1_N _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20582_ _20975_/D _21286_/B _21296_/B _20845_/D vssd1 vssd1 vccd1 vccd1 _20586_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout311_A _18851_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout409_A _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19646__B _20841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21203_ _21204_/A _21204_/B vssd1 vssd1 vccd1 vccd1 _21203_/X sky130_fd_sc_hd__and2_1
XFILLER_0_83_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13975__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16989__C _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17447__A _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21134_ _21134_/A _21134_/B vssd1 vssd1 vccd1 vccd1 _21137_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_100_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout400 _13157_/B vssd1 vssd1 vccd1 vccd1 _12426_/B sky130_fd_sc_hd__buf_4
Xfanout411 _14698_/A vssd1 vssd1 vccd1 vccd1 _15514_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__20592__A1_N _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout422 _12771_/C vssd1 vssd1 vccd1 vccd1 _12897_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout433 _14712_/B vssd1 vssd1 vccd1 vccd1 _14713_/B sky130_fd_sc_hd__buf_4
XFILLER_0_100_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21065_ _21065_/A _21065_/B vssd1 vssd1 vccd1 vccd1 _21067_/A sky130_fd_sc_hd__nand2_1
XANTENNA__20389__A1 _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout444 _12245_/B vssd1 vssd1 vccd1 vccd1 _12357_/C sky130_fd_sc_hd__buf_4
Xfanout455 _16380_/B vssd1 vssd1 vccd1 vccd1 _16286_/B sky130_fd_sc_hd__buf_4
Xfanout466 _14698_/D vssd1 vssd1 vccd1 vccd1 _15370_/B sky130_fd_sc_hd__clkbuf_8
Xfanout477 _21750_/Q vssd1 vssd1 vccd1 vccd1 _15093_/B sky130_fd_sc_hd__buf_4
X_20016_ _19879_/X _19885_/C _20125_/B _20015_/X vssd1 vssd1 vccd1 vccd1 _20168_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__19381__B _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout488 _21747_/Q vssd1 vssd1 vccd1 vccd1 _16328_/A sky130_fd_sc_hd__buf_4
Xfanout499 _21744_/Q vssd1 vssd1 vccd1 vccd1 _14365_/D sky130_fd_sc_hd__clkbuf_8
XANTENNA__15804__A2 _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21338__B1 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12618__A2 _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18203__B1 _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15414__B _15415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21967_ _21974_/CLK _21967_/D vssd1 vssd1 vccd1 vccd1 hold279/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13291__A2 _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11434__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _13018_/B _12780_/A _12780_/B _13017_/A vssd1 vssd1 vccd1 vccd1 _11722_/A
+ sky130_fd_sc_hd__a22oi_2
X_20918_ _20918_/A _20918_/B vssd1 vssd1 vccd1 vccd1 _20920_/A sky130_fd_sc_hd__xnor2_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21898_ _21948_/CLK hold23/X vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_84_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11651_ _11650_/A _11650_/B _11650_/C vssd1 vssd1 vccd1 vccd1 _11652_/C sky130_fd_sc_hd__a21o_1
X_20849_ _20849_/A _20849_/B vssd1 vssd1 vccd1 vccd1 _20852_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_83_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout40 _21390_/B vssd1 vssd1 vccd1 vccd1 fanout40/X sky130_fd_sc_hd__clkbuf_8
Xfanout51 _11122_/X vssd1 vssd1 vccd1 vccd1 fanout51/X sky130_fd_sc_hd__buf_4
XFILLER_0_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout62 _21853_/Q vssd1 vssd1 vccd1 vccd1 _20721_/C sky130_fd_sc_hd__buf_6
XFILLER_0_65_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14370_ _14370_/A _14370_/B _14370_/C vssd1 vssd1 vccd1 vccd1 _14373_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_107_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21151__B _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18444__C _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12251__B1 _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11582_ _12020_/A _14621_/D _12403_/A _12326_/D vssd1 vssd1 vccd1 vccd1 _11583_/B
+ sky130_fd_sc_hd__a22o_1
Xfanout73 _21849_/Q vssd1 vssd1 vccd1 vccd1 _20838_/C sky130_fd_sc_hd__buf_4
Xfanout84 _21846_/Q vssd1 vssd1 vccd1 vccd1 _20733_/C sky130_fd_sc_hd__buf_4
Xfanout95 fanout96/X vssd1 vssd1 vccd1 vccd1 _21278_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12773__B _21766_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13321_ _14712_/B _14391_/B _13913_/C _14712_/A vssd1 vssd1 vccd1 vccd1 _13322_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18741__A _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16040_ _16391_/A _16414_/A _16040_/C _16268_/B vssd1 vssd1 vccd1 vccd1 _16213_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ _13252_/A _13252_/B vssd1 vssd1 vccd1 vccd1 _13353_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_49_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ _12203_/A _12203_/B _12203_/C vssd1 vssd1 vccd1 vccd1 _12203_/X sky130_fd_sc_hd__or3_1
XFILLER_0_122_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16899__C _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13183_ _13183_/A _13183_/B vssd1 vssd1 vccd1 vccd1 _13184_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_0_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12134_ _12100_/A _12100_/C _12100_/B vssd1 vssd1 vccd1 vccd1 _12150_/B sky130_fd_sc_hd__a21o_1
XANTENNA__18690__B1 _21367_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17991_ _18849_/B _19185_/D _18732_/C _19221_/C vssd1 vssd1 vccd1 vccd1 _17991_/X
+ sky130_fd_sc_hd__and4_1
X_19730_ _19723_/A _21171_/B _19723_/C _19586_/X vssd1 vssd1 vccd1 vccd1 _19735_/A
+ sky130_fd_sc_hd__a31o_1
X_16942_ _16989_/C _17146_/C _16941_/B _16938_/X vssd1 vssd1 vccd1 vccd1 _16943_/B
+ sky130_fd_sc_hd__a31o_1
X_12065_ _12066_/A _12066_/B _12066_/C vssd1 vssd1 vccd1 vccd1 _12065_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__15308__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12857__A2 _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14212__C _14212_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11016_ mstream_o[90] hold3/X _11027_/S vssd1 vssd1 vccd1 vccd1 _21627_/D sky130_fd_sc_hd__mux2_1
XANTENNA__10868__A1 _10867_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19661_ _19661_/A _19661_/B vssd1 vssd1 vccd1 vccd1 _19669_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14059__A1 _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16873_ _16873_/A _16873_/B _16873_/C vssd1 vssd1 vccd1 vccd1 _16933_/A sky130_fd_sc_hd__nand3_1
XANTENNA__14059__B2 _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18188__A _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18612_ _18454_/A _18454_/Y _18610_/Y _18611_/X vssd1 vssd1 vccd1 vccd1 _18674_/A
+ sky130_fd_sc_hd__o211a_1
X_15824_ _15823_/B _15823_/C _15823_/A vssd1 vssd1 vccd1 vccd1 _15824_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__21329__B1 _21329_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19592_ _19291_/A _19291_/B _19589_/X _19590_/Y vssd1 vssd1 vccd1 vccd1 _19592_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12609__A2 _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18543_ _18543_/A _18543_/B vssd1 vssd1 vccd1 vccd1 _18576_/A sky130_fd_sc_hd__nor2_1
XTAP_3360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15755_ _15755_/A _15755_/B vssd1 vssd1 vccd1 vccd1 _15756_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_99_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12967_ _13250_/B _12967_/B vssd1 vssd1 vccd1 vccd1 _12969_/B sky130_fd_sc_hd__nor2_1
XTAP_3371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11344__S _11348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14706_ _14705_/B _14705_/C _14705_/A vssd1 vssd1 vccd1 vccd1 _14707_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11293__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11918_ _11917_/A _11917_/C _11917_/B vssd1 vssd1 vccd1 vccd1 _11924_/B sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_17_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18474_ _18475_/A _18475_/B vssd1 vssd1 vccd1 vccd1 _18474_/X sky130_fd_sc_hd__or2_1
X_15686_ _15683_/Y _15684_/X _15520_/X _15522_/X vssd1 vssd1 vccd1 vccd1 _15687_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12898_ _21743_/Q _12897_/C _12897_/D _14367_/A vssd1 vssd1 vccd1 vccd1 _12899_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17425_ _17425_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17427_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_129_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14637_ _15155_/C _15978_/B _14637_/C _14785_/A vssd1 vssd1 vccd1 vccd1 _14785_/B
+ sky130_fd_sc_hd__nand4_2
X_11849_ _11848_/A _11848_/C _11848_/B vssd1 vssd1 vccd1 vccd1 _11854_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14568_ _14568_/A _14568_/B _14568_/C vssd1 vssd1 vccd1 vccd1 _14568_/Y sky130_fd_sc_hd__nand3_1
X_17356_ _17356_/A _17356_/B _17356_/C _17356_/D vssd1 vssd1 vccd1 vccd1 _17356_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__16508__B1 _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16307_ _16406_/A _16404_/B vssd1 vssd1 vccd1 vccd1 _16308_/B sky130_fd_sc_hd__nand2_1
XANTENNA__19170__B2 _11550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13519_ _13361_/A _13361_/C _13512_/A vssd1 vssd1 vccd1 vccd1 _13520_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_42_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14499_ _14813_/A _14659_/A _15112_/D vssd1 vssd1 vccd1 vccd1 _14499_/X sky130_fd_sc_hd__and3_1
X_17287_ _17288_/A _17288_/B vssd1 vssd1 vccd1 vccd1 _17404_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19026_ _19023_/X _19024_/Y _18859_/D _18860_/B vssd1 vssd1 vccd1 vccd1 _19043_/B
+ sky130_fd_sc_hd__a211oi_2
X_16238_ _16119_/B _16120_/Y _16235_/A _16237_/Y vssd1 vssd1 vccd1 vccd1 _16348_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14534__A2 _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16169_ _16169_/A _16169_/B vssd1 vssd1 vccd1 vccd1 _16170_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18801__D _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19185__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16602__C _17443_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14298__A1 _12291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19928_ _19928_/A _19928_/B vssd1 vssd1 vccd1 vccd1 _19929_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__19225__A2 _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19859_ _19961_/A _20381_/A _19857_/Y _19858_/X vssd1 vssd1 vccd1 vccd1 _19863_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_138_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17787__A2 _17924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20791__A1 _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20791__B2 _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12858__B _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21821_ _21821_/CLK _21821_/D vssd1 vssd1 vccd1 vccd1 hold327/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__15234__B _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout261_A _19823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13680__D _14635_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18736__A1 _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout359_A _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18736__B2 _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21752_ _22049_/CLK _21752_/D vssd1 vssd1 vccd1 vccd1 _21752_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20543__A1 _20991_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18545__B _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20703_ _20705_/A vssd1 vssd1 vccd1 vccd1 _20836_/A sky130_fd_sc_hd__inv_2
XFILLER_0_149_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21683_ _21939_/CLK _21683_/D vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout526_A _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11036__A1 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20634_ _20501_/Y _20503_/Y _20632_/Y _20633_/X vssd1 vssd1 vccd1 vccd1 _20634_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_149_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20565_ _20565_/A _20685_/B vssd1 vssd1 vccd1 vccd1 _20567_/B sky130_fd_sc_hd__or2_1
XFILLER_0_62_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17711__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20496_ _20496_/A _20496_/B vssd1 vssd1 vccd1 vccd1 _20498_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_143_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18711__D _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17608__C _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21117_ _21188_/A _21116_/C _21116_/A vssd1 vssd1 vccd1 vccd1 _21117_/X sky130_fd_sc_hd__o21a_1
XANTENNA__19392__A _19692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22097_ _22105_/CLK _22097_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[33] sky130_fd_sc_hd__dfrtp_4
Xfanout230 _20273_/A vssd1 vssd1 vccd1 vccd1 _21296_/A sky130_fd_sc_hd__buf_4
Xfanout241 _21293_/A vssd1 vssd1 vccd1 vccd1 _20863_/C sky130_fd_sc_hd__buf_4
XANTENNA__19823__C _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout252 hold330/X vssd1 vssd1 vccd1 vccd1 _17334_/B sky130_fd_sc_hd__buf_4
X_21048_ _21048_/A _21048_/B vssd1 vssd1 vccd1 vccd1 _21050_/B sky130_fd_sc_hd__or2_1
Xfanout263 _21802_/Q vssd1 vssd1 vccd1 vccd1 _17433_/A sky130_fd_sc_hd__clkbuf_8
Xfanout274 _21800_/Q vssd1 vssd1 vccd1 vccd1 _17525_/A sky130_fd_sc_hd__buf_2
Xfanout285 _19487_/A vssd1 vssd1 vccd1 vccd1 _20032_/D sky130_fd_sc_hd__buf_4
XFILLER_0_156_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout296 _21796_/Q vssd1 vssd1 vccd1 vccd1 _18873_/A sky130_fd_sc_hd__clkbuf_8
X_13870_ _13868_/X _13870_/B vssd1 vssd1 vccd1 vccd1 _13871_/B sky130_fd_sc_hd__nand2b_1
X_12821_ _12831_/D _12831_/C _12947_/A vssd1 vssd1 vccd1 vccd1 _12822_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_1146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15540_ _15540_/A _15663_/B vssd1 vssd1 vccd1 vccd1 _15543_/A sky130_fd_sc_hd__or2_1
XFILLER_0_139_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12752_ _12877_/B _13152_/C _13152_/D _12637_/A vssd1 vssd1 vccd1 vccd1 _12752_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1023 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17997__D _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11703_ _11650_/A _11652_/B _12297_/A _11702_/Y vssd1 vssd1 vccd1 vccd1 _12297_/B
+ sky130_fd_sc_hd__a211oi_4
X_15471_ _15287_/Y _15289_/Y _15469_/Y _15470_/X vssd1 vssd1 vccd1 vccd1 _15473_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_84_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ _12572_/A _12572_/C _12572_/B vssd1 vssd1 vccd1 vccd1 _12684_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__12784__A _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14422_ _14422_/A _14422_/B vssd1 vssd1 vccd1 vccd1 _14423_/B sky130_fd_sc_hd__xor2_4
XANTENNA__11027__A1 hold247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17210_ _17210_/A _17210_/B vssd1 vssd1 vccd1 vccd1 _17213_/A sky130_fd_sc_hd__xnor2_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ _11683_/B _11631_/X _11625_/X _11787_/A vssd1 vssd1 vccd1 vccd1 _11635_/B
+ sky130_fd_sc_hd__a211o_1
X_18190_ _18789_/A _19089_/B _18187_/Y _18332_/A vssd1 vssd1 vccd1 vccd1 _18192_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14353_ _15695_/A _14508_/A _14354_/C _14817_/D vssd1 vssd1 vccd1 vccd1 _14353_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_108_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17141_ _17141_/A _17141_/B _17141_/C _17493_/A vssd1 vssd1 vccd1 vccd1 _17141_/X
+ sky130_fd_sc_hd__and4_1
X_11565_ _12750_/A _11564_/X _11563_/X vssd1 vssd1 vccd1 vccd1 _11566_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ _13304_/A _13304_/B _13304_/C vssd1 vssd1 vccd1 vccd1 _13306_/C sky130_fd_sc_hd__nand3_2
X_17072_ _17071_/B _17071_/C _17071_/A vssd1 vssd1 vccd1 vccd1 _17073_/C sky130_fd_sc_hd__a21bo_1
X_14284_ _14284_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14289_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11496_ _11502_/A1 t2x[15] v1z[15] fanout20/X _11495_/X vssd1 vssd1 vccd1 vccd1 _11496_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16023_ _16023_/A _16143_/B vssd1 vssd1 vccd1 vccd1 _21409_/B sky130_fd_sc_hd__or2_2
X_13235_ _13376_/A _13234_/Y _13394_/A _16328_/B vssd1 vssd1 vccd1 vccd1 _13376_/B
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__17087__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_990 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13166_ _13166_/A _13166_/B _13166_/C vssd1 vssd1 vccd1 vccd1 _13168_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_27_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12117_ _12020_/A _12302_/A _12312_/A _12326_/D vssd1 vssd1 vccd1 vccd1 _12118_/B
+ sky130_fd_sc_hd__a22oi_1
X_13097_ _13097_/A _13097_/B vssd1 vssd1 vccd1 vccd1 _13111_/A sky130_fd_sc_hd__and2_1
X_17974_ _17967_/A _17967_/B _17968_/Y vssd1 vssd1 vccd1 vccd1 _18101_/A sky130_fd_sc_hd__a21oi_2
X_19713_ _19711_/A _19711_/B _19711_/C vssd1 vssd1 vccd1 vccd1 _19715_/C sky130_fd_sc_hd__a21o_1
X_16925_ _17144_/A _17129_/B _17013_/C _17013_/D vssd1 vssd1 vccd1 vccd1 _16926_/B
+ sky130_fd_sc_hd__and4_1
X_12048_ _12048_/A _12048_/B vssd1 vssd1 vccd1 vccd1 _12050_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__21337__A _21349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19644_ _19644_/A _20032_/D _20838_/C _20838_/D vssd1 vssd1 vccd1 vccd1 _19645_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__21056__B _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16856_ _17165_/C _17168_/A _17165_/A _17165_/B vssd1 vssd1 vccd1 vccd1 _17372_/B
+ sky130_fd_sc_hd__o211ai_4
X_15807_ _15808_/C _16414_/B _15805_/Y _15927_/A vssd1 vssd1 vccd1 vccd1 _15809_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_19575_ _20650_/A _19866_/C _19575_/C _19575_/D vssd1 vssd1 vccd1 vccd1 _19575_/Y
+ sky130_fd_sc_hd__nand4_2
X_16787_ _16778_/X _16785_/X _16786_/X _16718_/Y vssd1 vssd1 vccd1 vccd1 _16790_/A
+ sky130_fd_sc_hd__o211ai_4
X_13999_ _14306_/A _14155_/D _13999_/C _14153_/A vssd1 vssd1 vccd1 vccd1 _14153_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12397__C _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18526_ _18542_/B _18525_/B _18525_/C _18525_/D vssd1 vssd1 vccd1 vccd1 _18526_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11266__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15738_ _15741_/C vssd1 vssd1 vccd1 vccd1 _15738_/Y sky130_fd_sc_hd__inv_2
XTAP_3190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11266__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20525__A1 _20249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19391__A1 _19692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18457_ _18454_/Y _18455_/X _18327_/X _18330_/Y vssd1 vssd1 vccd1 vccd1 _18457_/Y
+ sky130_fd_sc_hd__o211ai_4
X_15669_ _15669_/A _15669_/B vssd1 vssd1 vccd1 vccd1 _15680_/A sky130_fd_sc_hd__or2_1
XANTENNA_190 hold247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15070__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17408_ _17405_/Y _17406_/X _17316_/X _17319_/Y vssd1 vssd1 vccd1 vccd1 _17409_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18388_ _18388_/A _18388_/B vssd1 vssd1 vccd1 vccd1 _18389_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17339_ _17557_/B _17915_/D _17924_/B _17557_/A vssd1 vssd1 vccd1 vccd1 _17340_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20350_ _20498_/B _20350_/B vssd1 vssd1 vccd1 vccd1 _20352_/B sky130_fd_sc_hd__nor2_1
XANTENNA__15704__B2 _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20416__A _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19009_ _19008_/D _19185_/B _21261_/B _18857_/B vssd1 vssd1 vccd1 vccd1 _19010_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_141_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20281_ _20281_/A _20281_/B vssd1 vssd1 vccd1 vccd1 _20292_/A sky130_fd_sc_hd__or2_1
XANTENNA_fanout107_A _21267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22020_ _22020_/CLK _22020_/D vssd1 vssd1 vccd1 vccd1 hold179/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__15229__B _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14133__B _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold49/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout476_A _15093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18957__B2 _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout643_A _21329_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11257__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21804_ _22021_/CLK _21804_/D vssd1 vssd1 vccd1 vccd1 hold322/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20516__A1 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21735_ _21803_/CLK _21735_/D vssd1 vssd1 vccd1 vccd1 _21735_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_93_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16507__C _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21666_ _21906_/CLK _21666_/D vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold319_A hold319/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14308__B _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12757__A1 _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20617_ _20480_/Y _20484_/A _20614_/Y _20616_/X vssd1 vssd1 vccd1 vccd1 _20617_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15130__D _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21597_ _21888_/CLK _21597_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[60] sky130_fd_sc_hd__dfrtp_4
XANTENNA__19685__A2 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11350_ _11544_/A1 t1x[31] v2z[31] _11543_/B2 _11349_/X vssd1 vssd1 vccd1 vccd1 _11350_/X
+ sky130_fd_sc_hd__a221o_4
XFILLER_0_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20548_ _20679_/A vssd1 vssd1 vccd1 vccd1 _20550_/D sky130_fd_sc_hd__inv_2
XANTENNA__17619__B _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12509__A1 _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11281_ _11325_/A1 t2y[14] t0y[14] _11507_/A1 vssd1 vssd1 vccd1 vccd1 _11281_/X sky130_fd_sc_hd__a22o_1
XANTENNA__19437__A2 _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20479_ _20479_/A _20602_/B vssd1 vssd1 vccd1 vccd1 _20481_/B sky130_fd_sc_hd__or2_1
XFILLER_0_120_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17338__C _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13182__A1 _14712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13020_ _13020_/A _13020_/B _13020_/C vssd1 vssd1 vccd1 vccd1 _13023_/A sky130_fd_sc_hd__nand3_1
XANTENNA__13182__B2 _14712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11159__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14971_ _14974_/A _14974_/B _14971_/C vssd1 vssd1 vccd1 vccd1 _15085_/A sky130_fd_sc_hd__and3_2
XFILLER_0_22_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18948__A1 _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16710_ _16715_/A _16493_/Y _16492_/X _16484_/X vssd1 vssd1 vccd1 vccd1 _16712_/D
+ sky130_fd_sc_hd__a211o_1
X_13922_ _13920_/Y _13921_/X _14848_/A _14234_/C vssd1 vssd1 vccd1 vccd1 _13924_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_96_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11496__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17690_ _17689_/A _17689_/B _17689_/C _17689_/D vssd1 vssd1 vccd1 vccd1 _17690_/Y
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__11496__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17620__A1 _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16641_ _16622_/A _16622_/C _16622_/B vssd1 vssd1 vccd1 vccd1 _16642_/C sky130_fd_sc_hd__a21o_1
X_13853_ _13736_/Y _13739_/Y _13973_/B _13852_/X vssd1 vssd1 vccd1 vccd1 _13972_/A
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__17620__B2 _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19360_ _19204_/B _19206_/B _19519_/A _19359_/Y vssd1 vssd1 vccd1 vccd1 _19519_/B
+ sky130_fd_sc_hd__a211oi_1
X_12804_ _12803_/A _12803_/B _12803_/C _12803_/D vssd1 vssd1 vccd1 vccd1 _12804_/Y
+ sky130_fd_sc_hd__o22ai_4
X_16572_ _16572_/A _16572_/B vssd1 vssd1 vccd1 vccd1 _16580_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12445__B1 _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13784_ _13784_/A _13784_/B _13784_/C vssd1 vssd1 vccd1 vccd1 _13787_/A sky130_fd_sc_hd__nand3_1
X_10996_ mstream_o[70] hold42/X _11005_/S vssd1 vssd1 vccd1 vccd1 _21607_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_97_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18311_ _18307_/X _18308_/Y _18157_/A _18157_/Y vssd1 vssd1 vccd1 vccd1 _18373_/B
+ sky130_fd_sc_hd__a211oi_2
X_15523_ _15523_/A _15523_/B vssd1 vssd1 vccd1 vccd1 _15525_/B sky130_fd_sc_hd__xor2_1
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18616__D _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19291_ _19291_/A _19291_/B vssd1 vssd1 vccd1 vccd1 _19292_/B sky130_fd_sc_hd__xor2_2
X_12735_ _12856_/A _12734_/Y _13556_/A _13573_/D vssd1 vssd1 vccd1 vccd1 _12856_/B
+ sky130_fd_sc_hd__and4bb_1
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17520__D _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18242_ _17967_/A _17967_/B _18100_/A vssd1 vssd1 vccd1 vccd1 _18242_/Y sky130_fd_sc_hd__a21boi_2
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15454_ _16087_/A _15695_/A _15717_/C _15976_/D vssd1 vssd1 vccd1 vccd1 _15587_/A
+ sky130_fd_sc_hd__and4_1
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ _12667_/A _12667_/B vssd1 vssd1 vccd1 vccd1 _12766_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_26_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14218__B _14218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14405_ _14557_/B _15001_/B _15510_/B _14557_/A vssd1 vssd1 vccd1 vccd1 _14408_/C
+ sky130_fd_sc_hd__a22o_1
X_11617_ _12302_/A _12858_/C _12991_/D _12269_/D vssd1 vssd1 vccd1 vccd1 _11617_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_142_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18173_ _19379_/B _18624_/A _18170_/Y _18322_/A vssd1 vssd1 vccd1 vccd1 _18174_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_26_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15385_ _15386_/B _15386_/C _15386_/A vssd1 vssd1 vccd1 vccd1 _15385_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_52_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12597_ _12708_/A _12708_/B _12825_/A vssd1 vssd1 vccd1 vccd1 _12598_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_136_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17124_ _17146_/A _17146_/B _17124_/C _17141_/C vssd1 vssd1 vccd1 vccd1 _17126_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11420__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14336_ _14489_/A _14334_/Y _14160_/B _14162_/B vssd1 vssd1 vccd1 vccd1 _14337_/B
+ sky130_fd_sc_hd__o211ai_1
X_11548_ _11549_/A hold2/A vssd1 vssd1 vccd1 vccd1 _11548_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14267_ _14264_/Y _14265_/X _14105_/B _14105_/Y vssd1 vssd1 vccd1 vccd1 _14268_/C
+ sky130_fd_sc_hd__a211o_1
X_17055_ _17096_/A _17146_/C vssd1 vssd1 vccd1 vccd1 _17069_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_122_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11479_ _11478_/X _18319_/B _11521_/S vssd1 vssd1 vccd1 vccd1 _21831_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_64_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14234__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16006_ _16003_/Y _16004_/X _15876_/X _15878_/Y vssd1 vssd1 vccd1 vccd1 _16007_/B
+ sky130_fd_sc_hd__a211o_1
X_13218_ _13218_/A _13218_/B _13218_/C vssd1 vssd1 vccd1 vccd1 _13218_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__11577__B _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14198_ _14198_/A _14198_/B _14198_/C vssd1 vssd1 vccd1 vccd1 _14201_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_20_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13149_ _13040_/A _13040_/C _13040_/B vssd1 vssd1 vccd1 vccd1 _13164_/A sky130_fd_sc_hd__a21bo_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14249__B1_N hold313/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17957_ _17953_/X _17954_/Y _17812_/X _17815_/X vssd1 vssd1 vccd1 vccd1 _17958_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14673__A1 _14828_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14673__B2 _16173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16908_ _16909_/A _16908_/B _16908_/C vssd1 vssd1 vccd1 vccd1 _16916_/A sky130_fd_sc_hd__nand3_1
XANTENNA__11487__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17888_ _17747_/Y _17750_/X _17975_/A _17887_/Y vssd1 vssd1 vccd1 vccd1 _17975_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__21628__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_7 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19627_ _19465_/A _19465_/B _19463_/Y vssd1 vssd1 vccd1 vccd1 _19629_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__12839__D _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16839_ _16840_/A _16840_/B _16840_/C vssd1 vssd1 vccd1 vccd1 _16849_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_88_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11239__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19558_ _19424_/B _19426_/A _19556_/X _19557_/Y vssd1 vssd1 vccd1 vccd1 _19560_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_76_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18509_ _18508_/A _18508_/B _18508_/C vssd1 vssd1 vccd1 vccd1 _18511_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19489_ _19650_/D _20841_/B vssd1 vssd1 vccd1 vccd1 _19490_/B sky130_fd_sc_hd__nand2_2
XANTENNA__17375__B1 _21337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17914__A2 _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21520_ hold258/X sstream_i[97] _21528_/S vssd1 vssd1 vccd1 vccd1 _22047_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_63_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21451_ hold214/X sstream_i[28] _21481_/S vssd1 vssd1 vccd1 vccd1 _21978_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout224_A _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20402_ _20403_/B _20403_/A vssd1 vssd1 vccd1 vccd1 _20402_/X sky130_fd_sc_hd__and2b_1
XANTENNA__11411__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21382_ _14605_/B _19476_/Y _21420_/S vssd1 vssd1 vccd1 vccd1 _21382_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20146__A _20689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20333_ _20838_/B _20975_/D _21283_/B _21305_/B vssd1 vssd1 vccd1 vccd1 _20472_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_113_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16062__C _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20264_ _21291_/A _21278_/A _21301_/A _20863_/C vssd1 vssd1 vccd1 vccd1 _20267_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_347 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout593_A _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22003_ _22005_/CLK _22003_/D vssd1 vssd1 vccd1 vccd1 hold131/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13983__A _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19373__C _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20195_ _20196_/A _20196_/B vssd1 vssd1 vccd1 vccd1 _20195_/X sky130_fd_sc_hd__or2_1
XANTENNA__14664__A1 _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11478__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11478__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12675__B1 _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15704__A2_N _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10850_ _10805_/Y _11066_/A _10802_/X _10859_/A vssd1 vssd1 vccd1 vccd1 _10859_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_79_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17621__C _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_142 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12520_ _12521_/A _12521_/B _12521_/C vssd1 vssd1 vccd1 vccd1 _12522_/B sky130_fd_sc_hd__a21oi_4
X_21718_ _21724_/CLK _21718_/D _21422_/A vssd1 vssd1 vccd1 vccd1 _21718_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12451_ _12451_/A _12451_/B vssd1 vssd1 vccd1 vccd1 _12471_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_136_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21649_ _21722_/CLK _21649_/D fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[112]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11402_ _11124_/A hold282/A fanout47/X hold154/A vssd1 vssd1 vccd1 vccd1 _11402_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15170_ _15017_/A _15019_/B _15017_/B vssd1 vssd1 vccd1 vccd1 _15175_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__13877__B _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12382_ _12379_/Y _12380_/X _11802_/X _11805_/X vssd1 vssd1 vccd1 vccd1 _12382_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_90 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14121_ _14121_/A _14121_/B _13834_/A vssd1 vssd1 vccd1 vccd1 _14285_/B sky130_fd_sc_hd__or3b_2
XFILLER_0_104_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20673__B1 _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11333_ _11349_/A1 t2y[27] t0y[27] _21723_/D vssd1 vssd1 vccd1 vccd1 _11333_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_22_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18171__D _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13596__C _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14052_ _13919_/A _13918_/B _13916_/X vssd1 vssd1 vccd1 vccd1 _14068_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_104_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11264_ _12020_/A _11263_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21767_/D sky130_fd_sc_hd__mux2_1
X_13003_ _13003_/A vssd1 vssd1 vccd1 vccd1 _13003_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13893__A _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18860_ _18860_/A _18860_/B vssd1 vssd1 vccd1 vccd1 _18861_/A sky130_fd_sc_hd__or2_1
X_11195_ _14391_/B _11194_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21748_/D sky130_fd_sc_hd__mux2_1
XANTENNA__20976__B2 _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17811_ _17810_/B _17810_/C _17810_/A vssd1 vssd1 vccd1 vccd1 _17811_/Y sky130_fd_sc_hd__o21ai_2
X_18791_ _18790_/B _18947_/B _18790_/A vssd1 vssd1 vccd1 vccd1 _18792_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14501__B _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17742_ _21796_/Q _17741_/B _17870_/A _17741_/D vssd1 vssd1 vccd1 vccd1 _17743_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11469__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14954_ _14954_/A _14954_/B _14954_/C vssd1 vssd1 vccd1 vccd1 _14956_/B sky130_fd_sc_hd__nand3_2
XANTENNA__12302__A _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21037__D _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21721__RESET_B _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13905_ _14051_/A _13904_/C _13904_/A vssd1 vssd1 vccd1 vccd1 _13906_/C sky130_fd_sc_hd__a21o_1
X_17673_ _17673_/A _17673_/B _17673_/C vssd1 vssd1 vccd1 vccd1 _17676_/A sky130_fd_sc_hd__nand3_1
XANTENNA__14407__A1 _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14885_ _14705_/B _14707_/B _14883_/X _14884_/Y vssd1 vssd1 vccd1 vccd1 _14887_/C
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__18196__A _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19412_ _19412_/A _19412_/B vssd1 vssd1 vccd1 vccd1 _19420_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_134_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16624_ _16613_/A _16613_/C _16613_/B vssd1 vssd1 vccd1 vccd1 _16625_/C sky130_fd_sc_hd__a21o_1
X_13836_ _14306_/A _14477_/C _14155_/D _14138_/A vssd1 vssd1 vccd1 vccd1 _13839_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21334__B _21334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11860__B _12621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19343_ _19343_/A _19343_/B vssd1 vssd1 vccd1 vccd1 _19345_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16555_ _16870_/A _17223_/A vssd1 vssd1 vccd1 vccd1 _16644_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13767_ _13767_/A _13767_/B _13910_/B vssd1 vssd1 vccd1 vccd1 _13767_/X sky130_fd_sc_hd__and3_1
X_10979_ mstream_o[61] _10978_/Y _11005_/S vssd1 vssd1 vccd1 vccd1 _21598_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_130_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11352__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15506_ _15220_/B _15362_/B _15218_/X vssd1 vssd1 vccd1 vccd1 _16031_/A sky130_fd_sc_hd__a21o_4
XFILLER_0_57_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19274_ _19270_/X _19272_/Y _19099_/B _19101_/B vssd1 vssd1 vccd1 vccd1 _19275_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_45_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12718_ _13983_/B _14176_/C _13402_/D _13394_/A vssd1 vssd1 vccd1 vccd1 _12719_/A
+ sky130_fd_sc_hd__a22o_1
X_16486_ _17300_/C _17282_/A _17277_/A _17520_/D vssd1 vssd1 vccd1 vccd1 _16489_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13698_ _13698_/A _13698_/B _13698_/C vssd1 vssd1 vccd1 vccd1 _13698_/X sky130_fd_sc_hd__or3_2
XFILLER_0_85_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_19_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21682_/CLK sky130_fd_sc_hd__clkbuf_16
X_18225_ _18225_/A _18225_/B _18225_/C vssd1 vssd1 vccd1 vccd1 _18225_/X sky130_fd_sc_hd__or3_2
XFILLER_0_66_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15437_ _15437_/A _15437_/B vssd1 vssd1 vccd1 vccd1 _15438_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_5_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12649_ _12649_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _12651_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_115_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18156_ _18304_/B _18155_/B _18155_/C vssd1 vssd1 vccd1 vccd1 _18157_/B sky130_fd_sc_hd__a21oi_2
X_15368_ _15892_/A _15632_/B _15510_/B _15368_/D vssd1 vssd1 vccd1 vccd1 _15548_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_87_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16163__B _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17107_ _17106_/A _17120_/A _17078_/X _17083_/Y vssd1 vssd1 vccd1 vccd1 _17156_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold305 hold305/A vssd1 vssd1 vccd1 vccd1 hold305/X sky130_fd_sc_hd__dlygate4sd3_1
X_14319_ _14319_/A _14319_/B vssd1 vssd1 vccd1 vccd1 _14321_/B sky130_fd_sc_hd__or2_2
Xhold316 hold316/A vssd1 vssd1 vccd1 vccd1 hold316/X sky130_fd_sc_hd__dlygate4sd3_1
X_18087_ _18107_/B _18087_/B _18087_/C _18087_/D vssd1 vssd1 vccd1 vccd1 _18087_/X
+ sky130_fd_sc_hd__or4_2
X_15299_ _15702_/D _15829_/C _15954_/D _15435_/A vssd1 vssd1 vccd1 vccd1 _15303_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold327 hold327/A vssd1 vssd1 vccd1 vccd1 hold327/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17038_ _17038_/A _17038_/B _17038_/C vssd1 vssd1 vccd1 vccd1 _17038_/X sky130_fd_sc_hd__or3_2
XFILLER_0_1_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11738__D _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19821__A2 _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20413__B _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16610__C _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18989_ _18826_/C _18826_/Y _18987_/X _18988_/X vssd1 vssd1 vccd1 vccd1 _18991_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11527__S _11545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20951_ _20951_/A _20951_/B _20951_/C vssd1 vssd1 vccd1 vccd1 _20952_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_75_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21392__A1 _21390_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout174_A _18058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16619__A _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15523__A _15523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20882_ _20883_/A _20883_/B vssd1 vssd1 vccd1 vccd1 _20882_/Y sky130_fd_sc_hd__nand2_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15071__B2 fanout6/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18256__D _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13621__A2 _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout439_A _21761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13043__A _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21503_ hold285/X sstream_i[80] _21507_/S vssd1 vssd1 vccd1 vccd1 _22030_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_75_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12882__A _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21434_ hold244/X sstream_i[11] _21442_/S vssd1 vssd1 vccd1 vccd1 _21961_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18848__B1 _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18312__A2 _18929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__B1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19087__D _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21365_ _21412_/A _18537_/Y _21421_/S _21364_/Y vssd1 vssd1 vccd1 vccd1 _21365_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20316_ _20316_/A _20316_/B vssd1 vssd1 vccd1 vccd1 _20321_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_102_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20026__D _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21296_ _21296_/A _21296_/B vssd1 vssd1 vccd1 vccd1 _21297_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14024__D _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20247_ _21831_/Q _21832_/Q _20247_/C _20247_/D vssd1 vssd1 vccd1 vccd1 _20248_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA_fanout87_A _19053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20178_ _20032_/D _20178_/B _20721_/C _20178_/D vssd1 vssd1 vccd1 vccd1 _20328_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_122_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13863__D _14663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11951_ _12020_/A _12402_/A _12302_/A _12326_/D vssd1 vssd1 vccd1 vccd1 _11952_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21383__A1 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16529__A _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10902_ _10902_/A _10902_/B _10902_/C vssd1 vssd1 vccd1 vccd1 _10903_/B sky130_fd_sc_hd__and3_1
XTAP_3778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14670_ _14670_/A _14670_/B vssd1 vssd1 vccd1 vccd1 _14684_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_93_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11882_ _12319_/C _12302_/A _12312_/A _12420_/D vssd1 vssd1 vccd1 vccd1 _11883_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13621_ _14713_/B _14077_/B _14234_/C _14713_/A vssd1 vssd1 vccd1 vccd1 _13622_/B
+ sky130_fd_sc_hd__a22o_1
X_10833_ _11050_/B _11051_/A _11050_/A vssd1 vssd1 vccd1 vccd1 _11053_/B sky130_fd_sc_hd__o21ba_2
XANTENNA__11680__B _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18166__D _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17339__B1 _17924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13612__A2 _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16340_ _16340_/A _16340_/B vssd1 vssd1 vccd1 vccd1 _16341_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_149_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13552_ _13548_/A _13549_/X _13392_/Y _13395_/X vssd1 vssd1 vccd1 vccd1 _13652_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18585__A2_N _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12503_ _12503_/A _12503_/B vssd1 vssd1 vccd1 vccd1 _12505_/A sky130_fd_sc_hd__nand2_1
X_16271_ _16380_/A _16371_/A _16369_/B vssd1 vssd1 vccd1 vccd1 _16271_/X sky130_fd_sc_hd__and3_1
XFILLER_0_125_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13483_ _13483_/A _13483_/B _13483_/C vssd1 vssd1 vccd1 vccd1 _13486_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_54_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16562__A1 _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18010_ _18010_/A _20148_/C _18144_/A _18010_/D vssd1 vssd1 vccd1 vccd1 _18144_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_63_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15222_ _15363_/A _15222_/B vssd1 vssd1 vccd1 vccd1 _15225_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_63_871 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12434_ _12435_/A _12435_/B vssd1 vssd1 vccd1 vccd1 _12434_/X sky130_fd_sc_hd__and2_2
XFILLER_0_129_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15117__A2 _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15153_ _15435_/A _15153_/B _15829_/C _15954_/D vssd1 vssd1 vccd1 vccd1 _15305_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__19575__A _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12365_ _12364_/B _12364_/C _12364_/A vssd1 vssd1 vccd1 vccd1 _12367_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_121_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14104_ _14100_/X _14102_/Y _13939_/B _13939_/Y vssd1 vssd1 vccd1 vccd1 _14105_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14325__B1 _14635_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11316_ _13402_/D _11315_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21780_/D sky130_fd_sc_hd__mux2_1
X_15084_ _15085_/A _15502_/A _15085_/C _15085_/D vssd1 vssd1 vccd1 vccd1 _15087_/A
+ sky130_fd_sc_hd__o22ai_1
X_19961_ _19961_/A _20381_/A _19961_/C _19961_/D vssd1 vssd1 vccd1 vccd1 _20095_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_61_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12296_ _12289_/A _12289_/B _12294_/X vssd1 vssd1 vccd1 vccd1 _12296_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13679__A2 _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14035_ _14365_/A _21742_/Q _14537_/A _14516_/A vssd1 vssd1 vccd1 vccd1 _14190_/A
+ sky130_fd_sc_hd__nand4_2
X_18912_ _18912_/A _18912_/B _19065_/B vssd1 vssd1 vccd1 vccd1 _18914_/B sky130_fd_sc_hd__nand3_1
X_11247_ fanout59/X v0z[5] fanout19/X _11246_/X vssd1 vssd1 vccd1 vccd1 _11247_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17095__A _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19892_ _19892_/A _20671_/B vssd1 vssd1 vccd1 vccd1 _19893_/B sky130_fd_sc_hd__and2_1
XANTENNA__17526__C _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19803__A2 _20841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18843_ hold47/X fanout8/X _13967_/X _11550_/B _18842_/Y vssd1 vssd1 vccd1 vccd1
+ _18843_/X sky130_fd_sc_hd__a221o_1
X_11178_ hold279/X fanout51/X fanout47/X hold311/A vssd1 vssd1 vccd1 vccd1 _11178_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18774_ _18775_/A _18775_/B _18775_/C vssd1 vssd1 vccd1 vccd1 _18774_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_59_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15986_ _15986_/A _15986_/B _15986_/C vssd1 vssd1 vccd1 vccd1 _15986_/X sky130_fd_sc_hd__and3_1
XFILLER_0_98_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18638__B _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12103__A2 _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19567__A1 _19868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17725_ _17725_/A _17725_/B vssd1 vssd1 vccd1 vccd1 _17736_/A sky130_fd_sc_hd__or2_1
X_14937_ _14939_/A vssd1 vssd1 vccd1 vccd1 _15167_/A sky130_fd_sc_hd__inv_2
XANTENNA__17542__B _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21374__A1 _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11311__B1 _11310_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17656_ _17434_/B _19432_/A _17544_/X _17543_/X _19951_/A vssd1 vssd1 vccd1 vccd1
+ _17664_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14868_ _14868_/A _14868_/B _14868_/C vssd1 vssd1 vccd1 vccd1 _14887_/B sky130_fd_sc_hd__and3_1
X_16607_ _17557_/A _17915_/A _17557_/B _17657_/A vssd1 vssd1 vccd1 vccd1 _16608_/C
+ sky130_fd_sc_hd__a22o_1
X_13819_ _13819_/A _13819_/B vssd1 vssd1 vccd1 vccd1 _13956_/A sky130_fd_sc_hd__nor2_1
X_17587_ _17475_/A _17474_/B _17474_/A vssd1 vssd1 vccd1 vccd1 _17589_/B sky130_fd_sc_hd__o21bai_4
X_14799_ _14797_/Y _14799_/B vssd1 vssd1 vccd1 vccd1 _14802_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_9_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19326_ _19194_/A _19193_/Y _19192_/B vssd1 vssd1 vccd1 vccd1 _19469_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_85_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16538_ _16680_/A _16680_/B _16537_/A vssd1 vssd1 vccd1 vccd1 _16552_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21080__A _21293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19257_ _20101_/A _20101_/B _19703_/C _19906_/C vssd1 vssd1 vccd1 vccd1 _19258_/B
+ sky130_fd_sc_hd__nand4_1
X_16469_ _17300_/C _17124_/C _17282_/A _17520_/D vssd1 vssd1 vccd1 vccd1 _16472_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18208_ _18207_/A _18207_/B _18207_/C vssd1 vssd1 vccd1 vccd1 _18209_/C sky130_fd_sc_hd__a21o_1
XANTENNA__14564__B1 _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19188_ _19188_/A _19188_/B vssd1 vssd1 vccd1 vccd1 _19189_/B sky130_fd_sc_hd__nor2_1
XANTENNA__14406__B _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18139_ _17999_/A _17999_/C _17999_/B vssd1 vssd1 vccd1 vccd1 _18140_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold102 hold102/A vssd1 vssd1 vccd1 vccd1 hold102/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 hold113/A vssd1 vssd1 vccd1 vccd1 hold113/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 hold124/A vssd1 vssd1 vccd1 vccd1 hold124/X sky130_fd_sc_hd__dlygate4sd3_1
X_21150_ _21301_/A _21264_/B _21046_/B _21151_/A vssd1 vssd1 vccd1 vccd1 _21150_/X
+ sky130_fd_sc_hd__a22o_1
Xhold135 hold135/A vssd1 vssd1 vccd1 vccd1 hold135/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold146 hold146/A vssd1 vssd1 vccd1 vccd1 hold146/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 hold157/A vssd1 vssd1 vccd1 vccd1 hold157/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 hold168/A vssd1 vssd1 vccd1 vccd1 hold168/X sky130_fd_sc_hd__dlygate4sd3_1
X_20101_ _20101_/A _20101_/B _21816_/Q _21817_/Q vssd1 vssd1 vccd1 vccd1 _20282_/A
+ sky130_fd_sc_hd__nand4_2
Xhold179 hold179/A vssd1 vssd1 vccd1 vccd1 hold179/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21081_ _21194_/A vssd1 vssd1 vccd1 vccd1 _21083_/D sky130_fd_sc_hd__inv_2
Xfanout604 _11459_/B2 vssd1 vssd1 vccd1 vccd1 _11223_/A sky130_fd_sc_hd__buf_4
XFILLER_0_42_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout615 _21568_/S vssd1 vssd1 vccd1 vccd1 _10992_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_95_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout626 _21087_/D vssd1 vssd1 vccd1 vccd1 _19695_/A sky130_fd_sc_hd__clkbuf_8
X_20032_ _19810_/D _20178_/B _20721_/C _20032_/D vssd1 vssd1 vccd1 vccd1 _20035_/A
+ sky130_fd_sc_hd__and4b_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout637 _11089_/A vssd1 vssd1 vccd1 vccd1 fanout637/X sky130_fd_sc_hd__clkbuf_8
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20005__A2_N _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout291_A _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20797__C _21815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21983_ _22016_/CLK _21983_/D vssd1 vssd1 vccd1 vccd1 hold213/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21365__A1 _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20934_ _21110_/A _20934_/B vssd1 vssd1 vccd1 vccd1 _20936_/B sky130_fd_sc_hd__nand2_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20865_ _20866_/B _20866_/A vssd1 vssd1 vccd1 vccd1 _20865_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20192__A1_N _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20796_ _21258_/A _21264_/B _21046_/B _20797_/A vssd1 vssd1 vccd1 vccd1 _20800_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19379__B _19379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18283__B _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19730__A1 _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13858__D _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21417_ hold189/X fanout40/X _21415_/X _21416_/Y vssd1 vssd1 vccd1 vccd1 _21947_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11659__C _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16812__A _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14035__C _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ _12150_/A _12150_/B _12150_/C vssd1 vssd1 vccd1 vccd1 _12160_/A sky130_fd_sc_hd__and3_1
XFILLER_0_60_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21348_ hold163/X _21381_/B _21346_/X _21347_/Y vssd1 vssd1 vccd1 vccd1 _21923_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14858__A1 _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11101_ _10852_/X hold49/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21695_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18049__A1 _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18049__B2 _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12081_ _12078_/Y _12080_/X _12286_/C _12036_/X vssd1 vssd1 vccd1 vccd1 _12081_/X
+ sky130_fd_sc_hd__a211o_1
X_21279_ _21279_/A _21279_/B vssd1 vssd1 vccd1 vccd1 _21280_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_120_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11032_ mstream_o[106] hold299/X _11039_/S vssd1 vssd1 vccd1 vccd1 hold300/A sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15840_ _15971_/A _15841_/C _15841_/A vssd1 vssd1 vccd1 vccd1 _15842_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_21_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17272__A2 _12392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15771_ _15772_/A _16029_/A vssd1 vssd1 vccd1 vccd1 _15904_/B sky130_fd_sc_hd__nor2_1
XTAP_3520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12983_ _12983_/A _12983_/B vssd1 vssd1 vccd1 vccd1 _12986_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__21356__A1 _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17510_ _17510_/A _17510_/B vssd1 vssd1 vccd1 vccd1 _17512_/C sky130_fd_sc_hd__xnor2_1
XTAP_3553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14722_ _14571_/A _14974_/A _14717_/X _14719_/Y vssd1 vssd1 vccd1 vccd1 _14723_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18490_ _18491_/A _18491_/B vssd1 vssd1 vccd1 vccd1 _18632_/B sky130_fd_sc_hd__and2b_1
X_11934_ _12899_/B _12246_/C _11933_/B _11930_/X vssd1 vssd1 vccd1 vccd1 _11940_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_3575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17441_ _17441_/A _17441_/B vssd1 vssd1 vccd1 vccd1 _17461_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_68_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14653_ _14654_/A _14654_/B vssd1 vssd1 vccd1 vccd1 _14764_/B sky130_fd_sc_hd__and2b_1
XTAP_2874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11865_ _11865_/A _11865_/B vssd1 vssd1 vccd1 vccd1 _11867_/B sky130_fd_sc_hd__xnor2_2
XTAP_2885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13604_ _13605_/A _13605_/B _13605_/C vssd1 vssd1 vccd1 vccd1 _13604_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_131_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10816_ hold227/A hold229/A vssd1 vssd1 vccd1 vccd1 _10836_/A sky130_fd_sc_hd__and2_1
X_17372_ _17372_/A _17372_/B _17379_/B vssd1 vssd1 vccd1 vccd1 _17380_/B sky130_fd_sc_hd__or3_1
X_14584_ _14584_/A _14584_/B vssd1 vssd1 vccd1 vccd1 _14587_/A sky130_fd_sc_hd__xnor2_4
X_11796_ _11772_/A _11772_/B _11772_/C vssd1 vssd1 vccd1 vccd1 _11796_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19111_ _19432_/A _19866_/C _19111_/C _19276_/A vssd1 vssd1 vccd1 vccd1 _19276_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_55_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16323_ _16323_/A _16323_/B vssd1 vssd1 vccd1 vccd1 _16333_/A sky130_fd_sc_hd__or2_1
XFILLER_0_131_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13535_ _13536_/A _13536_/B vssd1 vssd1 vccd1 vccd1 _13535_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_32_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14507__A _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20331__A2 _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19042_ _19211_/B _19040_/Y _18878_/X _18881_/A vssd1 vssd1 vccd1 vccd1 _19043_/D
+ sky130_fd_sc_hd__a211oi_2
X_16254_ _16143_/A _16143_/B _16142_/A _16141_/Y vssd1 vssd1 vccd1 vccd1 _16256_/B
+ sky130_fd_sc_hd__o31ai_2
XFILLER_0_153_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13466_ _13466_/A _13466_/B vssd1 vssd1 vccd1 vccd1 _13486_/A sky130_fd_sc_hd__xor2_2
X_15205_ _14910_/A _15068_/A _15068_/B vssd1 vssd1 vccd1 vccd1 _15205_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13130__B _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12417_ _12309_/Y _12312_/X _12415_/X _12416_/Y vssd1 vssd1 vccd1 vccd1 _12479_/A
+ sky130_fd_sc_hd__o211a_1
X_16185_ _16185_/A _16185_/B vssd1 vssd1 vccd1 vccd1 _16185_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_140_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13397_ _13398_/B _13398_/A vssd1 vssd1 vccd1 vccd1 _13523_/A sky130_fd_sc_hd__and2b_1
X_15136_ _15282_/A _15135_/C _15135_/A vssd1 vssd1 vccd1 vccd1 _15138_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_121_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12348_ _12348_/A _12348_/B vssd1 vssd1 vccd1 vccd1 _12350_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__20244__A _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16441__B _16734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11780__B1 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_i_A _21806_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15067_ _15067_/A _15067_/B _15067_/C vssd1 vssd1 vccd1 vccd1 _15068_/B sky130_fd_sc_hd__and3_1
X_12279_ _12241_/X _12275_/X _12277_/X _12278_/Y _12238_/X vssd1 vssd1 vccd1 vccd1
+ _12279_/Y sky130_fd_sc_hd__a2111oi_1
X_19944_ _19944_/A _20081_/B vssd1 vssd1 vccd1 vccd1 _19944_/Y sky130_fd_sc_hd__xnor2_2
XANTENNA__14242__A _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16160__C _21753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14018_ _15435_/A _15153_/B _14018_/C _14176_/C vssd1 vssd1 vccd1 vccd1 _14020_/D
+ sky130_fd_sc_hd__nand4_4
X_19875_ _19753_/D _19753_/Y _19873_/Y _19874_/X vssd1 vssd1 vccd1 vccd1 _19877_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_156_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18826_ _18846_/B _18826_/B _18826_/C _18826_/D vssd1 vssd1 vccd1 vccd1 _18826_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_65_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18757_ _18757_/A _18757_/B _18757_/C vssd1 vssd1 vccd1 vccd1 _18758_/C sky130_fd_sc_hd__nand3_1
X_15969_ _15971_/B vssd1 vssd1 vccd1 vccd1 _15970_/B sky130_fd_sc_hd__inv_2
XANTENNA__21347__A1 _21349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17015__A2 _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17708_ _17705_/B _17590_/Y _17595_/A _17594_/B vssd1 vssd1 vccd1 vccd1 _17708_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18688_ _18688_/A _18839_/B vssd1 vssd1 vccd1 vccd1 _21367_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_148_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17639_ _18767_/B _17637_/X _17638_/X vssd1 vssd1 vccd1 vccd1 _17640_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_33_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13588__A1 _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_911 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13588__B2 _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20650_ _20650_/A _20650_/B vssd1 vssd1 vccd1 vccd1 _20651_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_86_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20419__A _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19309_ _19148_/A _19148_/C _19145_/Y vssd1 vssd1 vccd1 vccd1 _19311_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_74_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15520__B _15521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12260__A1 _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20581_ _20712_/B _20579_/X _20408_/B _20450_/X vssd1 vssd1 vccd1 vccd1 _20628_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout304_A _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21202_ _21090_/A _21206_/A _21089_/B _21086_/B _21086_/A vssd1 vssd1 vccd1 vccd1
+ _21204_/B sky130_fd_sc_hd__o32ai_4
XFILLER_0_44_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16989__D _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17447__B _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21133_ _21134_/B _21134_/A vssd1 vssd1 vccd1 vccd1 _21244_/B sky130_fd_sc_hd__and2b_1
Xfanout401 _21769_/Q vssd1 vssd1 vccd1 vccd1 _13157_/B sky130_fd_sc_hd__buf_4
Xfanout412 _21767_/Q vssd1 vssd1 vccd1 vccd1 _14698_/A sky130_fd_sc_hd__clkbuf_8
Xfanout423 _15076_/A vssd1 vssd1 vccd1 vccd1 _14557_/A sky130_fd_sc_hd__clkbuf_8
X_21064_ _21064_/A _21064_/B vssd1 vssd1 vccd1 vccd1 _21065_/B sky130_fd_sc_hd__or2_1
Xfanout434 _21762_/Q vssd1 vssd1 vccd1 vccd1 _14712_/B sky130_fd_sc_hd__buf_4
XFILLER_0_10_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout445 _12785_/B vssd1 vssd1 vccd1 vccd1 _12245_/B sky130_fd_sc_hd__buf_2
XANTENNA__20389__A2 _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout456 _14250_/B vssd1 vssd1 vccd1 vccd1 _16380_/B sky130_fd_sc_hd__clkbuf_8
X_20015_ _20125_/A _20014_/C _20014_/A vssd1 vssd1 vccd1 vccd1 _20015_/X sky130_fd_sc_hd__a21o_1
Xfanout467 _14698_/D vssd1 vssd1 vccd1 vccd1 _15001_/B sky130_fd_sc_hd__clkbuf_4
Xfanout478 _14217_/D vssd1 vssd1 vccd1 vccd1 _13913_/C sky130_fd_sc_hd__buf_4
Xfanout489 _21747_/Q vssd1 vssd1 vccd1 vccd1 _16399_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__21338__A1 _21407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21966_ _21974_/CLK _21966_/D vssd1 vssd1 vccd1 vccd1 hold282/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__16214__B1 _16418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20917_ _20917_/A _20917_/B vssd1 vssd1 vccd1 vccd1 _20918_/B sky130_fd_sc_hd__nand2_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21897_ _21932_/CLK _21897_/D vssd1 vssd1 vccd1 vccd1 hold151/A sky130_fd_sc_hd__dfxtp_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ _11650_/A _11650_/B _11650_/C vssd1 vssd1 vccd1 vccd1 _11652_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_77_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14776__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20848_ _20848_/A _20848_/B vssd1 vssd1 vccd1 vccd1 _20849_/B sky130_fd_sc_hd__nor2_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout30 _21489_/S vssd1 vssd1 vccd1 vccd1 _21442_/S sky130_fd_sc_hd__clkbuf_8
Xfanout41 _21329_/X vssd1 vssd1 vccd1 vccd1 _21421_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_36_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout52 _11121_/S vssd1 vssd1 vccd1 vccd1 _11108_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA__18444__D _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12251__A1 _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11581_ _12426_/B _12511_/A vssd1 vssd1 vccd1 vccd1 _11595_/A sky130_fd_sc_hd__nand2_1
Xfanout63 _19185_/B vssd1 vssd1 vccd1 vccd1 _21293_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21151__C _21815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20779_ _20912_/A _20780_/B vssd1 vssd1 vccd1 vccd1 _20916_/B sky130_fd_sc_hd__nor2_1
Xfanout74 _21849_/Q vssd1 vssd1 vccd1 vccd1 _19013_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12251__B2 _12242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout85 _19053_/B vssd1 vssd1 vccd1 vccd1 _19223_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13320_ _14712_/A _14712_/B _14391_/B _13913_/C vssd1 vssd1 vccd1 vccd1 _13320_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_80_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout96 _21843_/Q vssd1 vssd1 vccd1 vccd1 fanout96/X sky130_fd_sc_hd__buf_4
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18741__B _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13251_ _13252_/A _13252_/B vssd1 vssd1 vccd1 vccd1 _13251_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18555__A1_N _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12202_ _12203_/A _12203_/B _12203_/C vssd1 vssd1 vccd1 vccd1 _12202_/Y sky130_fd_sc_hd__nor3_1
X_13182_ _14712_/B _14384_/D _14391_/B _14712_/A vssd1 vssd1 vccd1 vccd1 _13183_/B
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__16899__D _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12133_ _12115_/A _12115_/C _12115_/B vssd1 vssd1 vccd1 vccd1 _12133_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17990_ _17990_/A _17990_/B vssd1 vssd1 vccd1 vccd1 _18091_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__18690__B2 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16941_ _16938_/X _16941_/B vssd1 vssd1 vccd1 vccd1 _16984_/B sky130_fd_sc_hd__and2b_1
X_12064_ _12053_/A _12053_/C _12053_/B vssd1 vssd1 vccd1 vccd1 _12066_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__21577__A1 _11061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15308__D _21735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11015_ mstream_o[89] hold62/X _11027_/S vssd1 vssd1 vccd1 vccd1 _21626_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14212__D _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19660_ _19542_/A _19541_/B _19539_/X vssd1 vssd1 vccd1 vccd1 _19660_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16872_ _16866_/A _16866_/C _16866_/B vssd1 vssd1 vccd1 vccd1 _16873_/C sky130_fd_sc_hd__a21o_1
XANTENNA__14059__A2 _14873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16453__B1 _16743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18188__B _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18611_ _18608_/Y _18609_/X _18476_/X _18516_/A vssd1 vssd1 vccd1 vccd1 _18611_/X
+ sky130_fd_sc_hd__a211o_1
X_15823_ _15823_/A _15823_/B _15823_/C vssd1 vssd1 vccd1 vccd1 _15823_/X sky130_fd_sc_hd__or3_4
X_19591_ _19589_/X _19590_/Y _19291_/A _19291_/B vssd1 vssd1 vccd1 vccd1 _19591_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__21329__A1 _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13406__A _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18542_ _18542_/A _18542_/B vssd1 vssd1 vccd1 vccd1 _18683_/A sky130_fd_sc_hd__or2_4
XTAP_3350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15754_ _15755_/A _15755_/B vssd1 vssd1 vccd1 vccd1 _15756_/A sky130_fd_sc_hd__or2_1
XFILLER_0_99_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12966_ _12966_/A _12966_/B _12966_/C vssd1 vssd1 vccd1 vccd1 _12967_/B sky130_fd_sc_hd__and3_1
XTAP_3361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14705_ _14705_/A _14705_/B _14705_/C vssd1 vssd1 vccd1 vccd1 _14707_/B sky130_fd_sc_hd__nand3_2
XTAP_3394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13019__B1 _21768_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18473_ _18473_/A _18473_/B vssd1 vssd1 vccd1 vccd1 _18475_/B sky130_fd_sc_hd__xor2_1
X_11917_ _11917_/A _11917_/B _11917_/C vssd1 vssd1 vccd1 vccd1 _11924_/A sky130_fd_sc_hd__nand3_1
X_15685_ _15520_/X _15522_/X _15683_/Y _15684_/X vssd1 vssd1 vccd1 vccd1 _15687_/B
+ sky130_fd_sc_hd__o211a_2
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ _21743_/Q _14367_/A _12897_/C _12897_/D vssd1 vssd1 vccd1 vccd1 _13032_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17424_ _17425_/A _17425_/B vssd1 vssd1 vccd1 vccd1 _17424_/X sky130_fd_sc_hd__and2_2
X_14636_ _15155_/C _15978_/B _14637_/C _14785_/A vssd1 vssd1 vccd1 vccd1 _14638_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14767__B1 _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11848_ _11848_/A _11848_/B _11848_/C vssd1 vssd1 vccd1 vccd1 _11854_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_56_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17355_ _17356_/A _17356_/B _17356_/C _17356_/D vssd1 vssd1 vccd1 vccd1 _17355_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_138_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14567_ _14568_/A _14568_/B _14568_/C vssd1 vssd1 vccd1 vccd1 _14567_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16508__A1 _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16508__B2 _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11779_ _12268_/A _12443_/A vssd1 vssd1 vccd1 vccd1 _11781_/B sky130_fd_sc_hd__and2_1
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18932__A _19092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16306_ _16306_/A _16306_/B vssd1 vssd1 vccd1 vccd1 _16308_/A sky130_fd_sc_hd__nor2_1
XANTENNA__19170__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13518_ _13518_/A _13518_/B _13518_/C _13518_/D vssd1 vssd1 vccd1 vccd1 _13518_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_82_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17286_ _17286_/A _17286_/B vssd1 vssd1 vccd1 vccd1 _17288_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14498_ _14813_/A _15653_/C _15112_/D _14659_/A vssd1 vssd1 vccd1 vccd1 _14498_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19025_ _18859_/D _18860_/B _19023_/X _19024_/Y vssd1 vssd1 vccd1 vccd1 _19174_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16237_ _16237_/A vssd1 vssd1 vccd1 vccd1 _16237_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13449_ _13449_/A _13449_/B vssd1 vssd1 vccd1 vccd1 _13451_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_113_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12980__A _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16452__A _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16168_ _16169_/A _16169_/B vssd1 vssd1 vccd1 vccd1 _16322_/B sky130_fd_sc_hd__or2_1
XFILLER_0_140_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18130__B1 _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19185__D _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11596__A _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15119_ _16196_/A _15022_/B _15120_/C _15266_/A vssd1 vssd1 vccd1 vccd1 _15122_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16602__D _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16099_ _16100_/A _16100_/B vssd1 vssd1 vccd1 vccd1 _16099_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_103_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14298__A2 _14296_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19927_ _19928_/B _19928_/A vssd1 vssd1 vccd1 vccd1 _19927_/X sky130_fd_sc_hd__and2b_1
XANTENNA__17283__A _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19858_ _19857_/B _19857_/C _19857_/A vssd1 vssd1 vccd1 vccd1 _19858_/X sky130_fd_sc_hd__a21o_1
X_18809_ _18658_/A _18658_/C _18658_/B vssd1 vssd1 vccd1 vccd1 _18810_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_78_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19789_ _19471_/X _19633_/X _19788_/C _19475_/A _19632_/Y vssd1 vssd1 vccd1 vccd1
+ _19789_/Y sky130_fd_sc_hd__o221ai_4
XANTENNA__20791__A2 _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12858__C _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21820_ _21821_/CLK _21820_/D vssd1 vssd1 vccd1 vccd1 hold294/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_92_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15234__C _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21751_ _22038_/CLK _21751_/D vssd1 vssd1 vccd1 vccd1 _21751_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__16747__A1 _21830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20543__A2 _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout254_A _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15531__A _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20702_ _20530_/Y _20532_/Y _20700_/A _20701_/Y vssd1 vssd1 vccd1 vccd1 _20705_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_148_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18545__C _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21682_ _21682_/CLK _21682_/D vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20633_ _20630_/Y _20631_/X _20496_/A _20499_/C vssd1 vssd1 vccd1 vccd1 _20633_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_135_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout421_A _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18842__A _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout519_A _21740_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20564_ _20685_/A _21264_/B _21171_/A _20564_/D vssd1 vssd1 vccd1 vccd1 _20685_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_74_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20495_ _20492_/A _20493_/Y _20299_/A _20300_/X vssd1 vssd1 vccd1 vccd1 _20496_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_131_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11339__A3 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17608__D _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold299_A hold299/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21116_ _21116_/A _21188_/A _21116_/C vssd1 vssd1 vccd1 vccd1 _21188_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_121_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19392__B _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22096_ _22096_/CLK _22096_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[32] sky130_fd_sc_hd__dfrtp_4
Xfanout220 _18789_/B vssd1 vssd1 vccd1 vccd1 _19906_/D sky130_fd_sc_hd__clkbuf_4
Xfanout231 _17670_/B vssd1 vssd1 vccd1 vccd1 _20273_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17193__A _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19823__D _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout242 _21808_/Q vssd1 vssd1 vccd1 vccd1 _21293_/A sky130_fd_sc_hd__clkbuf_4
X_21047_ _21047_/A _21161_/B vssd1 vssd1 vccd1 vccd1 _21050_/A sky130_fd_sc_hd__or2_1
Xfanout253 _18166_/A vssd1 vssd1 vccd1 vccd1 _19686_/B sky130_fd_sc_hd__buf_4
XFILLER_0_121_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout264 _19531_/A vssd1 vssd1 vccd1 vccd1 _19373_/B sky130_fd_sc_hd__buf_4
Xfanout275 _20317_/D vssd1 vssd1 vccd1 vccd1 _20026_/B sky130_fd_sc_hd__clkbuf_8
Xfanout286 _18010_/A vssd1 vssd1 vccd1 vccd1 _19487_/A sky130_fd_sc_hd__buf_4
Xfanout297 _21796_/Q vssd1 vssd1 vccd1 vccd1 _19650_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__15552__A1_N _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12820_ _12947_/B _12947_/C vssd1 vssd1 vccd1 vccd1 _12820_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_119_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ _12877_/B _12751_/B _13152_/D vssd1 vssd1 vccd1 vccd1 _12751_/X sky130_fd_sc_hd__and3_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21949_ _21949_/CLK _21949_/D vssd1 vssd1 vccd1 vccd1 hold187/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ _12318_/B _11701_/C _11701_/A vssd1 vssd1 vccd1 vccd1 _11702_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_139_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15470_ _15469_/B _15469_/C _15469_/A vssd1 vssd1 vccd1 vccd1 _15470_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_96_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12682_ _12681_/B _12681_/C _12681_/A vssd1 vssd1 vccd1 vccd1 _12684_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12784__B _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14421_ _14422_/A _14422_/B vssd1 vssd1 vccd1 vccd1 _14421_/Y sky130_fd_sc_hd__nand2b_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ _12109_/C _12619_/A _11563_/X _11564_/X _12750_/A vssd1 vssd1 vccd1 vccd1
+ _11793_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_38_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11180__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17140_ _17140_/A _17140_/B vssd1 vssd1 vccd1 vccd1 _17149_/A sky130_fd_sc_hd__nor2_1
X_14352_ _15695_/A _14354_/C _14817_/D _14508_/A vssd1 vssd1 vccd1 vccd1 _14357_/C
+ sky130_fd_sc_hd__a22o_1
X_11564_ _12229_/A _12155_/B _12528_/B vssd1 vssd1 vccd1 vccd1 _11564_/X sky130_fd_sc_hd__and3_1
XFILLER_0_52_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13303_ _13304_/A _13304_/B _13304_/C vssd1 vssd1 vccd1 vccd1 _13306_/B sky130_fd_sc_hd__a21o_2
X_17071_ _17071_/A _17071_/B _17071_/C vssd1 vssd1 vccd1 vccd1 _17101_/A sky130_fd_sc_hd__nand3_1
X_14283_ _14284_/A _14284_/B vssd1 vssd1 vccd1 vccd1 _14446_/B sky130_fd_sc_hd__and2_1
X_11495_ _11498_/A1 t1y[15] t0x[15] _11501_/B2 vssd1 vssd1 vccd1 vccd1 _11495_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_40_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16022_ _16021_/B _16021_/C _16021_/A vssd1 vssd1 vccd1 vccd1 _16143_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_33_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13234_ _13822_/B _14155_/C _14155_/D _13381_/C vssd1 vssd1 vccd1 vccd1 _13234_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_150_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17087__B _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14504__B _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13165_ _13287_/B _13164_/C _13164_/A vssd1 vssd1 vccd1 vccd1 _13166_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12116_ _12115_/A _12114_/Y _12066_/X _12085_/Y vssd1 vssd1 vccd1 vccd1 _12124_/A
+ sky130_fd_sc_hd__o211a_1
X_17973_ hold104/X _17972_/X fanout2/X vssd1 vssd1 vccd1 vccd1 hold105/A sky130_fd_sc_hd__mux2_1
X_13096_ _14294_/D _13092_/B _13089_/X vssd1 vssd1 vccd1 vccd1 _13224_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16924_ _17144_/A _17013_/C _17013_/D _17129_/B vssd1 vssd1 vccd1 vccd1 _16926_/A
+ sky130_fd_sc_hd__a22oi_2
X_12047_ _12781_/D _12214_/C vssd1 vssd1 vccd1 vccd1 _12048_/B sky130_fd_sc_hd__nand2_1
X_19712_ _19715_/B vssd1 vssd1 vccd1 vccd1 _19712_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21337__B _21337_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16855_ _16855_/A _17165_/C _16855_/C vssd1 vssd1 vccd1 vccd1 _17168_/A sky130_fd_sc_hd__nor3_2
X_19643_ _19644_/A _20838_/C _20838_/D _19487_/A vssd1 vssd1 vccd1 vccd1 _19645_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18927__A _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15806_ _15931_/A _15931_/B _16391_/B _16369_/B vssd1 vssd1 vccd1 vccd1 _15927_/A
+ sky130_fd_sc_hd__and4_1
X_19574_ _20650_/A _19866_/C _19575_/C _19575_/D vssd1 vssd1 vccd1 vccd1 _19574_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_88_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16786_ _16718_/A _16718_/C _16718_/B vssd1 vssd1 vccd1 vccd1 _16786_/X sky130_fd_sc_hd__a21o_1
X_13998_ _14306_/A _14155_/D _13999_/C _14153_/A vssd1 vssd1 vccd1 vccd1 _14000_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18525_ _18542_/B _18525_/B _18525_/C _18525_/D vssd1 vssd1 vccd1 vccd1 _18525_/Y
+ sky130_fd_sc_hd__nor4_2
X_15737_ _15737_/A _15737_/B _15737_/C vssd1 vssd1 vccd1 vccd1 _15741_/C sky130_fd_sc_hd__and3_2
XTAP_3180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12397__D _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12949_ _13091_/A _12950_/B _12950_/C vssd1 vssd1 vccd1 vccd1 _12949_/X sky130_fd_sc_hd__a21o_1
XTAP_3191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14776__A1_N _14774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16447__A _16813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17926__B1 _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20525__A2 _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19391__A2 _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18456_ _18327_/X _18330_/Y _18454_/Y _18455_/X vssd1 vssd1 vccd1 vccd1 _18456_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_47_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15668_ _15862_/B _15668_/B vssd1 vssd1 vccd1 vccd1 _15683_/A sky130_fd_sc_hd__and2_1
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_180 v2z[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_191 hold247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17407_ _17316_/X _17319_/Y _17405_/Y _17406_/X vssd1 vssd1 vccd1 vccd1 _17487_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_146_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15070__B _15070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14619_ _16084_/C _14457_/X _14460_/A _14460_/B vssd1 vssd1 vccd1 vccd1 _14620_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_145_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18387_ _18386_/A _18386_/B _18385_/A _18385_/B vssd1 vssd1 vccd1 vccd1 _18534_/A
+ sky130_fd_sc_hd__o211a_1
X_15599_ _15600_/A _15600_/B _15600_/C vssd1 vssd1 vccd1 vccd1 _15599_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_7_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17338_ _17557_/A _17557_/B _17915_/D _17924_/B vssd1 vssd1 vccd1 vccd1 _17340_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_44_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17269_ _17379_/B _17269_/B vssd1 vssd1 vccd1 vccd1 _17381_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_125_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19008_ _18857_/B _19185_/B _20721_/C _19008_/D vssd1 vssd1 vccd1 vccd1 _19194_/A
+ sky130_fd_sc_hd__and4b_1
XANTENNA__20416__B _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20280_ _20486_/B _20280_/B vssd1 vssd1 vccd1 vccd1 _20295_/A sky130_fd_sc_hd__and2_1
XFILLER_0_87_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18103__B1 _18101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12215__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19851__B1 _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15229__C _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14133__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19652__A2_N _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__21410__B1 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout371_A _21775_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17741__A _21796_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21803_ _21803_/CLK _21803_/D vssd1 vssd1 vccd1 vccd1 _21803_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_91_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout636_A _11089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21734_ _21803_/CLK _21734_/D vssd1 vssd1 vccd1 vccd1 _21734_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16507__D _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21665_ _21906_/CLK _21665_/D vssd1 vssd1 vccd1 vccd1 hold99/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12757__A2 _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20616_ _20616_/A _20616_/B _20616_/C vssd1 vssd1 vccd1 vccd1 _20616_/X sky130_fd_sc_hd__and3_1
XFILLER_0_149_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21596_ _21934_/CLK _21596_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[59] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_117_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13923__A1_N _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20547_ _20797_/A _21258_/A _21305_/A _21153_/B vssd1 vssd1 vccd1 vccd1 _20679_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_149_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18893__A1 _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14605__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17619__C _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13706__A1 _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12509__A2 _12402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11280_ _12420_/D _11279_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21771_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_43_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20478_ _20602_/A _21311_/B _20583_/A _20478_/D vssd1 vssd1 vccd1 vccd1 _20602_/B
+ sky130_fd_sc_hd__and4b_1
XANTENNA__17338__D _17924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13182__A2 _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14970_ _14970_/A _14970_/B vssd1 vssd1 vccd1 vccd1 _15056_/A sky130_fd_sc_hd__xnor2_1
X_22079_ _22096_/CLK _22079_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[15] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_22_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12142__B1 _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18948__A2 _19753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13921_ _14713_/A _14713_/B _15370_/B _15098_/B vssd1 vssd1 vccd1 vccd1 _13921_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__18246__A2_N fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16640_ _16639_/B _16639_/C _16639_/A vssd1 vssd1 vccd1 vccd1 _16642_/B sky130_fd_sc_hd__a21bo_1
X_13852_ _13973_/A _13851_/C _13851_/A vssd1 vssd1 vccd1 vccd1 _13852_/X sky130_fd_sc_hd__o21a_1
XANTENNA__17620__A2 _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15631__A1 _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15631__B2 _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12803_ _12803_/A _12803_/B _12803_/C _12803_/D vssd1 vssd1 vccd1 vccd1 _12803_/X
+ sky130_fd_sc_hd__or4_2
X_16571_ _16569_/X _16571_/B vssd1 vssd1 vccd1 vccd1 _16572_/B sky130_fd_sc_hd__and2b_1
XANTENNA__12445__A1 _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13783_ _13782_/A _13782_/B _13782_/C vssd1 vssd1 vccd1 vccd1 _13784_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12445__B2 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10995_ mstream_o[69] hold65/X _11005_/S vssd1 vssd1 vccd1 vccd1 _21606_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18310_ _18157_/A _18157_/Y _18307_/X _18308_/Y vssd1 vssd1 vccd1 vccd1 _18310_/Y
+ sky130_fd_sc_hd__o211ai_2
X_15522_ _15523_/B _15523_/A vssd1 vssd1 vccd1 vccd1 _15522_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_96_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12734_ _13860_/A _13269_/C _13269_/D _13554_/B vssd1 vssd1 vccd1 vccd1 _12734_/Y
+ sky130_fd_sc_hd__a22oi_1
X_19290_ _19445_/B _19126_/B _19445_/A vssd1 vssd1 vccd1 vccd1 _19291_/B sky130_fd_sc_hd__mux2_4
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18241_ _18241_/A _18241_/B vssd1 vssd1 vccd1 vccd1 _18394_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_32_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15453_ _15456_/D vssd1 vssd1 vccd1 vccd1 _15453_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_128_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ _12665_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _12667_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_139_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15321__D _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14404_ _14848_/A _15098_/B _14241_/X _14242_/X _14557_/D vssd1 vssd1 vccd1 vccd1
+ _14409_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_25_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18172_ _18170_/Y _18322_/A _19379_/B _18624_/A vssd1 vssd1 vccd1 vccd1 _18322_/B
+ sky130_fd_sc_hd__and4bb_1
X_11616_ _12302_/A _12858_/C _12991_/D _12312_/A vssd1 vssd1 vccd1 vccd1 _11667_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_65_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15384_ _15384_/A _15384_/B _15384_/C vssd1 vssd1 vccd1 vccd1 _15386_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_108_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12596_ _12831_/D _12596_/B vssd1 vssd1 vccd1 vccd1 _12825_/B sky130_fd_sc_hd__or2_1
XFILLER_0_154_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17123_ _17146_/A _17146_/B _17123_/C _17145_/B vssd1 vssd1 vccd1 vccd1 _17123_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_136_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14335_ _14160_/B _14162_/B _14489_/A _14334_/Y vssd1 vssd1 vccd1 vccd1 _14489_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_108_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11547_ _21725_/D _11555_/B vssd1 vssd1 vccd1 vccd1 _11547_/X sky130_fd_sc_hd__or2_2
XFILLER_0_53_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17054_ _17052_/X _17054_/B vssd1 vssd1 vccd1 vccd1 _17069_/A sky130_fd_sc_hd__and2b_1
X_14266_ _14105_/B _14105_/Y _14264_/Y _14265_/X vssd1 vssd1 vccd1 vccd1 _14268_/B
+ sky130_fd_sc_hd__o211ai_4
X_11478_ _11502_/A1 t2x[9] v1z[9] fanout20/X _11477_/X vssd1 vssd1 vccd1 vccd1 _11478_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__14234__B _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16005_ _15876_/X _15878_/Y _16003_/Y _16004_/X vssd1 vssd1 vccd1 vccd1 _16007_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_122_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13217_ _13218_/A _13218_/B _13218_/C vssd1 vssd1 vccd1 vccd1 _13217_/X sky130_fd_sc_hd__and3_1
XANTENNA__18636__A1 _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14197_ _14196_/B _14362_/B _14196_/A vssd1 vssd1 vccd1 vccd1 _14198_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_21_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11577__C _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13148_ _13148_/A _13148_/B vssd1 vssd1 vccd1 vccd1 _13166_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14250__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13079_ _12938_/B _12938_/Y _13077_/X _13078_/Y vssd1 vssd1 vccd1 vccd1 _13083_/B
+ sky130_fd_sc_hd__a211oi_2
X_17956_ _17958_/B vssd1 vssd1 vccd1 vccd1 _17956_/Y sky130_fd_sc_hd__inv_2
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14673__A2 _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16907_ _16843_/Y _16904_/X _16958_/A _16903_/A vssd1 vssd1 vccd1 vccd1 _16908_/C
+ sky130_fd_sc_hd__o211ai_2
X_17887_ _17884_/A _17885_/Y _17772_/Y _17776_/A vssd1 vssd1 vccd1 vccd1 _17887_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__11085__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19626_ _19626_/A _19626_/B vssd1 vssd1 vccd1 vccd1 _19629_/A sky130_fd_sc_hd__xnor2_1
X_16838_ _16838_/A _16838_/B vssd1 vssd1 vccd1 vccd1 _16840_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__21083__A _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16769_ _16769_/A _16849_/A vssd1 vssd1 vccd1 vccd1 _16838_/B sky130_fd_sc_hd__nor2_1
X_19557_ _19556_/B _19556_/C _19556_/A vssd1 vssd1 vccd1 vccd1 _19557_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16177__A _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18508_ _18508_/A _18508_/B _18508_/C vssd1 vssd1 vccd1 vccd1 _18511_/B sky130_fd_sc_hd__nand3_4
X_19488_ _20838_/C _19487_/X _19486_/X vssd1 vssd1 vccd1 vccd1 _19490_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__17375__A1 _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17375__B2 _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18439_ _18440_/A _18440_/B vssd1 vssd1 vccd1 vccd1 _18564_/B sky130_fd_sc_hd__or2_1
XFILLER_0_146_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_914 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21450_ hold220/X sstream_i[27] _21494_/S vssd1 vssd1 vccd1 vccd1 _21977_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_111_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20401_ _20913_/A _20401_/B vssd1 vssd1 vccd1 vccd1 _20403_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21381_ hold111/X _21381_/B vssd1 vssd1 vccd1 vccd1 _21381_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout217_A _21040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20146__B _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20332_ _20335_/D vssd1 vssd1 vccd1 vccd1 _20332_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_109_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20263_ _20157_/A _20157_/B _20155_/X vssd1 vssd1 vccd1 vccd1 _20301_/A sky130_fd_sc_hd__a21o_1
X_22002_ _22005_/CLK _22002_/D vssd1 vssd1 vccd1 vccd1 hold166/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__16638__B1 _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13983__B _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21258__A _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20194_ _20194_/A _20329_/B vssd1 vssd1 vccd1 vccd1 _20196_/B sky130_fd_sc_hd__or2_1
XANTENNA_fanout586_A _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19951__A _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19052__A1 _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12675__A1 _12785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12675__B2 _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17621__D _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10989__A1 _10988_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21717_ _21934_/CLK hold2/X fanout641/X vssd1 vssd1 vccd1 vccd1 _21717_/Q sky130_fd_sc_hd__dfrtp_4
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16815__A _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19107__A2 _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12450_ _12451_/A _12451_/B vssd1 vssd1 vccd1 vccd1 _12544_/B sky130_fd_sc_hd__nand2_1
X_21648_ _21722_/CLK _21648_/D fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[111]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11401_ _11400_/X _17334_/B _11401_/S vssd1 vssd1 vccd1 vccd1 _21805_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_152_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15129__B1 _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12381_ _11802_/X _11805_/X _12379_/Y _12380_/X vssd1 vssd1 vccd1 vccd1 _12381_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_62_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_80 hold234/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21579_ mstream_o[42] _11066_/Y _21579_/S vssd1 vssd1 vccd1 vccd1 _22106_/D sky130_fd_sc_hd__mux2_1
XANTENNA_91 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14120_ _14280_/B _14118_/Y _13956_/B _13958_/A vssd1 vssd1 vccd1 vccd1 _14121_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__12781__C _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20673__A1 _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11332_ _15174_/D _11331_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21784_/D sky130_fd_sc_hd__mux2_1
XANTENNA__20673__B2 _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13596__D _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14352__A1 _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14051_ _14051_/A _14051_/B vssd1 vssd1 vccd1 vccd1 _14070_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14352__B2 _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11263_ fanout59/X v0z[9] fanout19/X _11262_/X vssd1 vssd1 vccd1 vccd1 _11263_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13002_ _13002_/A _13002_/B _13002_/C vssd1 vssd1 vccd1 vccd1 _13003_/A sky130_fd_sc_hd__and3_1
XFILLER_0_31_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13893__B _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11194_ hold116/X fanout22/X _11193_/X vssd1 vssd1 vccd1 vccd1 _11194_/X sky130_fd_sc_hd__a21o_1
XANTENNA__10913__A1 _10912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11694__A _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17810_ _17810_/A _17810_/B _17810_/C vssd1 vssd1 vccd1 vccd1 _17810_/X sky130_fd_sc_hd__or3_2
XFILLER_0_100_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18790_ _18790_/A _18790_/B _18947_/B vssd1 vssd1 vccd1 vccd1 _18790_/X sky130_fd_sc_hd__and3_1
XFILLER_0_100_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17741_ _21796_/Q _17741_/B _17870_/A _17741_/D vssd1 vssd1 vccd1 vccd1 _17870_/B
+ sky130_fd_sc_hd__nand4_2
X_14953_ _14952_/B _15169_/B _14952_/A vssd1 vssd1 vccd1 vccd1 _14954_/C sky130_fd_sc_hd__a21o_1
XANTENNA__20800__A _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12302__B _12402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13904_ _13904_/A _14051_/A _13904_/C vssd1 vssd1 vccd1 vccd1 _14051_/B sky130_fd_sc_hd__nand3_1
X_17672_ _19123_/B _20270_/C _18789_/B _19123_/A vssd1 vssd1 vccd1 vccd1 _17673_/C
+ sky130_fd_sc_hd__a22o_1
X_14884_ _14883_/B _14883_/C _14883_/A vssd1 vssd1 vccd1 vccd1 _14884_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__14407__A2 _15091_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18196__B _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16623_ _16622_/B _16622_/C _16622_/A vssd1 vssd1 vccd1 vccd1 _16625_/B sky130_fd_sc_hd__a21bo_1
X_19411_ _20103_/A _19546_/D vssd1 vssd1 vccd1 vccd1 _19412_/B sky130_fd_sc_hd__nand2_1
X_13835_ _13835_/A _13835_/B vssd1 vssd1 vccd1 vccd1 _13844_/A sky130_fd_sc_hd__or2_1
XANTENNA__21088__A2_N _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16554_ _21825_/Q _16734_/B _17433_/A _17526_/B vssd1 vssd1 vccd1 vccd1 _16554_/X
+ sky130_fd_sc_hd__and4_1
X_19342_ _19189_/A _19188_/A _19188_/B _19184_/B _19184_/A vssd1 vssd1 vccd1 vccd1
+ _19343_/B sky130_fd_sc_hd__o32ai_4
X_13766_ _14859_/A _14218_/B _13766_/C _13910_/A vssd1 vssd1 vccd1 vccd1 _13910_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_84_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10978_ _10978_/A _10978_/B vssd1 vssd1 vccd1 vccd1 _10978_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_134_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15505_ _15380_/A _15380_/B _15378_/Y vssd1 vssd1 vccd1 vccd1 _15523_/A sky130_fd_sc_hd__o21bai_4
XFILLER_0_84_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19273_ _19099_/B _19101_/B _19270_/X _19272_/Y vssd1 vssd1 vccd1 vccd1 _19275_/A
+ sky130_fd_sc_hd__a211o_1
X_12717_ _12942_/A _12717_/B vssd1 vssd1 vccd1 vccd1 _12813_/A sky130_fd_sc_hd__or2_1
XFILLER_0_85_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16485_ _16485_/A _16485_/B vssd1 vssd1 vccd1 vccd1 _16771_/A sky130_fd_sc_hd__xor2_1
X_13697_ _13698_/A _13698_/B _13698_/C vssd1 vssd1 vccd1 vccd1 _13697_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16725__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18224_ _18225_/A _18225_/B _18225_/C vssd1 vssd1 vccd1 vccd1 _18224_/Y sky130_fd_sc_hd__nor3_2
X_15436_ _15436_/A _15577_/B vssd1 vssd1 vccd1 vccd1 _15438_/A sky130_fd_sc_hd__or2_2
XFILLER_0_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12648_ _12649_/A _12649_/B vssd1 vssd1 vccd1 vccd1 _12648_/X sky130_fd_sc_hd__and2_2
XANTENNA__20247__A _21831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18155_ _18304_/B _18155_/B _18155_/C vssd1 vssd1 vccd1 vccd1 _18157_/A sky130_fd_sc_hd__and3_2
X_15367_ _15632_/B _15510_/B _15368_/D _15892_/A vssd1 vssd1 vccd1 vccd1 _15370_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12579_ _12578_/B _12578_/C _12578_/A vssd1 vssd1 vccd1 vccd1 _12579_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_142_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17106_ _17106_/A _17106_/B _17106_/C vssd1 vssd1 vccd1 vccd1 _17120_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_29_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14318_ _14317_/A _14317_/B _14317_/C vssd1 vssd1 vccd1 vccd1 _14319_/B sky130_fd_sc_hd__o21a_1
X_18086_ _18107_/B _18087_/B _18087_/C _18087_/D vssd1 vssd1 vccd1 vccd1 _18086_/Y
+ sky130_fd_sc_hd__nor4_2
Xhold306 hold306/A vssd1 vssd1 vccd1 vccd1 hold306/X sky130_fd_sc_hd__buf_4
X_15298_ _15298_/A _15298_/B vssd1 vssd1 vccd1 vccd1 _15336_/A sky130_fd_sc_hd__nand2_2
Xhold317 hold317/A vssd1 vssd1 vccd1 vccd1 hold317/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold328 hold328/A vssd1 vssd1 vccd1 vccd1 hold328/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17037_ _17028_/A _17028_/B _17028_/C vssd1 vssd1 vccd1 vccd1 _17038_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14249_ _14248_/A _21759_/Q hold313/A vssd1 vssd1 vccd1 vccd1 _14251_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_123_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17556__A _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10904__A1 _10903_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15076__A _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16610__D _17334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18988_ _18987_/A _18987_/B _18985_/Y _18986_/X vssd1 vssd1 vccd1 vccd1 _18988_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17939_ _17799_/A _17799_/C _17799_/B vssd1 vssd1 vccd1 vccd1 _17940_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20950_ _20951_/A _20951_/B _20951_/C vssd1 vssd1 vccd1 vccd1 _20952_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_96_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16619__B _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19609_ _19609_/A _19609_/B vssd1 vssd1 vccd1 vccd1 _19612_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_95_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20881_ _20881_/A _20881_/B vssd1 vssd1 vccd1 vccd1 _20883_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout167_A _19732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13324__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11093__A0 _11051_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13043__B _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout334_A _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_700 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21502_ hold269/X sstream_i[79] _21507_/S vssd1 vssd1 vccd1 vccd1 _22029_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_9_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12882__B _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11779__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18848__A1 _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21433_ hold278/X sstream_i[10] _21442_/S vssd1 vssd1 vccd1 vccd1 _21960_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_12_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18848__B2 _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14155__A _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11396__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21364_ _21412_/A _21364_/B vssd1 vssd1 vccd1 vccd1 _21364_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20315_ _20316_/A _20316_/B vssd1 vssd1 vccd1 vccd1 _20466_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_43_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21295_ _21295_/A _21295_/B vssd1 vssd1 vccd1 vccd1 _21297_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20246_ _21832_/Q _20247_/C _20247_/D _21831_/Q vssd1 vssd1 vccd1 vccd1 _20248_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_101_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17284__B1 _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20177_ _20177_/A _20177_/B vssd1 vssd1 vccd1 vccd1 _20181_/A sky130_fd_sc_hd__xor2_2
XANTENNA__12403__A _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11950_ _11953_/A vssd1 vssd1 vccd1 vccd1 _11952_/C sky130_fd_sc_hd__inv_2
XTAP_3735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11320__A1 _11319_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16529__B _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10901_ _10902_/B _10902_/C _10902_/A vssd1 vssd1 vccd1 vccd1 _10911_/B sky130_fd_sc_hd__a21oi_1
XTAP_3768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11881_ _11881_/A _11881_/B vssd1 vssd1 vccd1 vccd1 _11958_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_93_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13620_ _14713_/A _14713_/B _14077_/B _14234_/C vssd1 vssd1 vccd1 vccd1 _13620_/X
+ sky130_fd_sc_hd__and4_1
X_10832_ _11047_/B _11048_/A _11047_/A vssd1 vssd1 vccd1 vccd1 _11051_/A sky130_fd_sc_hd__o21ba_2
XANTENNA__17339__A1 _17557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17339__B2 _17557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11084__A0 _10965_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13551_ _13392_/Y _13395_/X _13548_/A _13549_/X vssd1 vssd1 vccd1 vccd1 _13551_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12502_ _14133_/D _13258_/C _13258_/D _13983_/B vssd1 vssd1 vccd1 vccd1 _12503_/B
+ sky130_fd_sc_hd__a22o_1
X_16270_ _16371_/A _16369_/B _21755_/Q _16380_/A vssd1 vssd1 vccd1 vccd1 _16270_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20990__A1_N _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14022__B1 _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ _13332_/A _13332_/C _13332_/B vssd1 vssd1 vccd1 vccd1 _13483_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_81_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16562__A2 _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15221_ _15221_/A _15362_/A vssd1 vssd1 vccd1 vccd1 _15222_/B sky130_fd_sc_hd__xor2_2
X_12433_ _12433_/A _12433_/B vssd1 vssd1 vccd1 vccd1 _12435_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_63_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15152_ _15579_/D _15829_/C _15954_/D _15153_/B vssd1 vssd1 vccd1 vccd1 _15152_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12364_ _12364_/A _12364_/B _12364_/C vssd1 vssd1 vccd1 vccd1 _12367_/A sky130_fd_sc_hd__nand3_2
XANTENNA__19575__B _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14103_ _13939_/B _13939_/Y _14100_/X _14102_/Y vssd1 vssd1 vccd1 vccd1 _14105_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_121_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14325__A1 _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11315_ fanout58/X v0z[22] fanout17/X _11314_/X vssd1 vssd1 vccd1 vccd1 _11315_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15083_ _15082_/B _15082_/C _15082_/A vssd1 vssd1 vccd1 vccd1 _15085_/D sky130_fd_sc_hd__a21oi_1
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14325__B2 _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19960_ _19961_/A _20381_/A _19961_/C _19961_/D vssd1 vssd1 vccd1 vccd1 _19963_/A
+ sky130_fd_sc_hd__o22ai_1
X_12295_ _12289_/A _12289_/B _12294_/X vssd1 vssd1 vccd1 vccd1 _12391_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_121_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14034_ _14365_/A _14537_/A _14516_/A _21742_/Q vssd1 vssd1 vccd1 vccd1 _14037_/C
+ sky130_fd_sc_hd__a22o_1
X_18911_ _19686_/A _19238_/C _18911_/C _19065_/A vssd1 vssd1 vccd1 vccd1 _19065_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_120_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11246_ _11549_/A t1x[5] v2z[5] _21724_/D _11245_/X vssd1 vssd1 vccd1 vccd1 _11246_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__17095__B _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19891_ _19891_/A _19891_/B vssd1 vssd1 vccd1 vccd1 _19893_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17526__D _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18842_ _20770_/B _18842_/B vssd1 vssd1 vccd1 vccd1 _18842_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11177_ _13155_/A _11176_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21742_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15985_ _15986_/A _15986_/B _15986_/C vssd1 vssd1 vccd1 vccd1 _15985_/X sky130_fd_sc_hd__a21o_1
X_18773_ _20650_/A _18773_/B vssd1 vssd1 vccd1 vccd1 _18775_/C sky130_fd_sc_hd__and2_1
XFILLER_0_98_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14936_ _14774_/D _15838_/B _16314_/D _14936_/D vssd1 vssd1 vccd1 vccd1 _14939_/A
+ sky130_fd_sc_hd__and4b_1
X_17724_ _18703_/A _19053_/B _17720_/X _17722_/Y vssd1 vssd1 vccd1 vccd1 _17725_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_136_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21374__A2 _14126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15589__B1 _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14867_ _14868_/A _14868_/B _14868_/C vssd1 vssd1 vccd1 vccd1 _14887_/A sky130_fd_sc_hd__a21oi_2
X_17655_ _17651_/X _17652_/Y _17531_/X _17533_/X vssd1 vssd1 vccd1 vccd1 _17689_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_89_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13818_ _13806_/X _13818_/B vssd1 vssd1 vccd1 vccd1 _13960_/A sky130_fd_sc_hd__and2b_1
X_16606_ _17557_/A _17915_/A _17557_/B _17657_/A vssd1 vssd1 vccd1 vccd1 _16608_/B
+ sky130_fd_sc_hd__nand4_1
X_17586_ _17586_/A _17586_/B vssd1 vssd1 vccd1 vccd1 _17589_/A sky130_fd_sc_hd__nor2_2
X_14798_ _14795_/X _14796_/Y _14640_/B _14642_/B vssd1 vssd1 vccd1 vccd1 _14799_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_9_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11075__A0 _10903_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19325_ hold252/X _19324_/Y fanout3/X vssd1 vssd1 vccd1 vccd1 hold253/A sky130_fd_sc_hd__mux2_1
XANTENNA__21361__A _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16537_ _16537_/A _16537_/B vssd1 vssd1 vccd1 vccd1 _16680_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13749_ _15763_/A _14365_/D _13750_/C _13750_/D vssd1 vssd1 vccd1 vccd1 _13751_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21080__B _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16468_ _16468_/A _16468_/B vssd1 vssd1 vccd1 vccd1 _16476_/A sky130_fd_sc_hd__xor2_1
X_19256_ _20101_/B _19703_/C _18640_/B _20101_/A vssd1 vssd1 vccd1 vccd1 _19258_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_155_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16696__A1_N _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15419_ _15419_/A _15419_/B _15419_/C vssd1 vssd1 vccd1 vccd1 _15420_/C sky130_fd_sc_hd__nand3_1
XANTENNA__14564__A1 _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18207_ _18207_/A _18207_/B _18207_/C vssd1 vssd1 vccd1 vccd1 _18209_/B sky130_fd_sc_hd__nand3_1
XANTENNA__14564__B2 _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19187_ _19185_/D _19185_/B _21261_/B _17854_/B vssd1 vssd1 vccd1 vccd1 _19188_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16399_ _16399_/A _16399_/B vssd1 vssd1 vccd1 vccd1 _16400_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_115_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18138_ _18873_/A _19382_/B _18288_/A _18137_/D vssd1 vssd1 vccd1 vccd1 _18140_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold103 hold103/A vssd1 vssd1 vccd1 vccd1 hold103/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold114 hold114/A vssd1 vssd1 vccd1 vccd1 hold114/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18069_ _18069_/A _18069_/B _18069_/C vssd1 vssd1 vccd1 vccd1 _18071_/B sky130_fd_sc_hd__nand3_1
Xhold125 hold125/A vssd1 vssd1 vccd1 vccd1 hold125/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 hold136/A vssd1 vssd1 vccd1 vccd1 hold136/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold147 hold147/A vssd1 vssd1 vccd1 vccd1 hold147/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 hold158/A vssd1 vssd1 vccd1 vccd1 hold158/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12327__B1 _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20100_ _20101_/B _21816_/Q _20242_/C _20101_/A vssd1 vssd1 vccd1 vccd1 _20103_/C
+ sky130_fd_sc_hd__a22o_1
Xhold169 hold169/A vssd1 vssd1 vccd1 vccd1 hold169/X sky130_fd_sc_hd__dlygate4sd3_1
X_21080_ _21293_/A _21291_/A _21286_/B _21296_/B vssd1 vssd1 vccd1 vccd1 _21194_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_42_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12878__B2 _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout605 _11459_/B2 vssd1 vssd1 vccd1 vccd1 _11543_/B2 sky130_fd_sc_hd__buf_2
XFILLER_0_95_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout616 _21717_/Q vssd1 vssd1 vccd1 vccd1 _21568_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20031_ _20029_/X _20031_/B vssd1 vssd1 vccd1 vccd1 _20036_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__13319__A _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout627 _21087_/D vssd1 vssd1 vccd1 vccd1 _19535_/B sky130_fd_sc_hd__buf_2
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout638 fanout639/X vssd1 vssd1 vccd1 vccd1 _11089_/A sky130_fd_sc_hd__buf_4
XANTENNA__15718__A2_N _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12223__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout284_A _21798_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20797__D _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11302__A1 _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21982_ _22016_/CLK _21982_/D vssd1 vssd1 vccd1 vccd1 hold160/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__21365__A2 _18537_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18766__B1 _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12877__B _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20933_ _20932_/A _21048_/B _20931_/X vssd1 vssd1 vccd1 vccd1 _20934_/B sky130_fd_sc_hd__o21bai_1
XANTENNA_fanout451_A _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout549_A _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15275__A1_N _15933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20864_ _20864_/A _20985_/B vssd1 vssd1 vccd1 vccd1 _20866_/B sky130_fd_sc_hd__or2_1
XFILLER_0_7_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20795_ _20795_/A _20986_/B vssd1 vssd1 vccd1 vccd1 _20806_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19379__C _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19730__A2 _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14555__A1 _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12566__B1 _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21416_ _21412_/A _21142_/B fanout40/X vssd1 vssd1 vccd1 vccd1 _21416_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11659__D _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14307__A1 _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16812__B _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14035__D _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21347_ _21349_/A _17599_/B _21381_/B vssd1 vssd1 vccd1 vccd1 _21347_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11100_ _11066_/Y hold82/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21694_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18049__A2 _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _12080_/A _12083_/B _12073_/A vssd1 vssd1 vccd1 vccd1 _12080_/X sky130_fd_sc_hd__or3b_1
X_21278_ _21278_/A _21278_/B vssd1 vssd1 vccd1 vccd1 _21279_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_130_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11031_ mstream_o[105] hold270/X _11039_/S vssd1 vssd1 vccd1 vccd1 _21642_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_120_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20229_ _20770_/B _21396_/B vssd1 vssd1 vccd1 vccd1 _20229_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17924__A _18058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_18_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21722_/CLK sky130_fd_sc_hd__clkbuf_16
X_15770_ _15770_/A _16034_/A vssd1 vssd1 vccd1 vccd1 _16029_/A sky130_fd_sc_hd__or2_2
XTAP_3510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12982_ _12980_/X _12982_/B vssd1 vssd1 vccd1 vccd1 _12983_/B sky130_fd_sc_hd__and2b_1
XTAP_3521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21356__A2 _18101_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14721_ _14717_/X _14719_/Y _14571_/A _14974_/A vssd1 vssd1 vccd1 vccd1 _14721_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_99_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11933_ _11930_/X _11933_/B vssd1 vssd1 vccd1 vccd1 _12001_/B sky130_fd_sc_hd__and2b_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11183__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17440_ _17441_/A _17441_/B vssd1 vssd1 vccd1 vccd1 _17536_/B sky130_fd_sc_hd__nand2_2
XTAP_3598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14652_ _14652_/A _14652_/B vssd1 vssd1 vccd1 vccd1 _14654_/B sky130_fd_sc_hd__xnor2_4
XTAP_2864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11864_ _12781_/D _12528_/B _11851_/X _11556_/X _12637_/B vssd1 vssd1 vccd1 vccd1
+ _11867_/A sky130_fd_sc_hd__a32o_1
XTAP_2875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13603_ _13605_/A _13605_/B _13605_/C vssd1 vssd1 vccd1 vccd1 _13603_/X sky130_fd_sc_hd__o21a_1
XANTENNA__13899__A _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10815_ _10815_/A _10815_/B vssd1 vssd1 vccd1 vccd1 _11057_/A sky130_fd_sc_hd__nand2_2
X_17371_ _17479_/B _17371_/B vssd1 vssd1 vccd1 vccd1 _17381_/C sky130_fd_sc_hd__xnor2_4
XFILLER_0_156_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14583_ _14583_/A _14583_/B vssd1 vssd1 vccd1 vccd1 _14584_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_89_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11795_ _11795_/A _11795_/B _11795_/C vssd1 vssd1 vccd1 vccd1 _11795_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_68_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16322_ _16322_/A _16322_/B vssd1 vssd1 vccd1 vccd1 _16335_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_94_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19110_ _19432_/A _19866_/C _19111_/C _19276_/A vssd1 vssd1 vccd1 vccd1 _19112_/B
+ sky130_fd_sc_hd__a22o_1
X_13534_ _13534_/A _13534_/B vssd1 vssd1 vccd1 vccd1 _13536_/B sky130_fd_sc_hd__and2_1
XFILLER_0_125_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19041_ _18878_/X _18881_/A _19211_/B _19040_/Y vssd1 vssd1 vccd1 vccd1 _19176_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16253_ _16253_/A _16253_/B vssd1 vssd1 vccd1 vccd1 _16256_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13465_ _13466_/A _13466_/B vssd1 vssd1 vccd1 vccd1 _13605_/B sky130_fd_sc_hd__and2_1
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15204_ _15204_/A _15204_/B vssd1 vssd1 vccd1 vccd1 _15492_/A sky130_fd_sc_hd__or2_2
X_12416_ _12416_/A _12416_/B _12416_/C vssd1 vssd1 vccd1 vccd1 _12416_/Y sky130_fd_sc_hd__nand3_1
X_16184_ _16185_/A _16185_/B vssd1 vssd1 vccd1 vccd1 _16184_/X sky130_fd_sc_hd__and2_1
XANTENNA__13130__C _13269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13396_ _13396_/A _13396_/B vssd1 vssd1 vccd1 vccd1 _13398_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15135_ _15135_/A _15282_/A _15135_/C vssd1 vssd1 vccd1 vccd1 _15282_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12347_ _12348_/A _12348_/B vssd1 vssd1 vccd1 vccd1 _12437_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__20244__B _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16441__C _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15066_ _15067_/A _15067_/B _15067_/C vssd1 vssd1 vccd1 vccd1 _15068_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19237__A1 _19692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19943_ _19943_/A _19943_/B vssd1 vssd1 vccd1 vccd1 _20081_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12278_ _12238_/B _12238_/C _12238_/A vssd1 vssd1 vccd1 vccd1 _12278_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__19237__B2 _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14242__B _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14017_ _15435_/A _14018_/C _13858_/C _15153_/B vssd1 vssd1 vccd1 vccd1 _14020_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16160__D _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17834__A _19636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _11122_/A t2y[1] t0y[1] _11123_/A vssd1 vssd1 vccd1 vccd1 _11229_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19874_ _20650_/A _19874_/B _19874_/C _19874_/D vssd1 vssd1 vccd1 vccd1 _19874_/X
+ sky130_fd_sc_hd__and4_2
XANTENNA__11532__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18825_ _18822_/X _18823_/Y _18674_/C _18673_/Y vssd1 vssd1 vccd1 vccd1 _18826_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_65_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18756_ _18757_/A _18757_/B _18757_/C vssd1 vssd1 vccd1 vccd1 _18758_/B sky130_fd_sc_hd__a21o_1
X_15968_ _15968_/A _15968_/B vssd1 vssd1 vccd1 vccd1 _15971_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18748__B1 _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21347__A2 _17599_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11296__A0 _12402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17707_ _17830_/B _17707_/B vssd1 vssd1 vccd1 vccd1 _17837_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_72_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14919_ _21720_/Q hold174/A _10912_/X fanout5/X vssd1 vssd1 vccd1 vccd1 _14919_/X
+ sky130_fd_sc_hd__a22o_1
X_15899_ _16034_/B _15899_/B vssd1 vssd1 vccd1 vccd1 _15901_/B sky130_fd_sc_hd__nor2_1
X_18687_ _18687_/A _18687_/B vssd1 vssd1 vccd1 vccd1 _18839_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_37_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13037__A1 _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17638_ _18008_/A _18767_/B _18616_/D _18008_/B vssd1 vssd1 vccd1 vccd1 _17638_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13588__A2 _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17569_ _17570_/A _17570_/B _17570_/C vssd1 vssd1 vccd1 vccd1 _17569_/X sky130_fd_sc_hd__and3_1
XFILLER_0_74_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19199__C _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20419__B _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19308_ _19308_/A _19308_/B vssd1 vssd1 vccd1 vccd1 _19311_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_58_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20580_ _20408_/B _20450_/X _20712_/B _20579_/X vssd1 vssd1 vccd1 vccd1 _20628_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_116_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12260__A2 _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19239_ _19535_/B _20148_/C _19240_/C _19387_/A vssd1 vssd1 vccd1 vccd1 _19241_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11122__A _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21201_ _21201_/A _21201_/B vssd1 vssd1 vccd1 vccd1 _21204_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13975__C _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21132_ _20981_/A _20981_/B _20984_/A vssd1 vssd1 vccd1 vccd1 _21134_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__19228__A1 _19230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout402 _15763_/A vssd1 vssd1 vccd1 vccd1 _15375_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout499_A _21744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11268__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17239__B1 _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13049__A _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21063_ _21064_/A _21064_/B vssd1 vssd1 vccd1 vccd1 _21065_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout413 _12899_/B vssd1 vssd1 vccd1 vccd1 _12109_/C sky130_fd_sc_hd__buf_4
Xfanout424 _12771_/C vssd1 vssd1 vccd1 vccd1 _15076_/A sky130_fd_sc_hd__buf_6
Xfanout435 _12267_/A vssd1 vssd1 vccd1 vccd1 _12094_/A sky130_fd_sc_hd__buf_4
XANTENNA__11523__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout446 _21759_/Q vssd1 vssd1 vccd1 vccd1 _12785_/B sky130_fd_sc_hd__clkbuf_4
X_20014_ _20014_/A _20125_/A _20014_/C vssd1 vssd1 vccd1 vccd1 _20125_/B sky130_fd_sc_hd__nand3_1
Xfanout457 hold320/X vssd1 vssd1 vccd1 vccd1 _14250_/B sky130_fd_sc_hd__clkbuf_4
Xfanout468 _14698_/D vssd1 vssd1 vccd1 vccd1 _16414_/B sky130_fd_sc_hd__buf_4
XANTENNA__20170__A _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout479 _14217_/D vssd1 vssd1 vccd1 vccd1 _16418_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__15264__A _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21338__A2 _12493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11287__B1 _11286_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18203__A2 _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21965_ _21974_/CLK _21965_/D vssd1 vssd1 vccd1 vccd1 hold265/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__20546__B1 _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16214__A1 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16214__B2 _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20916_ _20916_/A _20916_/B _21033_/A vssd1 vssd1 vccd1 vccd1 _20917_/B sky130_fd_sc_hd__or3_1
XFILLER_0_16_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21896_ _21932_/CLK hold35/X vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__dfxtp_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14776__B2 _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20847_ _20845_/D _21293_/B _10798_/Y _20721_/D vssd1 vssd1 vccd1 vccd1 _20848_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xfanout20 _11224_/Y vssd1 vssd1 vccd1 vccd1 fanout20/X sky130_fd_sc_hd__clkbuf_8
Xfanout31 _21490_/S vssd1 vssd1 vccd1 vccd1 _21489_/S sky130_fd_sc_hd__clkbuf_8
Xfanout42 _21329_/X vssd1 vssd1 vccd1 vccd1 _21403_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout53 _11112_/S vssd1 vssd1 vccd1 vccd1 _11121_/S sky130_fd_sc_hd__clkbuf_8
X_11580_ _12020_/A _12326_/D _14621_/D _12403_/A vssd1 vssd1 vccd1 vccd1 _11580_/X
+ sky130_fd_sc_hd__and4_1
X_20778_ _20911_/A _20778_/B vssd1 vssd1 vccd1 vccd1 _20780_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12251__A2 _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout64 _19185_/B vssd1 vssd1 vccd1 vccd1 _20178_/B sky130_fd_sc_hd__buf_2
XFILLER_0_64_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout75 _21848_/Q vssd1 vssd1 vccd1 vccd1 _19201_/B sky130_fd_sc_hd__buf_4
XFILLER_0_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20048__C _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout86 _20671_/B vssd1 vssd1 vccd1 vccd1 _21264_/A sky130_fd_sc_hd__buf_4
XFILLER_0_92_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout9_A fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout97 _21843_/Q vssd1 vssd1 vccd1 vccd1 _21151_/A sky130_fd_sc_hd__buf_6
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13250_ _13244_/B _13250_/B _13250_/C vssd1 vssd1 vccd1 vccd1 _13252_/B sky130_fd_sc_hd__and3b_1
XFILLER_0_150_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12201_ _12195_/A _12195_/B _12195_/C vssd1 vssd1 vccd1 vccd1 _12203_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_150_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13181_ _14712_/A _14712_/B _14384_/D _14391_/B vssd1 vssd1 vccd1 vccd1 _13183_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_60_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12132_ _12124_/A _12124_/C _12124_/B vssd1 vssd1 vccd1 vccd1 _12132_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_103_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18690__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14700__A1 _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16940_ _17029_/A _17124_/C _17145_/B _17029_/B vssd1 vssd1 vccd1 vccd1 _16941_/B
+ sky130_fd_sc_hd__a22o_1
X_12063_ _12063_/A _12063_/B vssd1 vssd1 vccd1 vccd1 _12066_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11514__A1 _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11514__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ mstream_o[88] hold71/X _11027_/S vssd1 vssd1 vccd1 vccd1 _21625_/D sky130_fd_sc_hd__mux2_1
X_16871_ _16871_/A _16871_/B vssd1 vssd1 vccd1 vccd1 _16873_/B sky130_fd_sc_hd__xor2_2
XANTENNA__16453__A1 _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18610_ _18476_/X _18516_/A _18608_/Y _18609_/X vssd1 vssd1 vccd1 vccd1 _18610_/Y
+ sky130_fd_sc_hd__o211ai_4
X_15822_ _15819_/Y _15820_/X _15683_/B _15683_/Y vssd1 vssd1 vccd1 vccd1 _15823_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16453__B2 _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18188__C _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19590_ _19723_/A _21171_/B _19723_/B _19723_/C vssd1 vssd1 vccd1 vccd1 _19590_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_56_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21329__A2 _11549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15753_ _15753_/A _15753_/B vssd1 vssd1 vccd1 vccd1 _15755_/B sky130_fd_sc_hd__nor2_1
X_18541_ _18537_/A _18536_/B _18534_/Y vssd1 vssd1 vccd1 vccd1 _18688_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_35_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13406__B _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12965_ _12966_/A _12966_/B _12966_/C vssd1 vssd1 vccd1 vccd1 _13250_/B sky130_fd_sc_hd__a21oi_1
XTAP_3351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14704_ _14700_/X _14702_/Y _14541_/Y _14543_/X vssd1 vssd1 vccd1 vccd1 _14705_/C
+ sky130_fd_sc_hd__a211o_1
X_11916_ _11845_/A _11845_/C _11845_/B vssd1 vssd1 vccd1 vccd1 _11917_/C sky130_fd_sc_hd__a21o_1
X_15684_ _15683_/B _15683_/C _15683_/A vssd1 vssd1 vccd1 vccd1 _15684_/X sky130_fd_sc_hd__a21o_1
XTAP_3384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13019__A1 _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18472_ _18473_/A _18473_/B vssd1 vssd1 vccd1 vccd1 _18472_/Y sky130_fd_sc_hd__nand2b_1
XTAP_3395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_340 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14216__B1 _14217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13019__B2 _13018_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12896_ _12896_/A _12896_/B vssd1 vssd1 vccd1 vccd1 _12904_/A sky130_fd_sc_hd__nand2_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14635_ _15579_/D _15153_/B _15717_/C _14635_/D vssd1 vssd1 vccd1 vccd1 _14785_/A
+ sky130_fd_sc_hd__nand4_2
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14767__A1 _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17423_ _17423_/A _17423_/B vssd1 vssd1 vccd1 vccd1 _17425_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14767__B2 _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11847_ _11810_/A _11810_/C _11810_/B vssd1 vssd1 vccd1 vccd1 _11848_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_129_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14518__A _21743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14566_ _14716_/A _15234_/C vssd1 vssd1 vccd1 vccd1 _14568_/C sky130_fd_sc_hd__and2_1
XFILLER_0_83_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17354_ _17350_/X _17352_/Y _17251_/B _17251_/Y vssd1 vssd1 vccd1 vccd1 _17356_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16508__A2 _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11778_ _12261_/A _12357_/C _13017_/A _12444_/B vssd1 vssd1 vccd1 vccd1 _11781_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18932__B _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16305_ _16404_/A _16305_/B _16399_/B _16409_/B vssd1 vssd1 vccd1 vccd1 _16306_/B
+ sky130_fd_sc_hd__and4_1
X_13517_ _13518_/C _13518_/D vssd1 vssd1 vccd1 vccd1 _13517_/Y sky130_fd_sc_hd__nor2_1
X_17285_ _17283_/X _17285_/B vssd1 vssd1 vccd1 vccd1 _17286_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_67_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14497_ _14373_/A _14373_/B _14373_/C _14375_/X vssd1 vssd1 vccd1 vccd1 _14531_/A
+ sky130_fd_sc_hd__a31o_2
XANTENNA__12038__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16236_ _16302_/B _16233_/X _16075_/A _16077_/X vssd1 vssd1 vccd1 vccd1 _16237_/A
+ sky130_fd_sc_hd__o211a_1
X_19024_ _19024_/A _19024_/B _19024_/C vssd1 vssd1 vccd1 vccd1 _19024_/Y sky130_fd_sc_hd__nand3_1
X_13448_ _13449_/A _13449_/B vssd1 vssd1 vccd1 vccd1 _13448_/X sky130_fd_sc_hd__and2_1
XFILLER_0_24_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12980__B _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16452__B _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16167_ _16167_/A _16167_/B vssd1 vssd1 vccd1 vccd1 _16169_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_24_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13379_ _13682_/C _13822_/B _14155_/C _14155_/D vssd1 vssd1 vccd1 vccd1 _13527_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18130__A1 _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18130__B2 _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15118_ _15791_/A _16196_/B _16371_/A _16305_/B vssd1 vssd1 vccd1 vccd1 _15266_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11596__B _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16098_ _16098_/A _16098_/B vssd1 vssd1 vccd1 vccd1 _16100_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15049_ _15046_/Y _15047_/X _14837_/Y _14839_/X vssd1 vssd1 vccd1 vccd1 _15050_/D
+ sky130_fd_sc_hd__a211o_1
X_19926_ _19769_/A _19769_/B _19767_/X vssd1 vssd1 vccd1 vccd1 _19928_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_76_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11505__A1 _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11505__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17283__B _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19857_ _19857_/A _19857_/B _19857_/C vssd1 vssd1 vccd1 vccd1 _19857_/Y sky130_fd_sc_hd__nand3_1
X_18808_ _18807_/B _18807_/C _18807_/A vssd1 vssd1 vccd1 vccd1 _18810_/B sky130_fd_sc_hd__a21o_1
X_19788_ _19788_/A _19788_/B _19788_/C vssd1 vssd1 vccd1 vccd1 _19788_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__12501__A _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18739_ _20317_/D _19060_/B _18741_/C _18741_/D vssd1 vssd1 vccd1 vccd1 _18739_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14314__A1_N _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21750_ _22038_/CLK _21750_/D vssd1 vssd1 vccd1 vccd1 _21750_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16747__A2 _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19493__A_N _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20701_ _20699_/B _20699_/C _20699_/A vssd1 vssd1 vccd1 vccd1 _20701_/Y sky130_fd_sc_hd__a21oi_1
X_21681_ _21682_/CLK _21681_/D vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_47_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout247_A _21807_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20632_ _20496_/A _20499_/C _20630_/Y _20631_/X vssd1 vssd1 vccd1 vccd1 _20632_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_74_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18842__B _18842_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11441__B1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17739__A _18010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20563_ _21171_/A _21264_/B _20561_/Y _20685_/A vssd1 vssd1 vccd1 vccd1 _20565_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout414_A _21766_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20144__A1_N _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20494_ _20299_/A _20300_/X _20492_/A _20493_/Y vssd1 vssd1 vccd1 vccd1 _20496_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21115_ _21112_/X _21113_/Y _20998_/Y _21000_/Y vssd1 vssd1 vccd1 vccd1 _21116_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_1_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout210 _21815_/Q vssd1 vssd1 vccd1 vccd1 _21264_/B sky130_fd_sc_hd__buf_4
X_22095_ _22105_/CLK _22095_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[31] sky130_fd_sc_hd__dfrtp_4
Xfanout221 _21311_/A vssd1 vssd1 vccd1 vccd1 _18789_/B sky130_fd_sc_hd__buf_2
XFILLER_0_121_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout232 hold331/X vssd1 vssd1 vccd1 vccd1 _17670_/B sky130_fd_sc_hd__buf_4
X_21046_ _21256_/A _21046_/B _21046_/C _21046_/D vssd1 vssd1 vccd1 vccd1 _21161_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__17193__B _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout243 _19692_/A vssd1 vssd1 vccd1 vccd1 _19535_/A sky130_fd_sc_hd__buf_4
Xfanout254 _18166_/A vssd1 vssd1 vccd1 vccd1 _19382_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_22_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout265 _19531_/A vssd1 vssd1 vccd1 vccd1 _20590_/D sky130_fd_sc_hd__buf_4
Xfanout276 _18008_/A vssd1 vssd1 vccd1 vccd1 _20317_/D sky130_fd_sc_hd__buf_4
Xfanout287 _21798_/Q vssd1 vssd1 vccd1 vccd1 _18010_/A sky130_fd_sc_hd__buf_4
Xfanout298 _17063_/C vssd1 vssd1 vccd1 vccd1 _17013_/D sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout62_A _21853_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14997__A1 _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14997__B2 _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20519__B1 _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12750_ _12750_/A _15768_/A vssd1 vssd1 vccd1 vccd1 _12754_/A sky130_fd_sc_hd__nand2_1
X_21948_ _21948_/CLK _21948_/D vssd1 vssd1 vccd1 vccd1 hold195/A sky130_fd_sc_hd__dfxtp_1
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11701_ _11701_/A _12318_/B _11701_/C vssd1 vssd1 vccd1 vccd1 _12297_/A sky130_fd_sc_hd__and3_1
XFILLER_0_84_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ _12681_/A _12681_/B _12681_/C vssd1 vssd1 vccd1 vccd1 _12684_/A sky130_fd_sc_hd__nand3_2
X_21879_ _21945_/CLK _21879_/D vssd1 vssd1 vccd1 vccd1 hold78/A sky130_fd_sc_hd__dfxtp_2
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11461__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14420_ _14255_/A _14255_/C _14255_/B vssd1 vssd1 vccd1 vccd1 _14422_/B sky130_fd_sc_hd__a21bo_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ _11625_/X _11787_/A _11683_/B _11631_/X vssd1 vssd1 vccd1 vccd1 _11632_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14351_ _14351_/A _14351_/B vssd1 vssd1 vccd1 vccd1 _14361_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11563_ _12229_/A _12750_/A _12528_/B _12155_/B vssd1 vssd1 vccd1 vccd1 _11563_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13302_ _13302_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13304_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17070_ _17068_/A _17068_/B _17068_/C vssd1 vssd1 vccd1 vccd1 _17071_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_122_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14282_ _14282_/A _14282_/B vssd1 vssd1 vccd1 vccd1 _14284_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_80_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11494_ _11493_/X _18769_/B _11521_/S vssd1 vssd1 vccd1 vccd1 _21836_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_80_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16021_ _16021_/A _16021_/B _16021_/C vssd1 vssd1 vccd1 vccd1 _16023_/A sky130_fd_sc_hd__and3_1
XFILLER_0_134_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13233_ _13822_/B _13381_/C _14155_/C _14155_/D vssd1 vssd1 vccd1 vccd1 _13376_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_126_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13164_ _13164_/A _13287_/B _13164_/C vssd1 vssd1 vccd1 vccd1 _13166_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_62_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15319__D _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12115_ _12115_/A _12115_/B _12115_/C vssd1 vssd1 vccd1 vccd1 _12115_/X sky130_fd_sc_hd__or3_1
XANTENNA__17384__A _21792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13095_ hold107/X _13094_/X fanout2/X vssd1 vssd1 vccd1 vccd1 hold108/A sky130_fd_sc_hd__mux2_1
X_17972_ hold155/A fanout8/X _17970_/X _11550_/A _17971_/Y vssd1 vssd1 vccd1 vccd1
+ _17972_/X sky130_fd_sc_hd__a221o_1
X_19711_ _19711_/A _19711_/B _19711_/C vssd1 vssd1 vccd1 vccd1 _19715_/B sky130_fd_sc_hd__nand3_2
X_16923_ _16923_/A _16923_/B _16923_/C vssd1 vssd1 vccd1 vccd1 _16930_/A sky130_fd_sc_hd__nand3_1
X_12046_ _12044_/X _12046_/B vssd1 vssd1 vccd1 vccd1 _12048_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_137_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19642_ _19560_/A _19560_/C _19560_/B vssd1 vssd1 vccd1 vccd1 _19681_/A sky130_fd_sc_hd__a21bo_1
X_16854_ _16785_/X _16852_/Y _16859_/A _16851_/A vssd1 vssd1 vccd1 vccd1 _16855_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18927__B _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15805_ _15808_/D vssd1 vssd1 vccd1 vccd1 _15805_/Y sky130_fd_sc_hd__inv_2
X_19573_ _20650_/A _19414_/C _19575_/C _19575_/D vssd1 vssd1 vccd1 vccd1 _19573_/X
+ sky130_fd_sc_hd__a22o_1
X_13997_ _15159_/D _14936_/D _13997_/C _14155_/C vssd1 vssd1 vccd1 vccd1 _14153_/A
+ sky130_fd_sc_hd__nand4_2
X_16785_ _16785_/A _16785_/B _16785_/C vssd1 vssd1 vccd1 vccd1 _16785_/X sky130_fd_sc_hd__and3_2
XFILLER_0_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15632__A _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18524_ _18521_/X _18522_/Y _18373_/C _18372_/Y vssd1 vssd1 vccd1 vccd1 _18525_/D
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_38_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15736_ _15733_/X _15734_/Y _15563_/Y _15567_/B vssd1 vssd1 vccd1 vccd1 _15737_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_3170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12948_ _13091_/A _12950_/B _12950_/C vssd1 vssd1 vccd1 vccd1 _12951_/A sky130_fd_sc_hd__a21oi_1
XTAP_3181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16447__B _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18455_ _18454_/A _18454_/B _18441_/X vssd1 vssd1 vccd1 vccd1 _18455_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_34_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15674__A1_N _15933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15667_ _15667_/A _15667_/B vssd1 vssd1 vccd1 vccd1 _15668_/B sky130_fd_sc_hd__nand2_1
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ _13152_/C _12877_/X _12878_/X vssd1 vssd1 vccd1 vccd1 _12880_/B sky130_fd_sc_hd__a21bo_1
XANTENNA_170 v2z[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14248__A _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11371__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13152__A _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_181 v2z[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_192 hold247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17406_ _17405_/B _17405_/C _17405_/A vssd1 vssd1 vccd1 vccd1 _17406_/X sky130_fd_sc_hd__o21a_1
X_14618_ _14618_/A _14618_/B vssd1 vssd1 vccd1 vccd1 _14620_/A sky130_fd_sc_hd__xnor2_4
X_15598_ _15598_/A _15598_/B vssd1 vssd1 vccd1 vccd1 _15600_/C sky130_fd_sc_hd__xnor2_2
X_18386_ _18386_/A _18386_/B vssd1 vssd1 vccd1 vccd1 _18388_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_55_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14549_ _14551_/B vssd1 vssd1 vccd1 vccd1 _14549_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17337_ _17915_/A _19445_/A vssd1 vssd1 vccd1 vccd1 _17340_/A sky130_fd_sc_hd__and2_1
XFILLER_0_71_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12991__A _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17268_ _17372_/A _17372_/B _17379_/A vssd1 vssd1 vccd1 vccd1 _17269_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_71_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19007_ _19007_/A _19007_/B vssd1 vssd1 vccd1 vccd1 _19046_/A sky130_fd_sc_hd__nor2_2
XANTENNA__20416__C _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15079__A _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16219_ _16219_/A _16323_/B vssd1 vssd1 vccd1 vccd1 _16221_/B sky130_fd_sc_hd__or2_1
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17199_ _17199_/A _17199_/B vssd1 vssd1 vccd1 vccd1 _17219_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18103__B2 _11547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11726__B2 _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19851__A1 _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19493__B _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15229__D _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12215__B _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19851__B2 _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14133__D _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17862__B1 _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19909_ _19909_/A _19909_/B _20001_/B vssd1 vssd1 vccd1 vccd1 _19911_/B sky130_fd_sc_hd__nand3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12151__A1 _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16417__A1 _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21410__A1 _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17741__B _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout364_A _21778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21802_ _21803_/CLK _21802_/D vssd1 vssd1 vccd1 vccd1 _21802_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_91_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18556__C _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15261__B _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21733_ _21803_/CLK _21733_/D vssd1 vssd1 vccd1 vccd1 _21733_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_19_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout531_A _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20921__B1 _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout629_A _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13403__A1 _14463_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21664_ _21906_/CLK _21664_/D vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13997__A _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20615_ _20616_/A _20616_/B _20616_/C vssd1 vssd1 vccd1 vccd1 _20615_/X sky130_fd_sc_hd__a21o_1
X_21595_ _21934_/CLK _21595_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[58] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_959 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12109__C _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20546_ _21258_/A _21305_/A _21153_/B _20797_/A vssd1 vssd1 vccd1 vccd1 _20550_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18893__A2 _18894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14605__B _14605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17619__D _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13706__A2 _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20477_ _20583_/A _20193_/D _20475_/Y _20602_/A vssd1 vssd1 vccd1 vccd1 _20479_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_131_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22078_ _22080_/CLK _22078_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[14] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12142__A1 _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12142__B2 _12242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13920_ _14713_/B _15370_/B _15098_/B _14713_/A vssd1 vssd1 vccd1 vccd1 _13920_/Y
+ sky130_fd_sc_hd__a22oi_1
X_21029_ hold77/X fanout8/X _21027_/Y _11550_/A _21028_/Y vssd1 vssd1 vccd1 vccd1
+ _21029_/X sky130_fd_sc_hd__a221o_1
XANTENNA__15155__C _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13851_ _13851_/A _13973_/A _13851_/C vssd1 vssd1 vccd1 vccd1 _13973_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_18_1109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12802_ _12803_/A _12803_/B _12803_/C _12803_/D vssd1 vssd1 vccd1 vccd1 _12802_/Y
+ sky130_fd_sc_hd__nor4_2
X_13782_ _13782_/A _13782_/B _13782_/C vssd1 vssd1 vccd1 vccd1 _13784_/B sky130_fd_sc_hd__nand3_1
X_16570_ _17621_/C _17300_/C _17520_/D _17504_/C vssd1 vssd1 vccd1 vccd1 _16571_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10994_ mstream_o[68] hold86/X _11005_/S vssd1 vssd1 vccd1 vccd1 _21605_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12445__A2 _12771_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15521_ _16031_/A _15521_/B vssd1 vssd1 vccd1 vccd1 _15523_/B sky130_fd_sc_hd__xnor2_1
X_12733_ _13860_/A _13554_/B _12858_/C _13269_/D vssd1 vssd1 vccd1 vccd1 _12856_/A
+ sky130_fd_sc_hd__and4_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_128_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15452_ _16087_/A _15717_/C _15976_/D _16092_/D vssd1 vssd1 vccd1 vccd1 _15456_/D
+ sky130_fd_sc_hd__a22o_1
X_18240_ _18240_/A _18241_/A _18389_/A vssd1 vssd1 vccd1 vccd1 _18240_/X sky130_fd_sc_hd__or3b_2
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ _12665_/A _12665_/B vssd1 vssd1 vccd1 vccd1 _12766_/A sky130_fd_sc_hd__nand2b_2
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14403_ _14403_/A _14403_/B vssd1 vssd1 vccd1 vccd1 _14412_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_65_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11615_ _12302_/A _12858_/C _12991_/D _13985_/A vssd1 vssd1 vccd1 vccd1 _11615_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11405__B1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15383_ _15384_/A _15384_/B _15384_/C vssd1 vssd1 vccd1 vccd1 _15386_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_143_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18171_ _19535_/A _19695_/A _18319_/B _18622_/B vssd1 vssd1 vccd1 vccd1 _18322_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_53_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12595_ _12592_/X _12593_/Y _12481_/Y _12484_/X vssd1 vssd1 vccd1 vccd1 _12596_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_136_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18333__A1 _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14334_ _14333_/B _14333_/C _14322_/Y vssd1 vssd1 vccd1 vccd1 _14334_/Y sky130_fd_sc_hd__a21boi_1
X_17122_ _17089_/A _17089_/C _17089_/B vssd1 vssd1 vccd1 vccd1 _17122_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11546_ _21725_/D _11555_/B vssd1 vssd1 vccd1 vccd1 _20770_/B sky130_fd_sc_hd__nor2_8
XFILLER_0_29_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17053_ _17144_/A _17124_/C _17145_/B _17129_/B vssd1 vssd1 vccd1 vccd1 _17054_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14265_ _14264_/B _14264_/C _14264_/A vssd1 vssd1 vccd1 vccd1 _14265_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_34_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11477_ _11498_/A1 t1y[9] t0x[9] _11501_/B2 vssd1 vssd1 vccd1 vccd1 _11477_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_150_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16004_ _16001_/X _16002_/Y _15870_/Y _15874_/C vssd1 vssd1 vccd1 vccd1 _16004_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_33_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14234__C _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13216_ _13213_/Y _13214_/X _13074_/X _13077_/X vssd1 vssd1 vccd1 vccd1 _13218_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_122_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14196_ _14196_/A _14196_/B _14362_/B vssd1 vssd1 vccd1 vccd1 _14198_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13147_ _13230_/A _13145_/X _13002_/B _13003_/Y vssd1 vssd1 vccd1 vccd1 _13209_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12671__A1_N _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13078_ _13077_/B _13077_/C _13077_/A vssd1 vssd1 vccd1 vccd1 _13078_/Y sky130_fd_sc_hd__a21oi_1
X_17955_ _17812_/X _17815_/X _17953_/X _17954_/Y vssd1 vssd1 vccd1 vccd1 _17958_/B
+ sky130_fd_sc_hd__o211ai_4
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16906_ _16901_/A _16952_/A _16895_/X vssd1 vssd1 vccd1 vccd1 _16908_/B sky130_fd_sc_hd__a21o_1
X_12029_ _12029_/A _12029_/B _12029_/C vssd1 vssd1 vccd1 vccd1 _12030_/B sky130_fd_sc_hd__and3_1
X_17886_ _17772_/Y _17776_/A _17884_/A _17885_/Y vssd1 vssd1 vccd1 vccd1 _17975_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_75_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21364__A _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19625_ _19626_/A _19626_/B vssd1 vssd1 vccd1 vccd1 _19779_/B sky130_fd_sc_hd__nand2_1
X_16837_ _16894_/A _16894_/B vssd1 vssd1 vccd1 vccd1 _16837_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__16458__A _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19556_ _19556_/A _19556_/B _19556_/C vssd1 vssd1 vccd1 vccd1 _19556_/X sky130_fd_sc_hd__and3_1
X_16768_ _17300_/C _17520_/D _17277_/A _17387_/A vssd1 vssd1 vccd1 vccd1 _16849_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__11239__A3 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18507_ _18357_/A _18357_/C _18357_/B vssd1 vssd1 vccd1 vccd1 _18508_/C sky130_fd_sc_hd__a21bo_1
X_15719_ _15848_/A _15978_/B _16087_/A _15719_/D vssd1 vssd1 vccd1 vccd1 _15848_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_75_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19487_ _19487_/A _19487_/B _20838_/D vssd1 vssd1 vccd1 vccd1 _19487_/X sky130_fd_sc_hd__and3_1
XFILLER_0_75_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16699_ _16698_/B _16698_/C _16698_/A vssd1 vssd1 vccd1 vccd1 _16701_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__17375__A2 _12493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18438_ _18438_/A _18438_/B vssd1 vssd1 vccd1 vccd1 _18440_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_29_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_926 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18369_ _18368_/A _18368_/B _18368_/C _18368_/D vssd1 vssd1 vccd1 vccd1 _18369_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_28_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11947__A1 _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20400_ _20913_/A _20401_/B vssd1 vssd1 vccd1 vccd1 _20400_/X sky130_fd_sc_hd__and2_1
X_21380_ _21381_/B _21379_/X _21378_/Y vssd1 vssd1 vccd1 vccd1 _21934_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20146__C _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20331_ _20838_/B _21283_/B _21305_/B _20975_/D vssd1 vssd1 vccd1 vccd1 _20335_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19824__A1 _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20262_ _20096_/Y _20120_/Y _20259_/Y _20260_/X vssd1 vssd1 vccd1 vccd1 _20302_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_101_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16638__A1 _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22001_ _22005_/CLK _22001_/D vssd1 vssd1 vccd1 vccd1 hold142/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__17835__B1 _11553_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16638__B2 _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21258__B _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20193_ _20190_/Y _20329_/A _20721_/D _20193_/D vssd1 vssd1 vccd1 vccd1 _20329_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_110_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13983__C _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19951__B _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13321__B1 _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout579_A _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11276__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19588__B1 _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13872__A1 _13875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12675__A2 _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16087__B _21787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_94_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21716_ _21722_/CLK _21716_/D _21329_/B1 vssd1 vssd1 vccd1 vccd1 sstream_o sky130_fd_sc_hd__dfstp_4
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout25_A _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16815__B _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21647_ _21722_/CLK hold307/X fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[110]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18315__A1 _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11400_ hold269/X fanout28/X _11399_/X vssd1 vssd1 vccd1 vccd1 _11400_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_151_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15129__A1 _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15129__B2 _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12060__B1 _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12380_ _12379_/B _12379_/C _12379_/A vssd1 vssd1 vccd1 vccd1 _12380_/X sky130_fd_sc_hd__a21o_1
XANTENNA_70 hold268/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21578_ mstream_o[41] _11063_/X _21579_/S vssd1 vssd1 vccd1 vccd1 _22105_/D sky130_fd_sc_hd__mux2_1
XANTENNA_81 hold234/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_92 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12781__D _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ fanout58/X v0z[26] fanout18/X _11330_/X vssd1 vssd1 vccd1 vccd1 _11331_/X
+ sky130_fd_sc_hd__a31o_2
XANTENNA__16877__A1 _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20673__A2 _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16877__B2 _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20529_ _20529_/A _20529_/B vssd1 vssd1 vccd1 vccd1 _20531_/B sky130_fd_sc_hd__xnor2_1
X_14050_ _14132_/A _14048_/Y _13884_/B _13884_/Y vssd1 vssd1 vccd1 vccd1 _14109_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14352__A2 _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11262_ _11502_/A1 t1x[9] v2z[9] _11501_/B2 _11261_/X vssd1 vssd1 vccd1 vccd1 _11262_/X
+ sky130_fd_sc_hd__a221o_2
X_13001_ _13000_/A _13000_/B _13000_/C vssd1 vssd1 vccd1 vccd1 _13002_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13893__C _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11193_ hold297/X fanout51/X fanout47/X hold305/A vssd1 vssd1 vccd1 vccd1 _11193_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11694__B _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11186__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17740_ _18010_/A _17739_/C _17739_/D _17874_/A vssd1 vssd1 vccd1 vccd1 _17741_/D
+ sky130_fd_sc_hd__a22o_1
X_14952_ _14952_/A _14952_/B _15169_/B vssd1 vssd1 vccd1 vccd1 _14954_/B sky130_fd_sc_hd__nand3_2
XANTENNA__20189__A1 _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20189__B2 fanout96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20800__B _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13903_ _13900_/Y _13901_/X _13750_/D _13751_/B vssd1 vssd1 vccd1 vccd1 _13904_/C
+ sky130_fd_sc_hd__o211ai_2
X_17671_ _19123_/A _19123_/B _20270_/C _18789_/B vssd1 vssd1 vccd1 vccd1 _17673_/B
+ sky130_fd_sc_hd__nand4_1
X_14883_ _14883_/A _14883_/B _14883_/C vssd1 vssd1 vccd1 vccd1 _14883_/X sky130_fd_sc_hd__and3_2
XFILLER_0_138_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19410_ _19906_/D _19409_/X _19408_/X vssd1 vssd1 vccd1 vccd1 _19412_/A sky130_fd_sc_hd__a21bo_1
X_16622_ _16622_/A _16622_/B _16622_/C vssd1 vssd1 vccd1 vccd1 _16642_/A sky130_fd_sc_hd__nand3_1
X_13834_ _13834_/A _13834_/B vssd1 vssd1 vccd1 vccd1 _13851_/A sky130_fd_sc_hd__or2_1
XFILLER_0_58_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19341_ _19341_/A _19341_/B vssd1 vssd1 vccd1 vccd1 _19343_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13765_ _14859_/A _14218_/B _13766_/C _13910_/A vssd1 vssd1 vccd1 vccd1 _13767_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16553_ _16553_/A _16553_/B vssd1 vssd1 vccd1 vccd1 _16686_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11626__B1 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10977_ _10977_/A _10977_/B vssd1 vssd1 vccd1 vccd1 _10978_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_35_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15504_ _15907_/A _16261_/B vssd1 vssd1 vccd1 vccd1 _16036_/A sky130_fd_sc_hd__or2_4
X_19272_ _19406_/B _19271_/C _19271_/A vssd1 vssd1 vccd1 vccd1 _19272_/Y sky130_fd_sc_hd__a21oi_1
X_12716_ _12716_/A _12716_/B _12716_/C vssd1 vssd1 vccd1 vccd1 _12717_/B sky130_fd_sc_hd__and3_1
XFILLER_0_155_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13696_ _13691_/Y _13693_/X _13538_/Y _13541_/X vssd1 vssd1 vccd1 vccd1 _13698_/C
+ sky130_fd_sc_hd__o211a_1
X_16484_ _16485_/A _16485_/B vssd1 vssd1 vccd1 vccd1 _16484_/X sky130_fd_sc_hd__and2_1
XANTENNA__16725__B _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18223_ _18220_/X _18221_/Y _18082_/B _18081_/Y vssd1 vssd1 vccd1 vccd1 _18225_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15435_ _15435_/A _15698_/B _15435_/C _15435_/D vssd1 vssd1 vccd1 vccd1 _15577_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_66_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12647_ _12637_/A _13157_/B _12536_/B _12534_/X vssd1 vssd1 vccd1 vccd1 _12649_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20247__B _21832_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15366_ _15221_/A _15220_/B _15218_/X vssd1 vssd1 vccd1 vccd1 _15382_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_143_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18154_ _18014_/A _18014_/C _18014_/B vssd1 vssd1 vccd1 vccd1 _18155_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_25_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12578_ _12578_/A _12578_/B _12578_/C vssd1 vssd1 vccd1 vccd1 _12578_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_41_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17105_ _17101_/A _17101_/B _17101_/C vssd1 vssd1 vccd1 vccd1 _17106_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14317_ _14317_/A _14317_/B _14317_/C vssd1 vssd1 vccd1 vccd1 _14319_/A sky130_fd_sc_hd__nor3_1
X_11529_ _11544_/A1 t2x[26] v1z[26] fanout21/X _11528_/X vssd1 vssd1 vccd1 vccd1 _11529_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15297_ _15297_/A vssd1 vssd1 vccd1 vccd1 _15338_/A sky130_fd_sc_hd__inv_2
X_18085_ _18082_/X _18083_/Y _17948_/B _17947_/Y vssd1 vssd1 vccd1 vccd1 _18087_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_29_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold307 hold307/A vssd1 vssd1 vccd1 vccd1 hold307/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold318 hold318/A vssd1 vssd1 vccd1 vccd1 hold318/X sky130_fd_sc_hd__dlygate4sd3_1
X_14248_ _14248_/A _21759_/Q _16173_/B vssd1 vssd1 vccd1 vccd1 _14572_/B sky130_fd_sc_hd__and3_1
X_17036_ _17058_/A _17036_/B vssd1 vssd1 vccd1 vccd1 _17038_/B sky130_fd_sc_hd__xnor2_1
Xhold329 hold329/A vssd1 vssd1 vccd1 vccd1 hold329/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17556__B _17924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14179_ _14179_/A _14179_/B vssd1 vssd1 vccd1 vccd1 _14189_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_110_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15076__B _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18987_ _18987_/A _18987_/B _18985_/Y _18986_/X vssd1 vssd1 vccd1 vccd1 _18987_/X
+ sky130_fd_sc_hd__or4bb_2
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17938_ _17937_/B _17937_/C _17937_/A vssd1 vssd1 vccd1 vccd1 _17940_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12657__A2 _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17869_ _17869_/A _17869_/B vssd1 vssd1 vccd1 vccd1 _17883_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_75_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19608_ _19608_/A _19608_/B vssd1 vssd1 vccd1 vccd1 _19609_/B sky130_fd_sc_hd__and2_1
XFILLER_0_89_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16619__C _17334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20880_ _20881_/A _20880_/B _20880_/C vssd1 vssd1 vccd1 vccd1 _20880_/X sky130_fd_sc_hd__or3_1
XANTENNA__13324__B _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19539_ _19378_/X _19381_/X _19536_/X _19538_/Y vssd1 vssd1 vccd1 vccd1 _19539_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16556__B1 _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21501_ hold304/X sstream_i[78] _21510_/S vssd1 vssd1 vccd1 vccd1 _22028_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_5_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout327_A _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12882__C _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21432_ hold242/X sstream_i[9] _21442_/S vssd1 vssd1 vccd1 vccd1 _21959_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_146_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18848__A2 _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14155__B _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21363_ hold136/X fanout40/X _21362_/X vssd1 vssd1 vccd1 vccd1 _21928_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_32_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20314_ _20314_/A _20314_/B vssd1 vssd1 vccd1 vccd1 _20316_/B sky130_fd_sc_hd__or2_1
XFILLER_0_3_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21294_ _21294_/A _21294_/B vssd1 vssd1 vccd1 vccd1 _21295_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__20173__A _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20245_ _20245_/A _20428_/B vssd1 vssd1 vccd1 vccd1 _20255_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17284__A1 _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17284__B2 _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20176_ _20176_/A _20314_/B _20177_/B vssd1 vssd1 vccd1 vccd1 _20176_/X sky130_fd_sc_hd__or3b_1
XANTENNA__12403__B _12403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_hold274_A hold274/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21368__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10900_ _10885_/A _10885_/B _10885_/C _10892_/A vssd1 vssd1 vccd1 vccd1 _10902_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_3758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16529__C _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11880_ _11881_/A _11881_/B vssd1 vssd1 vccd1 vccd1 _11880_/X sky130_fd_sc_hd__and2_1
XTAP_3769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10831_ _11045_/A _10828_/Y _10830_/A vssd1 vssd1 vccd1 vccd1 _11048_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_79_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17339__A2 _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13550_ _13392_/Y _13395_/X _13548_/A _13549_/X vssd1 vssd1 vccd1 vccd1 _13652_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_55_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12501_ _14133_/D _13983_/B _13258_/C _13258_/D vssd1 vssd1 vccd1 vccd1 _12503_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_48_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13481_ _13480_/B _13480_/C _13480_/A vssd1 vssd1 vccd1 vccd1 _13483_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14022__A1 _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14022__B2 _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15220_ _15218_/X _15220_/B vssd1 vssd1 vccd1 vccd1 _15362_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12432_ _12433_/A _12433_/B vssd1 vssd1 vccd1 vccd1 _12432_/X sky130_fd_sc_hd__and2_2
XFILLER_0_152_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15151_ _15151_/A _15151_/B vssd1 vssd1 vccd1 vccd1 _15192_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_106_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17657__A _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12363_ _12362_/A _12362_/B _12362_/C vssd1 vssd1 vccd1 vccd1 _12364_/C sky130_fd_sc_hd__a21o_1
XANTENNA__16561__A _21830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14102_ _14101_/B _14101_/C _14101_/A vssd1 vssd1 vccd1 vccd1 _14102_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_22_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11314_ _11224_/A t1x[22] v2z[22] _11223_/A _11313_/X vssd1 vssd1 vccd1 vccd1 _11314_/X
+ sky130_fd_sc_hd__a221o_2
X_15082_ _15082_/A _15082_/B _15082_/C vssd1 vssd1 vccd1 vccd1 _15085_/C sky130_fd_sc_hd__and3_1
XANTENNA__14325__A2 _14477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12294_ _12035_/A _12294_/B _12294_/C _12294_/D vssd1 vssd1 vccd1 vccd1 _12294_/X
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14033_ _21742_/Q _14537_/A _13892_/X _13893_/X _14365_/D vssd1 vssd1 vccd1 vccd1
+ _14038_/A sky130_fd_sc_hd__a32o_1
X_18910_ _19379_/B _19238_/C _18911_/C _19065_/A vssd1 vssd1 vccd1 vccd1 _18912_/B
+ sky130_fd_sc_hd__a22o_1
X_11245_ _11122_/A t2y[5] t0y[5] _11123_/A vssd1 vssd1 vccd1 vccd1 _11245_/X sky130_fd_sc_hd__a22o_1
XANTENNA__19872__A _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19890_ _20838_/B _20975_/D _21278_/A _20265_/D vssd1 vssd1 vccd1 vccd1 _19891_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_129_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18841_ _18841_/A _18841_/B vssd1 vssd1 vccd1 vccd1 _18842_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_38_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11176_ hold154/X fanout22/X _11175_/X vssd1 vssd1 vccd1 vccd1 _11176_/X sky130_fd_sc_hd__a21o_1
X_18772_ _19972_/A _20394_/B _19546_/D _19906_/C vssd1 vssd1 vccd1 vccd1 _18775_/B
+ sky130_fd_sc_hd__nand4_1
X_15984_ _15986_/A _15986_/B _15986_/C vssd1 vssd1 vccd1 vccd1 _15984_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__13836__A1 _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21359__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13836__B2 _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17723_ _17720_/X _17723_/B _18703_/A _19053_/B vssd1 vssd1 vccd1 vccd1 _17725_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_145_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14935_ _14935_/A _14935_/B vssd1 vssd1 vccd1 vccd1 _14940_/A sky130_fd_sc_hd__or2_1
XFILLER_0_136_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15589__A1 _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17654_ _17531_/X _17533_/X _17651_/X _17652_/Y vssd1 vssd1 vccd1 vccd1 _17654_/Y
+ sky130_fd_sc_hd__o211ai_4
X_14866_ _14721_/X _14734_/A _14734_/B _14723_/B vssd1 vssd1 vccd1 vccd1 _14868_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__20582__A1 _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20582__B2 _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16605_ _19445_/A _17334_/B vssd1 vssd1 vccd1 vccd1 _16608_/A sky130_fd_sc_hd__and2_1
X_13817_ hold29/X _13816_/X fanout1/X vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__mux2_1
X_17585_ _17584_/B _17584_/C _17584_/A vssd1 vssd1 vccd1 vccd1 _17586_/B sky130_fd_sc_hd__a21oi_1
X_14797_ _14640_/B _14642_/B _14795_/X _14796_/Y vssd1 vssd1 vccd1 vccd1 _14797_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_147_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19324_ _20770_/B _19322_/Y _19323_/X vssd1 vssd1 vccd1 vccd1 _19324_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21361__B _21361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16536_ _16534_/B _16534_/C _16534_/A vssd1 vssd1 vccd1 vccd1 _16537_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_70_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21531__A0 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13748_ _15514_/A _15514_/B _14212_/C _14212_/D vssd1 vssd1 vccd1 vccd1 _13750_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_85_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19255_ _19115_/A _19114_/B _19112_/X vssd1 vssd1 vccd1 vccd1 _19271_/A sky130_fd_sc_hd__a21o_1
X_16467_ _17206_/B _17124_/C _16466_/B _16463_/X vssd1 vssd1 vccd1 vccd1 _16468_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_39_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13679_ _14138_/A _14155_/C _14155_/D _13975_/B vssd1 vssd1 vccd1 vccd1 _13679_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__18951__A _19732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18206_ _18066_/A _18066_/C _18066_/B vssd1 vssd1 vccd1 vccd1 _18207_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_143_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15418_ _15419_/A _15419_/B _15419_/C vssd1 vssd1 vccd1 vccd1 _15420_/B sky130_fd_sc_hd__a21o_2
XFILLER_0_115_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14564__A2 _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19186_ _19188_/A vssd1 vssd1 vccd1 vccd1 _19345_/A sky130_fd_sc_hd__inv_2
X_16398_ _16398_/A _16398_/B vssd1 vssd1 vccd1 vccd1 _16413_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13772__B1 _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18137_ _18873_/A _19382_/B _18288_/A _18137_/D vssd1 vssd1 vccd1 vccd1 _18288_/B
+ sky130_fd_sc_hd__nand4_1
X_15349_ _15350_/A _15350_/B vssd1 vssd1 vccd1 vccd1 _15349_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold104 hold104/A vssd1 vssd1 vccd1 vccd1 hold104/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold115 hold115/A vssd1 vssd1 vccd1 vccd1 hold115/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 hold126/A vssd1 vssd1 vccd1 vccd1 hold126/X sky130_fd_sc_hd__dlygate4sd3_1
X_18068_ _17932_/A _17932_/C _17932_/B vssd1 vssd1 vccd1 vccd1 _18069_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_106_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold137 hold137/A vssd1 vssd1 vccd1 vccd1 hold137/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12327__A1 _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13524__B1 _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold148 hold148/A vssd1 vssd1 vccd1 vccd1 hold148/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12327__B2 _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold159 hold159/A vssd1 vssd1 vccd1 vccd1 hold159/X sky130_fd_sc_hd__dlygate4sd3_1
X_17019_ _17144_/A _17129_/B _17019_/C _17124_/C vssd1 vssd1 vccd1 vccd1 _17019_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_10_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12504__A _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12878__A2 _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout606 _21719_/Q vssd1 vssd1 vccd1 vccd1 _11459_/B2 sky130_fd_sc_hd__clkbuf_8
Xfanout617 _21717_/Q vssd1 vssd1 vccd1 vccd1 _11005_/S sky130_fd_sc_hd__clkbuf_8
X_20030_ _19804_/D _19808_/B _20027_/X _20175_/B vssd1 vssd1 vccd1 vccd1 _20031_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13319__B _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout628 _21087_/D vssd1 vssd1 vccd1 vccd1 _20838_/B sky130_fd_sc_hd__buf_4
XFILLER_0_95_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout639 _21422_/A vssd1 vssd1 vccd1 vccd1 fanout639/X sky130_fd_sc_hd__clkbuf_8
XANTENNA__12223__B _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21981_ _22013_/CLK _21981_/D vssd1 vssd1 vccd1 vccd1 hold148/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout277_A _21800_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18766__A1 _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18766__B2 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20932_ _20932_/A _21048_/B _20931_/X vssd1 vssd1 vccd1 vccd1 _21110_/A sky130_fd_sc_hd__or3b_2
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20863_ _20985_/A _21311_/B _20863_/C _20863_/D vssd1 vssd1 vccd1 vccd1 _20985_/B
+ sky130_fd_sc_hd__and4b_1
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21522__A0 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20794_ _21286_/A _21264_/A _20794_/C _20986_/A vssd1 vssd1 vccd1 vccd1 _20986_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_77_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19379__D _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout611_A _21718_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16084__C _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14555__A2 _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12566__A1 _12785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13763__B1 _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21415_ _21720_/D _21415_/B vssd1 vssd1 vccd1 vccd1 _21415_/X sky130_fd_sc_hd__or2_1
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12566__B2 _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16812__C _17063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21346_ _21349_/A _21346_/B vssd1 vssd1 vccd1 vccd1 _21346_/X sky130_fd_sc_hd__or2_1
XFILLER_0_102_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13515__B1 _11066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19692__A _19692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21277_ _21277_/A _21277_/B vssd1 vssd1 vccd1 vccd1 _21279_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout92_A _21844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11030_ mstream_o[104] hold286/X _11039_/S vssd1 vssd1 vccd1 vccd1 hold287/A sky130_fd_sc_hd__mux2_1
X_20228_ _20372_/B _20228_/B vssd1 vssd1 vccd1 vccd1 _21396_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__17924__B _17924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20159_ _20159_/A _20159_/B vssd1 vssd1 vccd1 vccd1 _20161_/B sky130_fd_sc_hd__xnor2_2
XTAP_3500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12981_ _14306_/A _13258_/C _13258_/D _14138_/A vssd1 vssd1 vccd1 vccd1 _12982_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11464__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14720_ _14717_/X _14719_/Y _14571_/A _14974_/A vssd1 vssd1 vccd1 vccd1 _14723_/A
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11932_ _12897_/C _13556_/A _12214_/C _12897_/D vssd1 vssd1 vccd1 vccd1 _11933_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14651_ _14652_/B _14652_/A vssd1 vssd1 vccd1 vccd1 _14764_/A sky130_fd_sc_hd__and2b_1
X_11863_ _12109_/C _12621_/C _11862_/B _11859_/X vssd1 vssd1 vccd1 vccd1 _11869_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_3599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14243__A1 _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13602_ _13602_/A _13602_/B vssd1 vssd1 vccd1 vccd1 _13605_/C sky130_fd_sc_hd__xor2_1
X_10814_ hold221/A hold80/A vssd1 vssd1 vccd1 vccd1 _10815_/B sky130_fd_sc_hd__or2_1
XTAP_2898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17370_ _17379_/A _17379_/B _17479_/A vssd1 vssd1 vccd1 vccd1 _17371_/B sky130_fd_sc_hd__o21a_1
XANTENNA__13899__B _14212_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14582_ _14583_/A _14583_/B vssd1 vssd1 vccd1 vccd1 _14582_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11794_ _11795_/A _11795_/B _11795_/C vssd1 vssd1 vccd1 vccd1 _11794_/X sky130_fd_sc_hd__and3_1
X_16321_ _16321_/A _16321_/B vssd1 vssd1 vccd1 vccd1 _16341_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_27_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13533_ _13530_/X _13678_/B _13404_/D _13405_/B vssd1 vssd1 vccd1 vccd1 _13534_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_83_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19040_ _19037_/X _19038_/Y _18876_/B _18878_/B vssd1 vssd1 vccd1 vccd1 _19040_/Y
+ sky130_fd_sc_hd__o211ai_2
X_16252_ _16253_/A _16253_/B vssd1 vssd1 vccd1 vccd1 _16366_/B sky130_fd_sc_hd__and2b_1
X_13464_ _13464_/A _13464_/B vssd1 vssd1 vccd1 vccd1 _13466_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12006__B1 _12403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16940__B1 _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15203_ _15203_/A _15203_/B _15203_/C vssd1 vssd1 vccd1 vccd1 _15204_/B sky130_fd_sc_hd__and3_1
X_12415_ _12416_/A _12416_/B _12416_/C vssd1 vssd1 vccd1 vccd1 _12415_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17387__A _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16183_ _16183_/A _16183_/B vssd1 vssd1 vccd1 vccd1 _16185_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_140_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13395_ _13396_/A _13396_/B vssd1 vssd1 vccd1 vccd1 _13395_/X sky130_fd_sc_hd__or2_1
XFILLER_0_112_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15134_ _15133_/B _15271_/B _15133_/A vssd1 vssd1 vccd1 vccd1 _15135_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_106_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12346_ _12346_/A _12346_/B vssd1 vssd1 vccd1 vccd1 _12348_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_49_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11780__A2 _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15065_ _15065_/A _15065_/B vssd1 vssd1 vccd1 vccd1 _15067_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__16441__D _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19942_ _19942_/A _19942_/B _19942_/C vssd1 vssd1 vccd1 vccd1 _19943_/B sky130_fd_sc_hd__and3_1
XFILLER_0_65_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19237__A2 _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ _12241_/X _12275_/X _12276_/Y vssd1 vssd1 vccd1 vccd1 _12277_/X sky130_fd_sc_hd__o21a_1
XANTENNA__14242__C _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14016_ _14015_/B _14015_/C _14015_/A vssd1 vssd1 vccd1 vccd1 _14113_/B sky130_fd_sc_hd__a21oi_1
X_11228_ _12269_/A _11227_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21758_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_120_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19873_ _21833_/Q _19874_/B _19874_/C _19874_/D vssd1 vssd1 vccd1 vccd1 _19873_/Y
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__17834__B _17834_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15635__A _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18824_ _18674_/C _18673_/Y _18822_/X _18823_/Y vssd1 vssd1 vccd1 vccd1 _18826_/C
+ sky130_fd_sc_hd__o211a_1
X_11159_ _12877_/B _11158_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21736_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17553__C _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18755_ _18755_/A _18755_/B vssd1 vssd1 vccd1 vccd1 _18757_/C sky130_fd_sc_hd__xnor2_1
X_15967_ _15966_/A _15966_/B _15966_/C vssd1 vssd1 vccd1 vccd1 _15968_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__18748__A1 _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11374__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13155__A _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17706_ _17705_/A _17705_/B _17830_/A vssd1 vssd1 vccd1 vccd1 _17707_/B sky130_fd_sc_hd__o21a_1
XANTENNA__18748__B2 _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14918_ _15206_/A _14918_/B vssd1 vssd1 vccd1 vccd1 _14918_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__11296__A1 _11295_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18686_ _18686_/A _18686_/B vssd1 vssd1 vccd1 vccd1 _18687_/B sky130_fd_sc_hd__xnor2_4
X_15898_ _16029_/A _15898_/B vssd1 vssd1 vccd1 vccd1 _15899_/B sky130_fd_sc_hd__and2_1
XFILLER_0_72_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17637_ _18008_/A _18008_/B _18616_/D vssd1 vssd1 vccd1 vccd1 _17637_/X sky130_fd_sc_hd__and3_1
X_14849_ _14847_/X _14848_/Y _14418_/A _14418_/B vssd1 vssd1 vccd1 vccd1 _14974_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_72_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13037__A2 _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15431__B1 _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15370__A _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17568_ _17567_/A _17567_/B _17567_/C vssd1 vssd1 vccd1 vccd1 _17570_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_147_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19307_ _19307_/A _19307_/B vssd1 vssd1 vccd1 vccd1 _19308_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__19199__D _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16519_ _17206_/B _17621_/C vssd1 vssd1 vccd1 vccd1 _16522_/A sky130_fd_sc_hd__and2_1
XFILLER_0_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17499_ _18859_/A _21151_/A vssd1 vssd1 vccd1 vccd1 _17500_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19238_ _19692_/A _19906_/A _19238_/C _19692_/B vssd1 vssd1 vccd1 vccd1 _19387_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_6_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11122__B _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19169_ _19788_/A _19169_/B vssd1 vssd1 vccd1 vccd1 _19169_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_103_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21200_ _21200_/A _21287_/A vssd1 vssd1 vccd1 vccd1 _21201_/B sky130_fd_sc_hd__nand2_1
XANTENNA__15529__B _15529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13975__D _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15498__B1 _10941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21131_ _21131_/A _21131_/B vssd1 vssd1 vccd1 vccd1 _21134_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19228__A2 _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17239__A1 _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout403 _21769_/Q vssd1 vssd1 vccd1 vccd1 _15763_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__13049__B _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21062_ _21172_/A _21062_/B vssd1 vssd1 vccd1 vccd1 _21064_/B sky130_fd_sc_hd__xor2_1
XANTENNA__17239__B2 _17557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout414 _21766_/Q vssd1 vssd1 vccd1 vccd1 _12899_/B sky130_fd_sc_hd__clkbuf_8
Xfanout425 _21764_/Q vssd1 vssd1 vccd1 vccd1 _12771_/C sky130_fd_sc_hd__buf_4
XANTENNA_fanout394_A _21771_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout436 _12780_/A vssd1 vssd1 vccd1 vccd1 _12267_/A sky130_fd_sc_hd__buf_4
X_20013_ _20154_/B _20012_/B _20012_/C vssd1 vssd1 vccd1 vccd1 _20014_/C sky130_fd_sc_hd__a21o_1
Xfanout447 _21759_/Q vssd1 vssd1 vccd1 vccd1 _14087_/A sky130_fd_sc_hd__buf_4
Xfanout458 _21755_/Q vssd1 vssd1 vccd1 vccd1 _16177_/B sky130_fd_sc_hd__buf_4
Xfanout469 _21752_/Q vssd1 vssd1 vccd1 vccd1 _14698_/D sky130_fd_sc_hd__buf_4
XANTENNA__20170__B _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15264__B _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout561_A _12621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11284__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18739__A1 _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21964_ _21974_/CLK _21964_/D vssd1 vssd1 vccd1 vccd1 hold266/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__20546__A1 _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20546__B2 _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16214__A2 _16396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20915_ _20916_/A _20916_/B _21033_/A vssd1 vssd1 vccd1 vccd1 _20917_/A sky130_fd_sc_hd__o21ai_2
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21895_ _21932_/CLK _21895_/D vssd1 vssd1 vccd1 vccd1 hold122/A sky130_fd_sc_hd__dfxtp_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15280__A _15281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11039__A1 hold283/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20846_ _20848_/A vssd1 vssd1 vccd1 vccd1 _20983_/A sky130_fd_sc_hd__inv_2
XFILLER_0_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout10 _11547_/X vssd1 vssd1 vccd1 vccd1 _11550_/A sky130_fd_sc_hd__clkbuf_8
Xfanout21 _11224_/Y vssd1 vssd1 vccd1 vccd1 fanout21/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout32 _21481_/S vssd1 vssd1 vccd1 vccd1 _21494_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_64_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout43 _11548_/Y vssd1 vssd1 vccd1 vccd1 _21142_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout54 _11087_/S vssd1 vssd1 vccd1 vccd1 _11088_/S sky130_fd_sc_hd__clkbuf_8
X_20777_ _20910_/A _21171_/B vssd1 vssd1 vccd1 vccd1 _20778_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout65 hold321/X vssd1 vssd1 vccd1 vccd1 _19185_/B sky130_fd_sc_hd__buf_4
XFILLER_0_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout76 _20193_/D vssd1 vssd1 vccd1 vccd1 _21311_/B sky130_fd_sc_hd__buf_4
XFILLER_0_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout87 _19053_/B vssd1 vssd1 vccd1 vccd1 _20671_/B sky130_fd_sc_hd__buf_4
XANTENNA__20048__D _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout98 _21842_/Q vssd1 vssd1 vccd1 vccd1 _21256_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12200_ _12207_/A _12200_/B vssd1 vssd1 vccd1 vccd1 _12203_/B sky130_fd_sc_hd__nand2_1
X_13180_ _14716_/A _14384_/C vssd1 vssd1 vccd1 vccd1 _13184_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15439__B _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12131_ _12127_/B _12127_/C _12127_/A vssd1 vssd1 vccd1 vccd1 _12131_/Y sky130_fd_sc_hd__o21ai_1
X_21329_ _21412_/A _11549_/A _21329_/B1 vssd1 vssd1 vccd1 vccd1 _21329_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_130_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12062_ _12109_/C _12269_/C _12061_/B _12058_/X vssd1 vssd1 vccd1 vccd1 _12063_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11013_ mstream_o[87] hold7/X _11027_/S vssd1 vssd1 vccd1 vccd1 _21624_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18469__C _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16870_ _16870_/A _17013_/D vssd1 vssd1 vccd1 vccd1 _16871_/B sky130_fd_sc_hd__nand2_1
X_15821_ _15683_/B _15683_/Y _15819_/Y _15820_/X vssd1 vssd1 vccd1 vccd1 _15823_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_99_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18540_ hold151/X _18539_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _21897_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17670__A _21824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15752_ _15752_/A _15752_/B vssd1 vssd1 vccd1 vccd1 _15755_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11278__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12964_ _13244_/A _12964_/B vssd1 vssd1 vccd1 vccd1 _12966_/C sky130_fd_sc_hd__or2_1
XTAP_3352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14703_ _14541_/Y _14543_/X _14700_/X _14702_/Y vssd1 vssd1 vccd1 vccd1 _14705_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__21192__A _21293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18471_ _18321_/A _18321_/B _18320_/B vssd1 vssd1 vccd1 vccd1 _18473_/B sky130_fd_sc_hd__o21ai_1
X_11915_ _11914_/B _11914_/C _11914_/A vssd1 vssd1 vccd1 vccd1 _11917_/B sky130_fd_sc_hd__a21bo_1
X_15683_ _15683_/A _15683_/B _15683_/C vssd1 vssd1 vccd1 vccd1 _15683_/Y sky130_fd_sc_hd__nand3_4
XTAP_3385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14216__A1 _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13019__A2 _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16286__A _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_330 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14216__B2 _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ _12895_/A _12895_/B vssd1 vssd1 vccd1 vccd1 _12929_/A sky130_fd_sc_hd__nand2_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17422_ _17423_/A _17423_/B vssd1 vssd1 vccd1 vccd1 _17422_/X sky130_fd_sc_hd__and2_2
X_14634_ _15579_/D _15717_/C _15976_/D _15153_/B vssd1 vssd1 vccd1 vccd1 _14637_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14767__A2 _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11846_ _11845_/B _11845_/C _11845_/A vssd1 vssd1 vccd1 vccd1 _11848_/B sky130_fd_sc_hd__a21bo_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14518__B _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17353_ _17251_/B _17251_/Y _17350_/X _17352_/Y vssd1 vssd1 vccd1 vccd1 _17356_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_32_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14565_ _14712_/A _14712_/B _16380_/B _16173_/B vssd1 vssd1 vccd1 vccd1 _14568_/B
+ sky130_fd_sc_hd__nand4_1
X_11777_ _12297_/B _11776_/B _11776_/C _11776_/D vssd1 vssd1 vccd1 vccd1 _11777_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_56_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12319__A _13554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16304_ _16305_/B _16399_/B _16409_/B _16404_/A vssd1 vssd1 vccd1 vccd1 _16306_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_55_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13516_ hold88/X _13515_/X fanout2/X vssd1 vssd1 vccd1 vccd1 _21864_/D sky130_fd_sc_hd__mux2_1
XANTENNA__11450__A1 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17284_ _17504_/C _17739_/C _17739_/D _17490_/A vssd1 vssd1 vccd1 vccd1 _17285_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11450__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14496_ _14496_/A _14496_/B vssd1 vssd1 vccd1 vccd1 _14588_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_70_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12038__B _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16733__B _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19023_ _19024_/A _19024_/B _19024_/C vssd1 vssd1 vccd1 vccd1 _19023_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16235_ _16235_/A vssd1 vssd1 vccd1 vccd1 _16348_/A sky130_fd_sc_hd__inv_2
X_13447_ _13447_/A _13447_/B vssd1 vssd1 vccd1 vccd1 _13449_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_35_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12980__C _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16166_ _16167_/A _16167_/B vssd1 vssd1 vccd1 vccd1 _16322_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_140_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13378_ _13682_/C _14155_/C _14155_/D _13822_/B vssd1 vssd1 vccd1 vccd1 _13378_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__18130__A2 _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15117_ _16196_/B _16371_/A _16305_/B _15791_/A vssd1 vssd1 vccd1 vccd1 _15120_/C
+ sky130_fd_sc_hd__a22o_1
X_12329_ _12329_/A _12329_/B vssd1 vssd1 vccd1 vccd1 _12332_/A sky130_fd_sc_hd__xnor2_1
X_16097_ _15965_/A _15964_/A _15964_/B _15960_/B _15960_/A vssd1 vssd1 vccd1 vccd1
+ _16098_/B sky130_fd_sc_hd__o32ai_4
XFILLER_0_107_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11596__C _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21367__A _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15048_ _14837_/Y _14839_/X _15046_/Y _15047_/X vssd1 vssd1 vccd1 vccd1 _15050_/C
+ sky130_fd_sc_hd__o211ai_4
X_19925_ _19925_/A _19925_/B vssd1 vssd1 vccd1 vccd1 _19928_/A sky130_fd_sc_hd__and2_1
XFILLER_0_142_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19856_ _19855_/B _19950_/B _20091_/A vssd1 vssd1 vccd1 vccd1 _19857_/C sky130_fd_sc_hd__a21o_1
XANTENNA__17283__C _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18807_ _18807_/A _18807_/B _18807_/C vssd1 vssd1 vccd1 vccd1 _18810_/A sky130_fd_sc_hd__nand3_2
X_19787_ _19476_/A _19787_/B vssd1 vssd1 vccd1 vccd1 _19788_/C sky130_fd_sc_hd__nand2b_1
X_16999_ _16999_/A _16999_/B _16999_/C vssd1 vssd1 vccd1 vccd1 _17000_/B sky130_fd_sc_hd__or3_1
XANTENNA__12501__B _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11269__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18738_ _19531_/A _19051_/A _19227_/C _19057_/D vssd1 vssd1 vccd1 vccd1 _18741_/D
+ sky130_fd_sc_hd__nand4_1
X_18669_ _18669_/A _18669_/B _18669_/C _18669_/D vssd1 vssd1 vccd1 vccd1 _18669_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20700_ _20700_/A vssd1 vssd1 vccd1 vccd1 _20700_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13613__A _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21680_ _21682_/CLK _21680_/D vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20631_ _20628_/X _20629_/X _20499_/A _20499_/Y vssd1 vssd1 vccd1 vccd1 _20631_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_110_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout142_A _21833_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12229__A _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11441__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20562_ _21056_/A _20562_/B _21046_/B _21278_/B vssd1 vssd1 vccd1 vccd1 _20685_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__17739__B _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_17_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21949_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20493_ _20491_/B _20491_/C _20491_/A vssd1 vssd1 vccd1 vccd1 _20493_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout407_A _21768_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21114_ _20998_/Y _21000_/Y _21112_/X _21113_/Y vssd1 vssd1 vccd1 vccd1 _21188_/A
+ sky130_fd_sc_hd__o211a_1
Xfanout200 _21256_/B vssd1 vssd1 vccd1 vccd1 _19972_/C sky130_fd_sc_hd__clkbuf_4
X_22094_ _22105_/CLK _22094_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[30] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12899__A _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14694__A1 _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout211 _19866_/C vssd1 vssd1 vccd1 vccd1 _19414_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout222 _21311_/A vssd1 vssd1 vccd1 vccd1 _20924_/A sky130_fd_sc_hd__buf_4
XFILLER_0_121_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21045_ _21256_/A _21816_/Q _21046_/C _21046_/D vssd1 vssd1 vccd1 vccd1 _21047_/A
+ sky130_fd_sc_hd__a22oi_1
Xfanout233 _17924_/B vssd1 vssd1 vccd1 vccd1 _18773_/B sky130_fd_sc_hd__buf_4
Xfanout244 _21807_/Q vssd1 vssd1 vccd1 vccd1 _19692_/A sky130_fd_sc_hd__clkbuf_4
Xfanout255 _19892_/A vssd1 vssd1 vccd1 vccd1 _20845_/D sky130_fd_sc_hd__buf_4
Xfanout266 _18030_/B vssd1 vssd1 vccd1 vccd1 _19531_/A sky130_fd_sc_hd__clkbuf_4
Xfanout277 _21800_/Q vssd1 vssd1 vccd1 vccd1 _18008_/A sky130_fd_sc_hd__buf_4
Xfanout288 _17619_/A vssd1 vssd1 vccd1 vccd1 _16968_/C sky130_fd_sc_hd__buf_4
Xfanout299 _17621_/C vssd1 vssd1 vccd1 vccd1 _17063_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17490__A _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20519__A1 _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14997__A2 _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20519__B2 _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21947_ _21949_/CLK _21947_/D vssd1 vssd1 vccd1 vccd1 hold189/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__17396__B1 _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ _12318_/A _11699_/C _11699_/A vssd1 vssd1 vccd1 vccd1 _11701_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_16_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ _12679_/A _12679_/B _12679_/C vssd1 vssd1 vccd1 vccd1 _12681_/C sky130_fd_sc_hd__a21o_1
X_21878_ _21945_/CLK _21878_/D vssd1 vssd1 vccd1 vccd1 hold263/A sky130_fd_sc_hd__dfxtp_1
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _12109_/C _12528_/B _11630_/C _11683_/A vssd1 vssd1 vccd1 vccd1 _11631_/X
+ sky130_fd_sc_hd__a22o_1
X_20829_ _20826_/Y _20827_/X _20699_/B _20700_/Y vssd1 vssd1 vccd1 vccd1 _20830_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14350_ _15153_/B _15788_/B vssd1 vssd1 vccd1 vccd1 _14351_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_92_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11432__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11562_ _12109_/C _12619_/A vssd1 vssd1 vccd1 vccd1 _11566_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13709__B1 _14663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13301_ _13302_/A _13302_/B vssd1 vssd1 vccd1 vccd1 _13301_/X sky130_fd_sc_hd__and2_2
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14281_ _14282_/A _14282_/B vssd1 vssd1 vccd1 vccd1 _14446_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_18_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11493_ _11493_/A1 t2x[14] v1z[14] fanout20/X _11492_/X vssd1 vssd1 vccd1 vccd1 _11493_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__14354__A _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16020_ _16016_/X _16018_/Y _16019_/X vssd1 vssd1 vccd1 vccd1 _16021_/C sky130_fd_sc_hd__o21a_1
X_13232_ _13822_/B _13997_/C _13115_/B _13113_/X vssd1 vssd1 vccd1 vccd1 _13237_/A
+ sky130_fd_sc_hd__a31oi_2
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11189__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13163_ _13287_/A _13162_/C _13162_/A vssd1 vssd1 vccd1 vccd1 _13164_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_21_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14134__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12114_ _12115_/A _12115_/B _12115_/C vssd1 vssd1 vccd1 vccd1 _12114_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__17871__A1 _18008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13094_ _16363_/A hold155/A _11059_/Y fanout6/X _13093_/Y vssd1 vssd1 vccd1 vccd1
+ _13094_/X sky130_fd_sc_hd__a221o_1
X_17971_ _21142_/A _21352_/B vssd1 vssd1 vccd1 vccd1 _17971_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17384__B _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17871__B2 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19710_ _19551_/A _19551_/C _19551_/B vssd1 vssd1 vccd1 vccd1 _19711_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_100_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11499__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16922_ _16863_/A _16863_/C _16863_/B vssd1 vssd1 vccd1 vccd1 _16923_/C sky130_fd_sc_hd__a21o_1
X_12045_ _12094_/A _12530_/A _12512_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _12046_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11499__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19641_ _19522_/A _19522_/B _19520_/Y vssd1 vssd1 vccd1 vccd1 _19683_/A sky130_fd_sc_hd__o21ba_1
X_16853_ _16851_/A _16859_/A _16852_/Y _16785_/X vssd1 vssd1 vccd1 vccd1 _17165_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_102_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15804_ _15931_/B _16391_/B _16369_/B _15931_/A vssd1 vssd1 vccd1 vccd1 _15808_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19572_ _19575_/D vssd1 vssd1 vccd1 vccd1 _19572_/Y sky130_fd_sc_hd__inv_2
X_16784_ _16789_/A _16784_/B vssd1 vssd1 vccd1 vccd1 _16785_/C sky130_fd_sc_hd__nor2_1
X_13996_ _13858_/B _13997_/C _14155_/C _14936_/D vssd1 vssd1 vccd1 vccd1 _13999_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18523_ _18373_/C _18372_/Y _18521_/X _18522_/Y vssd1 vssd1 vccd1 vccd1 _18525_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15632__B _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15735_ _15563_/Y _15567_/B _15733_/X _15734_/Y vssd1 vssd1 vccd1 vccd1 _15737_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_133_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11120__A0 _10984_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12947_ _12947_/A _12947_/B _12947_/C vssd1 vssd1 vccd1 vccd1 _12950_/C sky130_fd_sc_hd__and3_1
XTAP_3182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17926__A2 _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18454_ _18454_/A _18454_/B _18441_/X vssd1 vssd1 vccd1 vccd1 _18454_/Y sky130_fd_sc_hd__nor3b_4
X_15666_ _15667_/A _15667_/B vssd1 vssd1 vccd1 vccd1 _15862_/B sky130_fd_sc_hd__or2_1
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ _12877_/A _13152_/C _13152_/D _12877_/B vssd1 vssd1 vccd1 vccd1 _12878_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA_160 v2z[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14248__B _21759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_171 v2z[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17405_ _17405_/A _17405_/B _17405_/C vssd1 vssd1 vccd1 vccd1 _17405_/Y sky130_fd_sc_hd__nor3_2
XANTENNA_182 v2z[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_193 hold247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14617_ _14774_/D _15698_/B vssd1 vssd1 vccd1 vccd1 _14618_/B sky130_fd_sc_hd__nand2_2
XANTENNA__13152__B _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18385_ _18385_/A _18385_/B vssd1 vssd1 vccd1 vccd1 _18388_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_28_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11829_ _11833_/B _11830_/B _11830_/C _11830_/D vssd1 vssd1 vccd1 vccd1 _11829_/X
+ sky130_fd_sc_hd__and4_1
X_15597_ _15598_/A _15598_/B vssd1 vssd1 vccd1 vccd1 _15597_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16744__A _21830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17336_ _17336_/A _17336_/B vssd1 vssd1 vccd1 vccd1 _17345_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11423__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14548_ _14548_/A _14690_/B _14548_/C vssd1 vssd1 vccd1 vccd1 _14551_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12620__B1 _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12991__B _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18351__A2 _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17267_ _17267_/A _17267_/B vssd1 vssd1 vccd1 vccd1 _17379_/B sky130_fd_sc_hd__xnor2_4
X_14479_ _15159_/D _15174_/D _14479_/C _14632_/A vssd1 vssd1 vccd1 vccd1 _14632_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_70_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19006_ _19006_/A _19006_/B vssd1 vssd1 vccd1 vccd1 _19048_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_52_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16218_ _16409_/A _16328_/B _16218_/C _16218_/D vssd1 vssd1 vccd1 vccd1 _16323_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__15079__B _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20416__D _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17198_ _17198_/A _17198_/B vssd1 vssd1 vccd1 vccd1 _17260_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18103__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11726__A2 _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16149_ _16029_/A _16029_/B _15764_/B vssd1 vssd1 vccd1 vccd1 _16150_/B sky130_fd_sc_hd__o21ai_4
XFILLER_0_140_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19493__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19851__A2 _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17862__A1 _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17862__B2 _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19908_ _20148_/C _20273_/A _19908_/C _20001_/A vssd1 vssd1 vccd1 vccd1 _20001_/B
+ sky130_fd_sc_hd__nand4_2
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12512__A _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16417__A2 _21784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12151__A2 _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19839_ _19840_/A _19840_/B vssd1 vssd1 vccd1 vccd1 _19839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_39_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_127_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21801_ _21803_/CLK _21801_/D vssd1 vssd1 vccd1 vccd1 _21801_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_79_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18556__D _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11111__A0 _10926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout357_A _16391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21732_ _21803_/CLK _21732_/D vssd1 vssd1 vccd1 vccd1 _21732_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15928__A1 _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20921__A1 _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20921__B2 _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21663_ _21906_/CLK _21663_/D vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_143_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13403__A2 hold241/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_359 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20614_ _20616_/A _20616_/B _20616_/C vssd1 vssd1 vccd1 vccd1 _20614_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11414__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13997__B _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21594_ _21888_/CLK _21594_/D _11041_/A vssd1 vssd1 vccd1 vccd1 mstream_o[57] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_145_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12109__D _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20545_ _20545_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20556_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_105_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16092__C hold319/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14364__B1 _21744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20476_ _21261_/A _20838_/B _21283_/B _21305_/B vssd1 vssd1 vccd1 vccd1 _20602_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_61_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17302__B1 _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17730__A2_N _19060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14621__B _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22077_ _22080_/CLK _22077_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[13] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12142__A2 _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21028_ _21142_/A _21412_/B vssd1 vssd1 vccd1 vccd1 _21028_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__21401__A2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15155__D _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13850_ _13847_/Y _13848_/X _13689_/Y _13692_/X vssd1 vssd1 vccd1 vccd1 _13851_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12801_ _12797_/X _12799_/Y _12687_/B _12687_/Y vssd1 vssd1 vccd1 vccd1 _12803_/D
+ sky130_fd_sc_hd__o211a_2
XANTENNA__11102__A0 _10860_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13781_ _13627_/A _13627_/C _13627_/B vssd1 vssd1 vccd1 vccd1 _13782_/C sky130_fd_sc_hd__a21bo_1
X_10993_ mstream_o[67] hold11/X _11005_/S vssd1 vssd1 vccd1 vccd1 _21604_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_69_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15520_ _16031_/A _15521_/B vssd1 vssd1 vccd1 vccd1 _15520_/X sky130_fd_sc_hd__and2_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ _12732_/A _12732_/B vssd1 vssd1 vccd1 vccd1 _12741_/A sky130_fd_sc_hd__or2_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15451_ _15451_/A _15451_/B vssd1 vssd1 vccd1 vccd1 _15459_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ _12663_/A _12663_/B vssd1 vssd1 vccd1 vccd1 _12665_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_38_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14402_ _14402_/A _14402_/B vssd1 vssd1 vccd1 vccd1 _14427_/A sky130_fd_sc_hd__and2_2
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18170_ _19535_/A _18319_/B _18622_/B _19695_/A vssd1 vssd1 vccd1 vccd1 _18170_/Y
+ sky130_fd_sc_hd__a22oi_1
X_11614_ _11897_/A _11897_/B vssd1 vssd1 vccd1 vccd1 _11623_/A sky130_fd_sc_hd__or2_1
XANTENNA__11405__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15382_ _15382_/A _15382_/B vssd1 vssd1 vccd1 vccd1 _15384_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_38_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12602__B1 _11051_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12594_ _12481_/Y _12484_/X _12592_/X _12593_/Y vssd1 vssd1 vccd1 vccd1 _12831_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__18333__A2 _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19530__A1 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17121_ _17099_/A _17099_/C _17099_/B vssd1 vssd1 vccd1 vccd1 _17134_/B sky130_fd_sc_hd__a21o_1
X_14333_ _14322_/Y _14333_/B _14333_/C vssd1 vssd1 vccd1 vccd1 _14489_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11545_ _11544_/X _20721_/C _11545_/S vssd1 vssd1 vccd1 vccd1 _21853_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_151_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14084__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13158__A1 _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17052_ _17144_/A _17129_/B _17124_/C _17145_/B vssd1 vssd1 vccd1 vccd1 _17052_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_29_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14264_ _14264_/A _14264_/B _14264_/C vssd1 vssd1 vccd1 vccd1 _14264_/Y sky130_fd_sc_hd__nand3_2
X_11476_ _11475_/X _18789_/A _11521_/S vssd1 vssd1 vccd1 vccd1 _21830_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_151_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11169__B1 fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16003_ _15870_/Y _15874_/C _16001_/X _16002_/Y vssd1 vssd1 vccd1 vccd1 _16003_/Y
+ sky130_fd_sc_hd__o211ai_4
X_13215_ _13074_/X _13077_/X _13213_/Y _13214_/X vssd1 vssd1 vccd1 vccd1 _13218_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__17395__A _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14195_ _14195_/A _16286_/A _14195_/C _14362_/A vssd1 vssd1 vccd1 vccd1 _14362_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_110_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17844__A1 _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13146_ _13002_/B _13003_/Y _13230_/A _13145_/X vssd1 vssd1 vccd1 vccd1 _13230_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13077_ _13077_/A _13077_/B _13077_/C vssd1 vssd1 vccd1 vccd1 _13077_/X sky130_fd_sc_hd__and3_2
X_17954_ _17953_/B _17953_/C _17953_/A vssd1 vssd1 vccd1 vccd1 _17954_/Y sky130_fd_sc_hd__o21ai_2
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16905_ _16903_/A _16958_/A _16904_/X _16843_/Y vssd1 vssd1 vccd1 vccd1 _16909_/A
+ sky130_fd_sc_hd__a211o_1
X_12028_ _12029_/A _12029_/B _12029_/C vssd1 vssd1 vccd1 vccd1 _12286_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_40_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17885_ _17883_/B _17883_/C _17883_/A vssd1 vssd1 vccd1 vccd1 _17885_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__15643__A _16031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16836_ _16836_/A _16836_/B vssd1 vssd1 vccd1 vccd1 _16894_/B sky130_fd_sc_hd__xor2_1
X_19624_ _19624_/A _19624_/B vssd1 vssd1 vccd1 vccd1 _19626_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__21364__B _21364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19349__A1 _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16458__B _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19349__B2 fanout96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19555_ _19554_/A _19554_/B _19554_/C vssd1 vssd1 vccd1 vccd1 _19556_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_88_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13094__B1 _11059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16767_ _16767_/A vssd1 vssd1 vccd1 vccd1 _16769_/A sky130_fd_sc_hd__inv_2
X_13979_ _13979_/A _13979_/B vssd1 vssd1 vccd1 vccd1 _13981_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_88_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18506_ _18505_/B _18505_/C _18505_/A vssd1 vssd1 vccd1 vccd1 _18508_/B sky130_fd_sc_hd__a21o_1
X_15718_ _16087_/A _15978_/B _15716_/Y _15848_/A vssd1 vssd1 vccd1 vccd1 _15720_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_19486_ _19487_/A _20838_/C _20838_/D _19487_/B vssd1 vssd1 vccd1 vccd1 _19486_/X
+ sky130_fd_sc_hd__a22o_1
X_16698_ _16698_/A _16698_/B _16698_/C vssd1 vssd1 vccd1 vccd1 _16741_/A sky130_fd_sc_hd__nand3_2
X_18437_ _18438_/A _18438_/B vssd1 vssd1 vccd1 vccd1 _18564_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15649_ _15907_/A _15648_/B _15648_/C vssd1 vssd1 vccd1 vccd1 _15650_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_111_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18368_ _18368_/A _18368_/B _18368_/C _18368_/D vssd1 vssd1 vccd1 vccd1 _18368_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_127_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17319_ _17212_/X _17214_/X _17316_/X _17317_/Y vssd1 vssd1 vccd1 vccd1 _17319_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11947__A2 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18299_ _18296_/X _18442_/B _18167_/D _18169_/A vssd1 vssd1 vccd1 vccd1 _18300_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_154_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20330_ _20330_/A _20330_/B vssd1 vssd1 vccd1 vccd1 _20338_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20146__D _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20261_ _20259_/Y _20260_/X _20096_/Y _20120_/Y vssd1 vssd1 vccd1 vccd1 _20302_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_12_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout105_A _19691_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19824__A2 _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22000_ _22005_/CLK _22000_/D vssd1 vssd1 vccd1 vccd1 hold162/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_40_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16638__A2 _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20192_ _20721_/D _20193_/D _20190_/Y _20329_/A vssd1 vssd1 vccd1 vccd1 _20194_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__13983__D _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12242__A _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19951__C _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13321__A1 _14712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13321__B2 _14712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11332__A0 _15174_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13872__A2 _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout474_A _15093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15074__A1 _14968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11292__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21715_ _22105_/CLK _21715_/D vssd1 vssd1 vccd1 vccd1 hold67/A sky130_fd_sc_hd__dfxtp_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16574__A1 _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16574__B2 _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21646_ _21722_/CLK _21646_/D fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[109]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout18_A fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18315__A2 _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12060__A1 _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19695__A _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15129__A2 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12060__B2 _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21577_ mstream_o[40] _11061_/X _21579_/S vssd1 vssd1 vccd1 vccd1 _22104_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_60 hold270/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_71 hold268/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_82 hold234/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _11544_/A1 t1x[26] v2z[26] _11223_/A _11329_/X vssd1 vssd1 vccd1 vccd1 _11330_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_144_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_93 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16877__A2 _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20528_ _20528_/A _20686_/B _20529_/B vssd1 vssd1 vccd1 vccd1 _20651_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_133_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11261_ _11325_/A1 t2y[9] t0y[9] _11498_/A1 vssd1 vssd1 vccd1 vccd1 _11261_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20459_ _20459_/A _20588_/B vssd1 vssd1 vccd1 vccd1 _20461_/A sky130_fd_sc_hd__or2_2
XFILLER_0_127_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13000_ _13000_/A _13000_/B _13000_/C vssd1 vssd1 vccd1 vccd1 _13002_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_24_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11192_ _14384_/D _11191_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21747_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_24_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11467__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14951_ _15579_/D _15174_/D _14951_/C _15169_/A vssd1 vssd1 vccd1 vccd1 _15169_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__20189__A2 _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11323__B1 _11322_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13902_ _13750_/D _13751_/B _13900_/Y _13901_/X vssd1 vssd1 vccd1 vccd1 _14051_/A
+ sky130_fd_sc_hd__a211o_1
X_17670_ _21824_/Q _17670_/B vssd1 vssd1 vccd1 vccd1 _17673_/A sky130_fd_sc_hd__and2_1
X_14882_ _14881_/B _14881_/C _14881_/A vssd1 vssd1 vccd1 vccd1 _14883_/C sky130_fd_sc_hd__a21o_1
X_16621_ _17146_/A _17334_/B _18166_/A _17146_/B vssd1 vssd1 vccd1 vccd1 _16622_/C
+ sky130_fd_sc_hd__a22o_1
X_13833_ _13833_/A _13833_/B vssd1 vssd1 vccd1 vccd1 _13834_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19340_ _19340_/A _19340_/B vssd1 vssd1 vccd1 vccd1 _19341_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_74_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16552_ _16552_/A _16552_/B vssd1 vssd1 vccd1 vccd1 _16553_/B sky130_fd_sc_hd__xnor2_1
X_13764_ _14557_/A _14557_/B _14873_/B _13913_/C vssd1 vssd1 vccd1 vccd1 _13910_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_85_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10976_ hold128/A hold146/A vssd1 vssd1 vccd1 vccd1 _10977_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_84_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15503_ _15907_/A _16261_/B vssd1 vssd1 vccd1 vccd1 _16151_/A sky130_fd_sc_hd__nor2_2
X_19271_ _19271_/A _19406_/B _19271_/C vssd1 vssd1 vccd1 vccd1 _19271_/Y sky130_fd_sc_hd__nand3_1
X_12715_ _12716_/A _12716_/B _12716_/C vssd1 vssd1 vccd1 vccd1 _12942_/A sky130_fd_sc_hd__a21oi_2
X_16483_ _17206_/B _17141_/C _16482_/B _16479_/X vssd1 vssd1 vccd1 vccd1 _16485_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13695_ _13698_/B vssd1 vssd1 vccd1 vccd1 _13695_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_84_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18222_ _18082_/B _18081_/Y _18220_/X _18221_/Y vssd1 vssd1 vccd1 vccd1 _18225_/B
+ sky130_fd_sc_hd__o211a_2
X_15434_ _15435_/A _15698_/B _15435_/C _15435_/D vssd1 vssd1 vccd1 vccd1 _15436_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_72_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17622__A2_N _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12646_ _12646_/A _12646_/B vssd1 vssd1 vccd1 vccd1 _12649_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18153_ _18304_/A _18152_/C _18152_/A vssd1 vssd1 vccd1 vccd1 _18155_/B sky130_fd_sc_hd__a21o_1
XANTENNA__20247__C _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15365_ _15365_/A _15365_/B vssd1 vssd1 vccd1 vccd1 _15386_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_142_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12577_ _12578_/A _12578_/B _12578_/C vssd1 vssd1 vccd1 vccd1 _12577_/X sky130_fd_sc_hd__and3_1
XFILLER_0_142_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17104_ _17110_/A _17104_/B vssd1 vssd1 vccd1 vccd1 _17106_/B sky130_fd_sc_hd__or2_1
X_14316_ _14316_/A _14316_/B vssd1 vssd1 vccd1 vccd1 _14317_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18084_ _17948_/B _17947_/Y _18082_/X _18083_/Y vssd1 vssd1 vccd1 vccd1 _18087_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_13_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11528_ _21723_/D t1y[26] t0x[26] _11223_/A vssd1 vssd1 vccd1 vccd1 _11528_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_40_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15296_ _15296_/A _15296_/B vssd1 vssd1 vccd1 vccd1 _15297_/A sky130_fd_sc_hd__or2_1
XFILLER_0_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20544__A _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold308 hold308/A vssd1 vssd1 vccd1 vccd1 hold308/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17035_ _17035_/A _17035_/B vssd1 vssd1 vccd1 vccd1 _17036_/B sky130_fd_sc_hd__xnor2_1
Xhold319 hold319/A vssd1 vssd1 vccd1 vccd1 hold319/X sky130_fd_sc_hd__dlygate4sd3_1
X_14247_ _14248_/A _21759_/Q vssd1 vssd1 vccd1 vccd1 _14251_/A sky130_fd_sc_hd__or2_1
XFILLER_0_150_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11459_ _11123_/A t1y[3] t0x[3] _11459_/B2 vssd1 vssd1 vccd1 vccd1 _11459_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_111_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16460__C _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14178_ _15155_/C _16377_/A vssd1 vssd1 vccd1 vccd1 _14179_/B sky130_fd_sc_hd__nand2_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15828__B1 _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11377__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13129_ _13867_/A _15768_/A _13014_/X _13013_/X _13152_/C vssd1 vssd1 vccd1 vccd1
+ _13134_/A sky130_fd_sc_hd__a32o_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15076__C _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18986_ _18983_/X _18984_/X _18822_/C _18821_/Y vssd1 vssd1 vccd1 vccd1 _18986_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17937_ _17937_/A _17937_/B _17937_/C vssd1 vssd1 vccd1 vccd1 _17940_/A sky130_fd_sc_hd__nand3_2
XANTENNA__15373__A _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18242__A1 _17967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17868_ _17869_/A _17869_/B vssd1 vssd1 vccd1 vccd1 _17982_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_84_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19607_ _19606_/B _19606_/C _19606_/A vssd1 vssd1 vccd1 vccd1 _19608_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_75_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16819_ _16820_/A _16820_/B vssd1 vssd1 vccd1 vccd1 _16840_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16619__D _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17799_ _17799_/A _17799_/B _17799_/C vssd1 vssd1 vccd1 vccd1 _17802_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_36_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19538_ _19686_/A _20419_/A _19538_/C _19538_/D vssd1 vssd1 vccd1 vccd1 _19538_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19469_ _19469_/A _19469_/B vssd1 vssd1 vccd1 vccd1 _19472_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__16556__A1 _21825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16556__B2 _16734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21500_ hold292/X sstream_i[77] _21510_/S vssd1 vssd1 vccd1 vccd1 _22027_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_9_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12882__D _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21431_ hold248/X sstream_i[8] _21442_/S vssd1 vssd1 vccd1 vccd1 _21958_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout222_A _21311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14155__C _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21362_ _21412_/A _18390_/Y _21421_/S _21361_/Y vssd1 vssd1 vccd1 vccd1 _21362_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20313_ _20313_/A _20460_/B vssd1 vssd1 vccd1 vccd1 _20316_/A sky130_fd_sc_hd__or2_1
XFILLER_0_141_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21293_ _21293_/A _21293_/B vssd1 vssd1 vccd1 vccd1 _21294_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_114_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20173__B _20841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20244_ _20910_/A _21046_/B _20244_/C _20428_/A vssd1 vssd1 vccd1 vccd1 _20428_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_130_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout591_A _11549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11553__B1 _21329_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18859__A _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17284__A2 _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17763__A _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20175_ _20175_/A _20175_/B vssd1 vssd1 vccd1 vccd1 _20177_/B sky130_fd_sc_hd__or2_1
XFILLER_0_122_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12403__C _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21368__A1 _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18297__C _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16529__D _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17992__B1 _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10830_ _10830_/A _10830_/B vssd1 vssd1 vccd1 vccd1 _11045_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_95_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_156_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19733__A1 _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12500_ _12414_/A _12414_/B _12412_/X vssd1 vssd1 vccd1 vccd1 _12526_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13480_ _13480_/A _13480_/B _13480_/C vssd1 vssd1 vccd1 vccd1 _13483_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_81_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14022__A2 _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12431_ _12528_/B _12426_/B _12328_/B _12326_/X vssd1 vssd1 vccd1 vccd1 _12433_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21629_ _21682_/CLK _21629_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[92] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15150_ _15147_/X _15148_/X _15013_/X _15050_/X vssd1 vssd1 vccd1 vccd1 _15151_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_23_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12362_ _12362_/A _12362_/B _12362_/C vssd1 vssd1 vccd1 vccd1 _12364_/B sky130_fd_sc_hd__nand3_2
XANTENNA__17657__B _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16561__B _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14101_ _14101_/A _14101_/B _14101_/C vssd1 vssd1 vccd1 vccd1 _14101_/Y sky130_fd_sc_hd__nand3_2
X_11313_ _11349_/A1 t2y[22] t0y[22] _21723_/D vssd1 vssd1 vccd1 vccd1 _11313_/X sky130_fd_sc_hd__a22o_1
X_15081_ _15080_/B _15215_/B _15218_/A vssd1 vssd1 vccd1 vccd1 _15082_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_120_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12293_ hold212/X _12292_/X fanout3/X vssd1 vssd1 vccd1 vccd1 _21854_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_120_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14032_ _14032_/A _14032_/B vssd1 vssd1 vccd1 vccd1 _14040_/A sky130_fd_sc_hd__nand2_1
X_11244_ _12242_/B _11243_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21762_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19872__B _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18769__A _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18840_ _18537_/A _18839_/Y _18838_/Y vssd1 vssd1 vccd1 vccd1 _18841_/B sky130_fd_sc_hd__o21ba_2
X_11175_ hold282/X fanout51/X fanout47/X hold285/A vssd1 vssd1 vccd1 vccd1 _11175_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18771_ _19092_/B _19546_/D _19906_/C _19972_/A vssd1 vssd1 vccd1 vccd1 _18775_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15983_ _15983_/A _15983_/B vssd1 vssd1 vccd1 vccd1 _15986_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21359__A1 _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13836__A2 _14477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17722_ _17723_/B vssd1 vssd1 vccd1 vccd1 _17722_/Y sky130_fd_sc_hd__inv_2
X_14934_ _14934_/A _14934_/B _14934_/C vssd1 vssd1 vccd1 vccd1 _14935_/B sky130_fd_sc_hd__and3_1
XANTENNA__12610__A _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17653_ _17531_/X _17533_/X _17651_/X _17652_/Y vssd1 vssd1 vccd1 vccd1 _17689_/A
+ sky130_fd_sc_hd__o211a_1
X_14865_ _14865_/A _14865_/B _14865_/C _14865_/D vssd1 vssd1 vccd1 vccd1 _14868_/B
+ sky130_fd_sc_hd__nand4_1
X_16604_ _16604_/A _16604_/B vssd1 vssd1 vccd1 vccd1 _16617_/A sky130_fd_sc_hd__xnor2_2
X_13816_ _16363_/A hold150/A _10860_/Y fanout5/X _13815_/Y vssd1 vssd1 vccd1 vccd1
+ _13816_/X sky130_fd_sc_hd__a221o_1
X_17584_ _17584_/A _17584_/B _17584_/C vssd1 vssd1 vccd1 vccd1 _17586_/A sky130_fd_sc_hd__and3_1
X_14796_ _14795_/B _14795_/C _14784_/Y vssd1 vssd1 vccd1 vccd1 _14796_/Y sky130_fd_sc_hd__a21boi_1
X_19323_ hold57/A fanout7/X _14449_/B _19636_/A vssd1 vssd1 vccd1 vccd1 _19323_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_35_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16535_ _16468_/A _16468_/B _16475_/X vssd1 vssd1 vccd1 vccd1 _16680_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13747_ _15514_/B _14212_/C _14212_/D _15514_/A vssd1 vssd1 vccd1 vccd1 _13750_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10959_ _10959_/A _10959_/B vssd1 vssd1 vccd1 vccd1 _10959_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_128_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14537__A _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19254_ _19254_/A _19254_/B vssd1 vssd1 vccd1 vccd1 _19304_/A sky130_fd_sc_hd__nor2_1
X_16466_ _16463_/X _16466_/B vssd1 vssd1 vccd1 vccd1 _16478_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_156_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13678_ _13678_/A _13678_/B vssd1 vssd1 vccd1 vccd1 _13687_/A sky130_fd_sc_hd__or2_1
XFILLER_0_155_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18205_ _18204_/B _18204_/C _18204_/A vssd1 vssd1 vccd1 vccd1 _18207_/B sky130_fd_sc_hd__a21o_1
XANTENNA__18951__B _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15417_ _15417_/A _15417_/B vssd1 vssd1 vccd1 vccd1 _15419_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_128_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19185_ _17854_/B _19185_/B _20721_/C _19185_/D vssd1 vssd1 vccd1 vccd1 _19188_/A
+ sky130_fd_sc_hd__and4b_2
X_12629_ _12629_/A _12629_/B _12629_/C vssd1 vssd1 vccd1 vccd1 _12630_/C sky130_fd_sc_hd__nand3_1
X_16397_ _16341_/A _16340_/B _16340_/A vssd1 vssd1 vccd1 vccd1 _16398_/B sky130_fd_sc_hd__o21ba_1
XANTENNA__13772__A1 _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18136_ _19487_/A _19227_/C _19227_/D _19487_/B vssd1 vssd1 vccd1 vccd1 _18137_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13772__B2 _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15348_ _15196_/A _15196_/B _15194_/Y vssd1 vssd1 vccd1 vccd1 _15350_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_79_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15368__A _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold105 hold105/A vssd1 vssd1 vccd1 vccd1 hold105/X sky130_fd_sc_hd__dlygate4sd3_1
X_18067_ _18066_/B _18066_/C _18066_/A vssd1 vssd1 vccd1 vccd1 _18069_/B sky130_fd_sc_hd__a21o_1
X_15279_ _15279_/A _15279_/B vssd1 vssd1 vccd1 vccd1 _15281_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_124_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold116 hold116/A vssd1 vssd1 vccd1 vccd1 hold116/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold127 hold127/A vssd1 vssd1 vccd1 vccd1 hold127/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 hold138/A vssd1 vssd1 vccd1 vccd1 hold138/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13524__A1 _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17018_ _17018_/A _17018_/B _17018_/C vssd1 vssd1 vccd1 vccd1 _17025_/A sky130_fd_sc_hd__nand3_1
Xhold149 hold149/A vssd1 vssd1 vccd1 vccd1 hold149/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12327__A2 _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13524__B2 _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12504__B _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18463__A1 _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout607 _21718_/Q vssd1 vssd1 vccd1 vccd1 _11123_/A sky130_fd_sc_hd__clkbuf_8
Xfanout618 _21717_/Q vssd1 vssd1 vccd1 vccd1 _11012_/S sky130_fd_sc_hd__clkbuf_4
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout629 _17657_/A vssd1 vssd1 vccd1 vccd1 _21087_/D sky130_fd_sc_hd__clkbuf_8
XANTENNA__20721__B _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13288__B1 _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18969_ _18969_/A _18969_/B _18969_/C vssd1 vssd1 vccd1 vccd1 _18972_/A sky130_fd_sc_hd__nand3_2
XANTENNA__16199__A _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21980_ _22013_/CLK _21980_/D vssd1 vssd1 vccd1 vccd1 hold120/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__18766__A2 _19087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20931_ _20931_/A _20931_/B vssd1 vssd1 vccd1 vccd1 _20931_/X sky130_fd_sc_hd__or2_1
XANTENNA_fanout172_A _21827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16927__A _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20862_ _20863_/C _21311_/B _20860_/Y _20985_/A vssd1 vssd1 vccd1 vccd1 _20864_/A
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18445__A1_N _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12263__A1 _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20793_ _21286_/A _21264_/A _20794_/C _20986_/A vssd1 vssd1 vccd1 vccd1 _20795_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout437_A _21761_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16084__D _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17758__A _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout604_A _11459_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13763__A1 _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12566__A2 _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21621__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21414_ hold77/X fanout40/X _21413_/X vssd1 vssd1 vccd1 vccd1 _21946_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_72_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13763__B2 _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15278__A _15279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21345_ hold60/X _21381_/B _21344_/X vssd1 vssd1 vccd1 vccd1 _21922_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_102_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16812__D _17086_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14182__A _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13515__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13515__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21276_ _21206_/A _21205_/Y _21203_/X vssd1 vssd1 vccd1 vccd1 _21277_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17493__A _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20227_ _20372_/A _20083_/B _20079_/A vssd1 vssd1 vccd1 vccd1 _20228_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_21_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16465__B1 _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout85_A _19053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20158_ _20159_/A _20159_/B vssd1 vssd1 vccd1 vccd1 _20307_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_99_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12980_ _14306_/A _14138_/A _13258_/C _13258_/D vssd1 vssd1 vccd1 vccd1 _12980_/X
+ sky130_fd_sc_hd__and4_1
X_20089_ _20089_/A _20089_/B vssd1 vssd1 vccd1 vccd1 _20091_/B sky130_fd_sc_hd__xnor2_2
XTAP_3501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21210__B1 _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19954__A1 _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11931_ _12109_/C _12403_/B vssd1 vssd1 vccd1 vccd1 _12001_/A sky130_fd_sc_hd__nand2_1
XTAP_3545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14650_ _14650_/A _14650_/B vssd1 vssd1 vccd1 vccd1 _14652_/B sky130_fd_sc_hd__xnor2_4
XTAP_3589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11862_ _11859_/X _11862_/B vssd1 vssd1 vccd1 vccd1 _11936_/B sky130_fd_sc_hd__and2b_1
XTAP_2855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13601_ _13602_/A _13602_/B vssd1 vssd1 vccd1 vccd1 _13601_/X sky130_fd_sc_hd__or2_1
XFILLER_0_138_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10813_ hold221/A hold80/A vssd1 vssd1 vccd1 vccd1 _10815_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14581_ _14427_/A _14427_/B _14425_/X vssd1 vssd1 vccd1 vccd1 _14583_/B sky130_fd_sc_hd__a21o_2
XTAP_2888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14357__A _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11793_ _11793_/A _11793_/B vssd1 vssd1 vccd1 vccd1 _11795_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_67_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16320_ _16321_/B vssd1 vssd1 vccd1 vccd1 _16320_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_95_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13532_ _13404_/D _13405_/B _13530_/X _13678_/B vssd1 vssd1 vccd1 vccd1 _13534_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_39_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16251_ _16251_/A _16251_/B vssd1 vssd1 vccd1 vccd1 _16253_/B sky130_fd_sc_hd__or2_1
XANTENNA__12006__A1 _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13463_ _13464_/B _13464_/A vssd1 vssd1 vccd1 vccd1 _13605_/A sky130_fd_sc_hd__and2b_1
XANTENNA__12006__B2 _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16940__A1 _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16940__B2 _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19586__C _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15202_ _15203_/A _15203_/B _15203_/C vssd1 vssd1 vccd1 vccd1 _15204_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_36_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12414_ _12414_/A _12414_/B vssd1 vssd1 vccd1 vccd1 _12416_/C sky130_fd_sc_hd__xnor2_1
X_16182_ _16067_/A _16067_/B _16064_/X vssd1 vssd1 vccd1 vccd1 _16183_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13394_ _13394_/A _16399_/B vssd1 vssd1 vccd1 vccd1 _13396_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17387__B _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15133_ _15133_/A _15133_/B _15271_/B vssd1 vssd1 vccd1 vccd1 _15282_/A sky130_fd_sc_hd__or3_2
XANTENNA__12962__C1 _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12345_ _12343_/X _12345_/B vssd1 vssd1 vccd1 vccd1 _12346_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_23_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15064_ _15065_/A _15065_/B vssd1 vssd1 vccd1 vccd1 _15203_/B sky130_fd_sc_hd__nand2_1
X_19941_ _19941_/A vssd1 vssd1 vccd1 vccd1 _19943_/A sky130_fd_sc_hd__inv_2
XANTENNA__15932__A2_N _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12276_ _12258_/A _12258_/C _12258_/B vssd1 vssd1 vccd1 vccd1 _12276_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14015_ _14015_/A _14015_/B _14015_/C vssd1 vssd1 vccd1 vccd1 _14113_/A sky130_fd_sc_hd__and3_1
XANTENNA__15916__A _16380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11227_ fanout59/X v0z[0] fanout19/X _11226_/X vssd1 vssd1 vccd1 vccd1 _11227_/X
+ sky130_fd_sc_hd__a31o_1
X_19872_ _19972_/A _20394_/B _19872_/C _19972_/C vssd1 vssd1 vccd1 vccd1 _19874_/D
+ sky130_fd_sc_hd__nand4_1
XANTENNA__14820__A _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18823_ _18822_/A _18822_/B _18822_/C _18822_/D vssd1 vssd1 vccd1 vccd1 _18823_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_156_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15635__B _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158_ hold210/X fanout23/X _11157_/X vssd1 vssd1 vccd1 vccd1 _11158_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13436__A _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15966_ _15966_/A _15966_/B _15966_/C vssd1 vssd1 vccd1 vccd1 _15968_/A sky130_fd_sc_hd__or3_1
X_18754_ _18752_/X _18754_/B vssd1 vssd1 vccd1 vccd1 _18755_/B sky130_fd_sc_hd__and2b_1
X_11089_ _11089_/A _11089_/B vssd1 vssd1 vccd1 vccd1 _11112_/S sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18748__A2 _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14917_ _14918_/B _15206_/A vssd1 vssd1 vccd1 vccd1 _14922_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__13155__B _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17705_ _17705_/A _17705_/B vssd1 vssd1 vccd1 vccd1 _17705_/X sky130_fd_sc_hd__or2_1
X_15897_ _16029_/A _15898_/B vssd1 vssd1 vccd1 vccd1 _16034_/B sky130_fd_sc_hd__nor2_1
X_18685_ _18686_/A _18686_/B vssd1 vssd1 vccd1 vccd1 _18837_/A sky130_fd_sc_hd__or2_2
XFILLER_0_136_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14848_ _14848_/A _14848_/B _14848_/C vssd1 vssd1 vccd1 vccd1 _14848_/Y sky130_fd_sc_hd__nand3_1
X_17636_ _18010_/A _17636_/B vssd1 vssd1 vccd1 vccd1 _17640_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15431__A1 _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15431__B2 _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15370__B _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17567_ _17567_/A _17567_/B _17567_/C vssd1 vssd1 vccd1 vccd1 _17570_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_129_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14779_ _14625_/A _14624_/A _14624_/B _14620_/B _14620_/A vssd1 vssd1 vccd1 vccd1
+ _14780_/B sky130_fd_sc_hd__o32ai_4
XANTENNA__10795__A _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16518_ _16674_/A _16517_/B _16514_/X vssd1 vssd1 vccd1 vccd1 _16534_/A sky130_fd_sc_hd__a21o_1
XANTENNA__19173__A2 _19169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19306_ _19307_/A _19307_/B vssd1 vssd1 vccd1 vccd1 _19306_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_129_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17498_ _17498_/A _17498_/B vssd1 vssd1 vccd1 vccd1 _17500_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16449_ _16449_/A _16449_/B vssd1 vssd1 vccd1 vccd1 _16456_/B sky130_fd_sc_hd__xor2_2
X_19237_ _19692_/A _19238_/C _19692_/B _19068_/C vssd1 vssd1 vccd1 vccd1 _19240_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_874 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12548__A2 _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_121_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19168_ _17841_/Y _18394_/Y _19164_/X _19167_/X vssd1 vssd1 vccd1 vccd1 _19169_/B
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_147_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18119_ _18119_/A _18119_/B vssd1 vssd1 vccd1 vccd1 _18120_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__15098__A _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19793__A _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19099_ _19099_/A _19099_/B _19099_/C vssd1 vssd1 vccd1 vccd1 _19101_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_44_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15498__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21130_ _21238_/B _21130_/B _21131_/B vssd1 vssd1 vccd1 vccd1 _21244_/A sky130_fd_sc_hd__and3_1
XFILLER_0_83_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21061_ _21061_/A _21061_/B vssd1 vssd1 vccd1 vccd1 _21062_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__17239__A2 _17557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout404 _13155_/D vssd1 vssd1 vccd1 vccd1 _12326_/D sky130_fd_sc_hd__buf_4
XFILLER_0_111_297 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13049__C _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout415 _15217_/A vssd1 vssd1 vccd1 vccd1 _14859_/A sky130_fd_sc_hd__clkbuf_8
Xfanout426 _12781_/D vssd1 vssd1 vccd1 vccd1 _12223_/A sky130_fd_sc_hd__buf_4
X_20012_ _20154_/B _20012_/B _20012_/C vssd1 vssd1 vccd1 vccd1 _20125_/A sky130_fd_sc_hd__nand3_1
XANTENNA__20243__A1 _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout437 _21761_/Q vssd1 vssd1 vccd1 vccd1 _12780_/A sky130_fd_sc_hd__buf_4
Xfanout448 _12458_/A vssd1 vssd1 vccd1 vccd1 _12261_/A sky130_fd_sc_hd__buf_4
Xfanout459 _21755_/Q vssd1 vssd1 vccd1 vccd1 _15234_/C sky130_fd_sc_hd__buf_4
XANTENNA_fanout387_A _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20170__C _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18739__A2 _19060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11786__A1_N _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21963_ _21963_/CLK _21963_/D vssd1 vssd1 vccd1 vccd1 hold254/A sky130_fd_sc_hd__dfxtp_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout554_A _14774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20546__A2 _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20914_ _20914_/A _20914_/B vssd1 vssd1 vccd1 vccd1 _21033_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_7_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15422__A1 _15243_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21894_ _21938_/CLK _21894_/D vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20845_ _20721_/D _21293_/B _21853_/Q _20845_/D vssd1 vssd1 vccd1 vccd1 _20848_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_76_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout11 _11446_/S vssd1 vssd1 vccd1 vccd1 _11401_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_65_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout22 fanout23/X vssd1 vssd1 vccd1 vccd1 fanout22/X sky130_fd_sc_hd__buf_4
XFILLER_0_119_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13984__A1 _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout33 _21490_/S vssd1 vssd1 vccd1 vccd1 _21481_/S sky130_fd_sc_hd__clkbuf_8
Xfanout44 _11548_/Y vssd1 vssd1 vccd1 vccd1 _19636_/A sky130_fd_sc_hd__buf_2
X_20776_ _20776_/A _20776_/B vssd1 vssd1 vccd1 vccd1 _20911_/A sky130_fd_sc_hd__nor2_2
XANTENNA__20907__A _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout55 _11084_/S vssd1 vssd1 vccd1 vccd1 _11087_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_147_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout66 _20841_/B vssd1 vssd1 vccd1 vccd1 _21291_/B sky130_fd_sc_hd__buf_4
XFILLER_0_107_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout77 _21848_/Q vssd1 vssd1 vccd1 vccd1 _20193_/D sky130_fd_sc_hd__buf_4
Xfanout88 _21845_/Q vssd1 vssd1 vccd1 vccd1 _19053_/B sky130_fd_sc_hd__buf_4
XFILLER_0_52_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout99 _19060_/B vssd1 vssd1 vccd1 vccd1 _19382_/B sky130_fd_sc_hd__buf_4
XFILLER_0_52_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11211__A2 _11122_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15439__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12130_ _12130_/A _12130_/B vssd1 vssd1 vccd1 vccd1 _12130_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21328_ hold121/X _11553_/Y _21326_/X _21327_/X vssd1 vssd1 vccd1 vccd1 _21917_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21259_ _21259_/A _21259_/B vssd1 vssd1 vccd1 vccd1 _21260_/B sky130_fd_sc_hd__xnor2_2
X_12061_ _12058_/X _12061_/B vssd1 vssd1 vccd1 vccd1 _12104_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16438__B1 _12291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ mstream_o[86] hold18/X _11012_/S vssd1 vssd1 vccd1 vccd1 _21623_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18469__D _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15820_ _15817_/A _15818_/Y _15642_/Y _15644_/Y vssd1 vssd1 vccd1 vccd1 _15820_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13256__A _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15174__C _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15751_ _15752_/A _15752_/B vssd1 vssd1 vccd1 vccd1 _15751_/X sky130_fd_sc_hd__or2_1
XFILLER_0_99_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12963_ _13394_/A _14155_/C _12839_/X _12844_/A vssd1 vssd1 vccd1 vccd1 _12964_/B
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__17670__B _17670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14702_ _15375_/A _16268_/B _14702_/C _14702_/D vssd1 vssd1 vccd1 vccd1 _14702_/Y
+ sky130_fd_sc_hd__nand4_2
XTAP_3364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18470_ _18470_/A _18626_/B vssd1 vssd1 vccd1 vccd1 _18473_/A sky130_fd_sc_hd__or2_1
X_11914_ _11914_/A _11914_/B _11914_/C vssd1 vssd1 vccd1 vccd1 _11989_/A sky130_fd_sc_hd__nand3_1
X_15682_ _15682_/A _15682_/B _15682_/C vssd1 vssd1 vccd1 vccd1 _15683_/C sky130_fd_sc_hd__nand3_2
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_320 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12894_ _12891_/Y _12892_/X _12761_/X _12763_/X vssd1 vssd1 vccd1 vccd1 _12895_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_3386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_331 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14216__A2 _14873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17421_ _17520_/B _20249_/A _17309_/B _17307_/X vssd1 vssd1 vccd1 vccd1 _17423_/B
+ sky130_fd_sc_hd__a31o_1
X_14633_ _15435_/A _15788_/B _14498_/X _14499_/X _15653_/C vssd1 vssd1 vccd1 vccd1
+ _14638_/A sky130_fd_sc_hd__a32o_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _11845_/A _11845_/B _11845_/C vssd1 vssd1 vccd1 vccd1 _11917_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_68_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14087__A _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17352_ _17351_/B _17351_/C _17351_/A vssd1 vssd1 vccd1 vccd1 _17352_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_32_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14564_ _14713_/B _16380_/B _16173_/B _14713_/A vssd1 vssd1 vccd1 vccd1 _14568_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ _12297_/B _11776_/B _11776_/C _11776_/D vssd1 vssd1 vccd1 vccd1 _11776_/X
+ sky130_fd_sc_hd__or4_2
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16303_ _16303_/A _16303_/B vssd1 vssd1 vccd1 vccd1 _16343_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_144_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12319__B _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13515_ _16363_/A hold136/X _11066_/Y fanout6/X _13514_/Y vssd1 vssd1 vccd1 vccd1
+ _13515_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11223__B _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17283_ _17504_/C _17490_/A _17739_/C _17739_/D vssd1 vssd1 vccd1 vccd1 _17283_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_27_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14495_ _14496_/A _14496_/B vssd1 vssd1 vccd1 vccd1 _14611_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_27_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19022_ _19024_/A _19024_/B _19024_/C vssd1 vssd1 vccd1 vccd1 _19174_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16234_ _16075_/A _16077_/X _16302_/B _16233_/X vssd1 vssd1 vccd1 vccd1 _16235_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__16733__C _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13446_ _13447_/A _13447_/B vssd1 vssd1 vccd1 vccd1 _13446_/X sky130_fd_sc_hd__and2_1
XFILLER_0_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12980__D _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16165_ _16165_/A _16165_/B vssd1 vssd1 vccd1 vccd1 _16167_/B sky130_fd_sc_hd__or2_1
XFILLER_0_3_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14619__A1_N _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13377_ _13682_/C _13997_/C _13253_/X _13254_/X _13858_/C vssd1 vssd1 vccd1 vccd1
+ _13384_/A sky130_fd_sc_hd__a32oi_4
XFILLER_0_51_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15116_ _15116_/A _15116_/B vssd1 vssd1 vccd1 vccd1 _15126_/A sky130_fd_sc_hd__or2_1
XFILLER_0_2_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12328_ _12326_/X _12328_/B vssd1 vssd1 vccd1 vccd1 _12329_/B sky130_fd_sc_hd__and2b_1
X_16096_ _16096_/A _16207_/B vssd1 vssd1 vccd1 vccd1 _16098_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11596__D _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15646__A _16036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15047_ _15044_/Y _15045_/X _14883_/X _14887_/C vssd1 vssd1 vccd1 vccd1 _15047_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19924_ _19923_/A _19923_/B _19921_/Y _19922_/X vssd1 vssd1 vccd1 vccd1 _19925_/B
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__21367__B _21367_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12259_ _12259_/A _12259_/B vssd1 vssd1 vccd1 vccd1 _12259_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__19091__A1 _19092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19855_ _20091_/A _19855_/B _19950_/B vssd1 vssd1 vccd1 vccd1 _19857_/B sky130_fd_sc_hd__nand3_1
XANTENNA__19091__B2 _19092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17283__D _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk_i clk_i vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk_i/X sky130_fd_sc_hd__clkbuf_16
XANTENNA__17861__A _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18806_ _18805_/A _18805_/B _18805_/C vssd1 vssd1 vccd1 vccd1 _18807_/C sky130_fd_sc_hd__a21o_1
X_19786_ _19796_/A _19786_/B vssd1 vssd1 vccd1 vccd1 _20081_/A sky130_fd_sc_hd__and2_1
X_16998_ _16999_/A _16999_/B _16999_/C vssd1 vssd1 vccd1 vccd1 _17005_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__12501__C _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18737_ _19373_/B _19051_/A _19057_/C _19057_/D vssd1 vssd1 vccd1 vccd1 _18737_/X
+ sky130_fd_sc_hd__and4_1
X_15949_ _15948_/B _15948_/C _15948_/A vssd1 vssd1 vccd1 vccd1 _15949_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18668_ _18669_/A _18669_/B _18669_/C _18669_/D vssd1 vssd1 vccd1 vccd1 _18668_/Y
+ sky130_fd_sc_hd__nor4_2
XANTENNA__16601__B1 _17443_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13613__B _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17619_ _17619_/A _17619_/B _17739_/C _17739_/D vssd1 vssd1 vccd1 vccd1 _17737_/A
+ sky130_fd_sc_hd__and4_1
X_18599_ _18464_/D _18465_/B _18597_/Y _18598_/X vssd1 vssd1 vccd1 vccd1 _18757_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20630_ _20499_/A _20499_/Y _20628_/X _20629_/X vssd1 vssd1 vccd1 vccd1 _20630_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_129_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12229__B _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20561_ _20564_/D vssd1 vssd1 vccd1 vccd1 _20561_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_156_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17739__C _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20492_ _20492_/A vssd1 vssd1 vccd1 vccd1 _20492_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15839__A2_N _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout302_A _21795_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14465__A2_N _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21113_ _21109_/Y _21110_/X _20993_/Y _20997_/A vssd1 vssd1 vccd1 vccd1 _21113_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15556__A _15556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22093_ _22105_/CLK _22093_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[29] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout201 _21818_/Q vssd1 vssd1 vccd1 vccd1 _21256_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__12899__B _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22072__RESET_B fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout212 _21283_/A vssd1 vssd1 vccd1 vccd1 _19866_/C sky130_fd_sc_hd__buf_4
XANTENNA__21413__B1 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21044_ _21161_/A vssd1 vssd1 vccd1 vccd1 _21046_/D sky130_fd_sc_hd__inv_2
Xfanout223 hold328/X vssd1 vssd1 vccd1 vccd1 _21311_/A sky130_fd_sc_hd__clkbuf_4
Xfanout234 _17924_/B vssd1 vssd1 vccd1 vccd1 _19705_/B sky130_fd_sc_hd__buf_2
Xfanout245 _21261_/A vssd1 vssd1 vccd1 vccd1 _21199_/A sky130_fd_sc_hd__buf_4
Xfanout256 _18166_/A vssd1 vssd1 vccd1 vccd1 _19892_/A sky130_fd_sc_hd__clkbuf_8
Xfanout267 _21802_/Q vssd1 vssd1 vccd1 vccd1 _18030_/B sky130_fd_sc_hd__clkbuf_4
Xfanout278 _21799_/Q vssd1 vssd1 vccd1 vccd1 _16860_/C sky130_fd_sc_hd__clkbuf_8
Xfanout289 _17874_/A vssd1 vssd1 vccd1 vccd1 _17619_/A sky130_fd_sc_hd__buf_6
XANTENNA__21293__A _21293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17490__B _21792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16387__A _16387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20519__A2 _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21946_ _21949_/CLK _21946_/D vssd1 vssd1 vccd1 vccd1 hold77/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__17396__A1 _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout48_A fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17396__B2 _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21877_ _21942_/CLK _21877_/D vssd1 vssd1 vccd1 vccd1 hold79/A sky130_fd_sc_hd__dfxtp_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ _12109_/C _12528_/B _11630_/C _11683_/A vssd1 vssd1 vccd1 vccd1 _11683_/B
+ sky130_fd_sc_hd__nand4_2
X_20828_ _20699_/B _20700_/Y _20826_/Y _20827_/X vssd1 vssd1 vccd1 vccd1 _20830_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18896__A1 _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11561_ _12223_/A _12637_/B _11560_/B _11557_/X vssd1 vssd1 vccd1 vccd1 _11573_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__18896__B2 _19230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20759_ _20623_/X _20627_/C _20757_/X _20758_/Y vssd1 vssd1 vccd1 vccd1 _20759_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_147_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13709__A1 _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13300_ _13300_/A _13300_/B vssd1 vssd1 vccd1 vccd1 _13302_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13709__B2 _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14280_ _14117_/B _14280_/B vssd1 vssd1 vccd1 vccd1 _14282_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_150_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11492_ _11507_/A1 t1y[14] t0x[14] _11501_/B2 vssd1 vssd1 vccd1 vccd1 _11492_/X sky130_fd_sc_hd__a22o_1
XANTENNA__14354__B _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ _13127_/A _13126_/B _13126_/A vssd1 vssd1 vccd1 vccd1 _13242_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__18648__A1 _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12155__A _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12393__B1 _11045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13162_ _13162_/A _13287_/A _13162_/C vssd1 vssd1 vccd1 vccd1 _13287_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_20_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12113_ _12102_/A _12102_/B _12102_/C vssd1 vssd1 vccd1 vccd1 _12115_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__14134__B2 _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ fanout9/X _21352_/B vssd1 vssd1 vccd1 vccd1 _13093_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17871__A2 _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17970_ _17968_/Y _17970_/B vssd1 vssd1 vccd1 vccd1 _17970_/X sky130_fd_sc_hd__and2b_2
XFILLER_0_20_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17384__C _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16921_ _16920_/B _16920_/C _16920_/A vssd1 vssd1 vccd1 vccd1 _16923_/B sky130_fd_sc_hd__a21bo_1
X_12044_ _12094_/A _12094_/B _12530_/A _12512_/A vssd1 vssd1 vccd1 vccd1 _12044_/X
+ sky130_fd_sc_hd__and4_1
X_19640_ _19640_/A _19640_/B vssd1 vssd1 vccd1 vccd1 _19777_/A sky130_fd_sc_hd__or2_1
X_16852_ _16785_/A _16785_/B _16785_/C vssd1 vssd1 vccd1 vccd1 _16852_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__15634__A1 _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16831__B1 _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15803_ _15803_/A _15803_/B vssd1 vssd1 vccd1 vccd1 _15811_/A sky130_fd_sc_hd__nor2_1
XANTENNA__21407__S _21407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16783_ _16783_/A _16783_/B _16783_/C vssd1 vssd1 vccd1 vccd1 _16784_/B sky130_fd_sc_hd__and3_1
X_19571_ _19972_/A _20394_/B _19866_/D _19874_/B vssd1 vssd1 vccd1 vccd1 _19575_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_137_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13995_ _13859_/A _13861_/B _13859_/B vssd1 vssd1 vccd1 vccd1 _14000_/A sky130_fd_sc_hd__o21bai_2
X_15734_ _15733_/B _15733_/C _15733_/A vssd1 vssd1 vccd1 vccd1 _15734_/Y sky130_fd_sc_hd__o21ai_2
X_18522_ _18521_/A _18521_/B _18521_/C _18521_/D vssd1 vssd1 vccd1 vccd1 _18522_/Y
+ sky130_fd_sc_hd__o22ai_1
XTAP_3150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21724__RESET_B _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12946_ _12961_/B _12945_/B _12945_/C vssd1 vssd1 vccd1 vccd1 _12950_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_137_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15665_ _15665_/A _15665_/B vssd1 vssd1 vccd1 vccd1 _15667_/B sky130_fd_sc_hd__xor2_1
XTAP_3194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18453_ _18453_/A _18453_/B _18453_/C vssd1 vssd1 vccd1 vccd1 _18454_/B sky130_fd_sc_hd__and3_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12877_ _12877_/A _12877_/B _13152_/D vssd1 vssd1 vccd1 vccd1 _12877_/X sky130_fd_sc_hd__and3_1
XANTENNA_150 v1z[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_161 v2z[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14248__C _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14616_ _15829_/C _14615_/X _14614_/X vssd1 vssd1 vccd1 vccd1 _14618_/A sky130_fd_sc_hd__a21bo_2
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17404_ _17404_/A _17404_/B _17404_/C vssd1 vssd1 vccd1 vccd1 _17405_/C sky130_fd_sc_hd__and3_1
XANTENNA_172 v2z[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_183 _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18384_ _18380_/Y _18381_/X _18125_/Y _18128_/Y vssd1 vssd1 vccd1 vccd1 _18385_/B
+ sky130_fd_sc_hd__o211ai_2
X_11828_ _11833_/A _11610_/Y _11609_/X _11601_/X vssd1 vssd1 vccd1 vccd1 _11830_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15596_ _15596_/A _15596_/B vssd1 vssd1 vccd1 vccd1 _15598_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_194 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13152__C _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17139__A1 _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20547__A _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16744__B _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17335_ _17335_/A _17335_/B vssd1 vssd1 vccd1 vccd1 _17336_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_44_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14547_ _14690_/A _14546_/C _14546_/A vssd1 vssd1 vccd1 vccd1 _14548_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_83_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11759_ _11758_/B _11758_/C _11758_/A vssd1 vssd1 vccd1 vccd1 _11761_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__12620__A1 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12620__B2 _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12991__C _13269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16463__C _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17266_ _17267_/A _17267_/B vssd1 vssd1 vccd1 vccd1 _17479_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14478_ _15159_/D _15174_/D _14479_/C _14632_/A vssd1 vssd1 vccd1 vccd1 _14480_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_141_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16217_ _16409_/A _21784_/Q _16218_/C _16218_/D vssd1 vssd1 vccd1 vccd1 _16219_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_113_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19005_ _18889_/A _18889_/C _18889_/B vssd1 vssd1 vccd1 vccd1 _19152_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_148_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13429_ _13428_/A _13428_/B _13415_/Y vssd1 vssd1 vccd1 vccd1 _13429_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__18639__A1 _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15570__B1 _15426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17197_ _17197_/A _17197_/B vssd1 vssd1 vccd1 vccd1 _17198_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16760__A _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16148_ _16036_/A _16036_/B _15907_/A vssd1 vssd1 vccd1 vccd1 _16152_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_23_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17311__A1 _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19493__D _19493_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16079_ _16079_/A _16079_/B _16079_/C vssd1 vssd1 vccd1 vccd1 _16079_/X sky130_fd_sc_hd__or3_2
XANTENNA__17862__A2 _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19907_ _20148_/C _20273_/A _19908_/C _20001_/A vssd1 vssd1 vccd1 vccd1 _19909_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12512__B _12621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19838_ _19840_/A _19840_/B vssd1 vssd1 vccd1 vccd1 _19838_/X sky130_fd_sc_hd__or2_1
XFILLER_0_39_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19769_ _19769_/A _19769_/B vssd1 vssd1 vccd1 vccd1 _19772_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_155_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13624__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21800_ _21803_/CLK _21800_/D vssd1 vssd1 vccd1 vccd1 _21800_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21731_ _22020_/CLK _21731_/D vssd1 vssd1 vccd1 vccd1 _21731_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20921__A2 _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21662_ _21934_/CLK _21662_/D vssd1 vssd1 vccd1 vccd1 hold81/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20613_ _20613_/A _20613_/B vssd1 vssd1 vccd1 vccd1 _20616_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__12611__A1 _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13997__C _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21593_ _21888_/CLK _21593_/D _11041_/A vssd1 vssd1 vccd1 vccd1 mstream_o[56] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout517_A _21740_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20544_ _21291_/A _21264_/A _20544_/C _20730_/A vssd1 vssd1 vccd1 vccd1 _20730_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_116_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14364__A1 _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14364__B2 _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20475_ _20478_/D vssd1 vssd1 vccd1 vccd1 _20475_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17302__A1 _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17302__B2 _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_381 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14621__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22076_ _22080_/CLK _22076_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[12] sky130_fd_sc_hd__dfrtp_4
XANTENNA__19055__B2 _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21027_ _21027_/A _21027_/B vssd1 vssd1 vccd1 vccd1 _21027_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12800_ _12687_/B _12687_/Y _12797_/X _12799_/Y vssd1 vssd1 vccd1 vccd1 _12803_/C
+ sky130_fd_sc_hd__a211oi_4
X_13780_ _13779_/B _13779_/C _13779_/A vssd1 vssd1 vccd1 vccd1 _13782_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_69_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10992_ mstream_o[66] hold143/X _10992_/S vssd1 vssd1 vccd1 vccd1 _21603_/D sky130_fd_sc_hd__mux2_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12731_ _12731_/A _12731_/B vssd1 vssd1 vccd1 vccd1 _12744_/A sky130_fd_sc_hd__xor2_2
X_21929_ _21932_/CLK _21929_/D vssd1 vssd1 vccd1 vccd1 hold94/A sky130_fd_sc_hd__dfxtp_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15450_ _15450_/A _15450_/B vssd1 vssd1 vccd1 vccd1 _15461_/A sky130_fd_sc_hd__or2_1
XANTENNA__19221__A _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12662_ _12897_/C _12660_/X _12661_/X vssd1 vssd1 vccd1 vccd1 _12663_/B sky130_fd_sc_hd__a21bo_1
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18318__B1 _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14401_ _14397_/X _14399_/Y _14224_/B _14226_/B vssd1 vssd1 vccd1 vccd1 _14402_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _12858_/C _12312_/A vssd1 vssd1 vccd1 vccd1 _11897_/B sky130_fd_sc_hd__nand2_1
X_15381_ _15382_/A _15382_/B vssd1 vssd1 vccd1 vccd1 _15381_/Y sky130_fd_sc_hd__nand2_2
XANTENNA__12602__A1 _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12593_ _12589_/X _12590_/Y _12415_/X _12418_/Y vssd1 vssd1 vccd1 vccd1 _12593_/Y
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12602__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14365__A _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17120_ _17120_/A _17120_/B vssd1 vssd1 vccd1 vccd1 _17120_/X sky130_fd_sc_hd__or2_1
XFILLER_0_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14332_ _14331_/B _14331_/C _14331_/A vssd1 vssd1 vccd1 vccd1 _14333_/C sky130_fd_sc_hd__a21o_1
XANTENNA__20676__A1 _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11544_ _11544_/A1 t2x[31] v1z[31] fanout21/X _11543_/X vssd1 vssd1 vccd1 vccd1 _11544_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14084__B _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14355__A1 _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13158__A2 _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17051_ _17049_/B _17049_/C _17049_/A vssd1 vssd1 vccd1 vccd1 _17117_/B sky130_fd_sc_hd__a21o_1
X_14263_ _14260_/X _14261_/Y _14101_/B _14101_/Y vssd1 vssd1 vccd1 vccd1 _14264_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_64_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11475_ _11502_/A1 t2x[8] v1z[8] fanout20/X _11474_/X vssd1 vssd1 vccd1 vccd1 _11475_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16002_ _15999_/Y _16000_/X _15826_/Y _15874_/X vssd1 vssd1 vccd1 vccd1 _16002_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__20814__B _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13214_ _13213_/B _13213_/C _13213_/A vssd1 vssd1 vccd1 vccd1 _13214_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_61_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14194_ _14195_/A _16286_/A _14195_/C _14362_/A vssd1 vssd1 vccd1 vccd1 _14196_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17395__B _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13145_ _13142_/X _13143_/Y _13029_/B _13031_/A vssd1 vssd1 vccd1 vccd1 _13145_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_131_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17844__A2 _19030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13076_ _13072_/X _13073_/Y _12931_/X _12934_/X vssd1 vssd1 vccd1 vccd1 _13077_/C
+ sky130_fd_sc_hd__a211o_1
X_17953_ _17953_/A _17953_/B _17953_/C vssd1 vssd1 vccd1 vccd1 _17953_/X sky130_fd_sc_hd__or3_2
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17057__B1 _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16904_ _16844_/A _16844_/B _16849_/C _16844_/D vssd1 vssd1 vccd1 vccd1 _16904_/X
+ sky130_fd_sc_hd__o22a_1
X_12027_ _12027_/A _12027_/B vssd1 vssd1 vccd1 vccd1 _12029_/C sky130_fd_sc_hd__xnor2_1
X_17884_ _17884_/A vssd1 vssd1 vccd1 vccd1 _17884_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_40_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11341__B2 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19623_ _19624_/B _19624_/A vssd1 vssd1 vccd1 vccd1 _19779_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__15643__B _15643_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16835_ _17300_/C _17387_/A vssd1 vssd1 vccd1 vccd1 _16894_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_16_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21788_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__19349__A2 _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19554_ _19554_/A _19554_/B _19554_/C vssd1 vssd1 vccd1 vccd1 _19556_/B sky130_fd_sc_hd__nand3_1
X_13978_ _13980_/A _14142_/B vssd1 vssd1 vccd1 vccd1 _13981_/A sky130_fd_sc_hd__nor2_1
XANTENNA__13094__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16766_ _17300_/C _17277_/A _17387_/A _17520_/D vssd1 vssd1 vccd1 vccd1 _16767_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19008__A_N _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13094__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18505_ _18505_/A _18505_/B _18505_/C vssd1 vssd1 vccd1 vccd1 _18508_/A sky130_fd_sc_hd__nand3_2
X_15717_ _16084_/A _15717_/B _15717_/C _15976_/D vssd1 vssd1 vccd1 vccd1 _15848_/A
+ sky130_fd_sc_hd__and4_1
X_12929_ _12929_/A _12929_/B _12929_/C vssd1 vssd1 vccd1 vccd1 _12929_/X sky130_fd_sc_hd__or3_2
XFILLER_0_76_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16697_ _16697_/A _16697_/B vssd1 vssd1 vccd1 vccd1 _16698_/C sky130_fd_sc_hd__nor2_1
X_19485_ _19405_/A _19405_/B _19404_/A vssd1 vssd1 vccd1 vccd1 _19524_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_88_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18436_ _18287_/A _18287_/B _18286_/B vssd1 vssd1 vccd1 vccd1 _18438_/B sky130_fd_sc_hd__o21ai_1
X_15648_ _15907_/A _15648_/B _15648_/C vssd1 vssd1 vccd1 vccd1 _15650_/A sky130_fd_sc_hd__nor3_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15579_ _15439_/D _21788_/Q _16314_/D _15579_/D vssd1 vssd1 vccd1 vccd1 _15712_/A
+ sky130_fd_sc_hd__and4b_2
X_18367_ _18368_/A _18368_/B _18368_/C _18368_/D vssd1 vssd1 vccd1 vccd1 _18367_/Y
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_90_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17318_ _17212_/X _17214_/X _17316_/X _17317_/Y vssd1 vssd1 vccd1 vccd1 _17356_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_83_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18298_ _18167_/D _18169_/A _18296_/X _18442_/B vssd1 vssd1 vccd1 vccd1 _18453_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_71_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17249_ _17248_/A _17248_/B _17248_/C vssd1 vssd1 vccd1 vccd1 _17251_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20260_ _20260_/A _20260_/B _20260_/C vssd1 vssd1 vccd1 vccd1 _20260_/X sky130_fd_sc_hd__and3_1
XFILLER_0_113_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13619__A _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17835__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20191_ _20975_/D _20845_/D _20733_/C _20606_/D vssd1 vssd1 vccd1 vccd1 _20329_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_45_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13857__B1 _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12242__B _12242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13321__A2 _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11332__A1 _11331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21395__A2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13872__A3 _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_600 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout467_A _14698_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11096__A0 _11057_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout634_A _16380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21714_ _22105_/CLK _21714_/D vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14034__B1 _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1068 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21721__D _21721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21645_ _21722_/CLK _21645_/D fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[108]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__14185__A _14659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_50 hold275/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17523__A1 _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12060__A2 _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19695__B _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21576_ mstream_o[39] _11059_/Y _21579_/S vssd1 vssd1 vccd1 vccd1 _22103_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_74_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_61 hold270/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_72 hold268/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_83 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20527_ _20249_/A _20526_/X _20657_/A vssd1 vssd1 vccd1 vccd1 _20529_/B sky130_fd_sc_hd__a21oi_1
XANTENNA_94 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12136__C _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ _12109_/C _11259_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21766_/D sky130_fd_sc_hd__mux2_1
X_20458_ _20590_/D _21291_/B _20458_/C _20458_/D vssd1 vssd1 vccd1 vccd1 _20588_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_123_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11191_ hold131/X fanout22/X _11190_/X vssd1 vssd1 vccd1 vccd1 _11191_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20389_ _20910_/A _21278_/B _20390_/C _20559_/A vssd1 vssd1 vccd1 vccd1 _20391_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20650__A _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14950_ _15579_/D _15174_/D _14951_/C _15169_/A vssd1 vssd1 vccd1 vccd1 _14952_/B
+ sky130_fd_sc_hd__a22o_1
X_22059_ _22063_/CLK _22059_/D vssd1 vssd1 vccd1 vccd1 hold262/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__11323__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21386__A2 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13901_ _13901_/A _13901_/B _13901_/C vssd1 vssd1 vccd1 vccd1 _13901_/X sky130_fd_sc_hd__and3_1
X_14881_ _14881_/A _14881_/B _14881_/C vssd1 vssd1 vccd1 vccd1 _14883_/B sky130_fd_sc_hd__nand3_2
XANTENNA__16262__A1 _15907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13832_ _13833_/A _13833_/B vssd1 vssd1 vccd1 vccd1 _13834_/A sky130_fd_sc_hd__and2_1
X_16620_ _17145_/A _17434_/B vssd1 vssd1 vccd1 vccd1 _16622_/B sky130_fd_sc_hd__and2_1
XANTENNA__18539__B1 _18537_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11087__A0 _10984_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16551_ _16552_/A _16552_/B vssd1 vssd1 vccd1 vccd1 _16551_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13763_ _14557_/B _14873_/B _13913_/C _14557_/A vssd1 vssd1 vccd1 vccd1 _13766_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10975_ hold128/A hold146/A vssd1 vssd1 vccd1 vccd1 _10977_/A sky130_fd_sc_hd__or2_1
XANTENNA__16575__A _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15502_ _15502_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _16261_/B sky130_fd_sc_hd__and2_1
XANTENNA__18493__C _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12714_ _13394_/A _14176_/C _12617_/A _12614_/X vssd1 vssd1 vccd1 vccd1 _12716_/C
+ sky130_fd_sc_hd__a31oi_2
X_16482_ _16479_/X _16482_/B vssd1 vssd1 vccd1 vccd1 _16758_/B sky130_fd_sc_hd__and2b_1
X_19270_ _19271_/A _19406_/B _19271_/C vssd1 vssd1 vccd1 vccd1 _19270_/X sky130_fd_sc_hd__and3_1
X_13694_ _13538_/Y _13541_/X _13691_/Y _13693_/X vssd1 vssd1 vccd1 vccd1 _13698_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_85_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15433_ _15577_/A vssd1 vssd1 vccd1 vccd1 _15435_/D sky130_fd_sc_hd__inv_2
X_18221_ _18220_/A _18220_/B _18220_/C _18220_/D vssd1 vssd1 vccd1 vccd1 _18221_/Y
+ sky130_fd_sc_hd__o22ai_2
X_12645_ _12643_/X _12645_/B vssd1 vssd1 vccd1 vccd1 _12646_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_127_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15364_ _15365_/B vssd1 vssd1 vccd1 vccd1 _15364_/Y sky130_fd_sc_hd__inv_2
X_18152_ _18152_/A _18304_/A _18152_/C vssd1 vssd1 vccd1 vccd1 _18304_/B sky130_fd_sc_hd__nand3_4
XANTENNA__20247__D _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12576_ _12575_/A _12575_/B _12575_/C vssd1 vssd1 vccd1 vccd1 _12578_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_92_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21420__S _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14315_ _14315_/A _14315_/B vssd1 vssd1 vccd1 vccd1 _14316_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_4_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17103_ _17029_/A _17146_/D _17094_/B _17096_/X vssd1 vssd1 vccd1 vccd1 _17104_/B
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__15919__A _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18083_ _18082_/B _18082_/C _18082_/A vssd1 vssd1 vccd1 vccd1 _18083_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_13_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11527_ _11526_/X _19199_/D _11545_/S vssd1 vssd1 vccd1 vccd1 _21847_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15295_ _15295_/A _15295_/B vssd1 vssd1 vccd1 vccd1 _15342_/A sky130_fd_sc_hd__or2_2
XFILLER_0_151_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20544__B _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17034_ _17035_/A _17035_/B vssd1 vssd1 vccd1 vccd1 _17034_/Y sky130_fd_sc_hd__nand2_1
X_14246_ _14090_/A _14090_/B _14090_/C vssd1 vssd1 vccd1 vccd1 _14254_/A sky130_fd_sc_hd__o21bai_1
Xhold309 hold309/A vssd1 vssd1 vccd1 vccd1 hold309/X sky130_fd_sc_hd__buf_4
XFILLER_0_151_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11458_ _11457_/X _19445_/A _11470_/S vssd1 vssd1 vccd1 vccd1 _21824_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_21_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14177_ _15112_/D _14176_/X _14175_/X vssd1 vssd1 vccd1 vccd1 _14179_/A sky130_fd_sc_hd__a21bo_1
X_11389_ _11388_/X _17526_/B _11401_/S vssd1 vssd1 vccd1 vccd1 _21801_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12343__A _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15828__B2 _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13128_ _13128_/A _13128_/B vssd1 vssd1 vccd1 vccd1 _13136_/A sky130_fd_sc_hd__nand2_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18949__B _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_43_clk_i_A _21822_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18985_ _18822_/C _18821_/Y _18983_/X _18984_/X vssd1 vssd1 vccd1 vccd1 _18985_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14500__A1 _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ _13059_/A _13059_/B _13059_/C vssd1 vssd1 vccd1 vccd1 _13062_/B sky130_fd_sc_hd__nand3_4
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17936_ _17935_/A _17935_/B _17935_/C vssd1 vssd1 vccd1 vccd1 _17937_/C sky130_fd_sc_hd__a21o_1
XANTENNA__18030__A _19823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11314__A1 _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15373__B _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17867_ _17867_/A _17867_/B vssd1 vssd1 vccd1 vccd1 _17869_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__10798__A _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19606_ _19606_/A _19606_/B _19606_/C vssd1 vssd1 vccd1 vccd1 _19608_/A sky130_fd_sc_hd__nand3_1
X_16818_ _16818_/A _16818_/B vssd1 vssd1 vccd1 vccd1 _16820_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17798_ _17797_/A _17797_/B _17797_/C vssd1 vssd1 vccd1 vccd1 _17799_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11078__A0 _10926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19537_ _19686_/A _20419_/A _19538_/C _19538_/D vssd1 vssd1 vccd1 vccd1 _19537_/X
+ sky130_fd_sc_hd__and4_1
X_16749_ _16749_/A _16749_/B vssd1 vssd1 vccd1 vccd1 _16751_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__17202__B1 _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19468_ _19468_/A _19468_/B vssd1 vssd1 vccd1 vccd1 _19469_/B sky130_fd_sc_hd__and2_1
XFILLER_0_9_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16556__A2 _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18419_ _18415_/Y _18417_/X _18264_/X _18266_/Y vssd1 vssd1 vccd1 vccd1 _18420_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19399_ _19398_/A _19398_/B _19398_/C vssd1 vssd1 vccd1 vccd1 _19400_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_51_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21430_ hold260/X sstream_i[7] _21489_/S vssd1 vssd1 vccd1 vccd1 _21957_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15829__A _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21361_ _21412_/A _21361_/B vssd1 vssd1 vccd1 vccd1 _21361_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout215_A _19868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20312_ _20462_/D _21291_/B _20312_/C _20312_/D vssd1 vssd1 vccd1 vccd1 _20460_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_13_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21292_ _21259_/A _21179_/A _21179_/B _21181_/Y vssd1 vssd1 vccd1 vccd1 _21294_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_3_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20243_ _20910_/A _21046_/B _20244_/C _20428_/A vssd1 vssd1 vccd1 vccd1 _20245_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11553__A1 _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18859__B _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20174_ _20176_/A _20314_/B vssd1 vssd1 vccd1 vccd1 _20177_/A sky130_fd_sc_hd__or2_1
XFILLER_0_110_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17763__B _19823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12403__D _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21368__A2 _18689_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11305__B2 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__B1 _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15283__B _15284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18297__D _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11069__A0 _10860_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17992__A1 _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17992__B2 _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14558__A1 _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12430_ _12430_/A _12430_/B vssd1 vssd1 vccd1 vccd1 _12433_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21628_ _21682_/CLK _21628_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[91] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12361_ _11727_/A _11727_/C _11727_/B vssd1 vssd1 vccd1 vccd1 _12362_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_117_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21559_ mstream_o[22] hold168/X _21562_/S vssd1 vssd1 vccd1 vccd1 _22086_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17657__C _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14100_ _14101_/A _14101_/B _14101_/C vssd1 vssd1 vccd1 vccd1 _14100_/X sky130_fd_sc_hd__and3_1
XFILLER_0_106_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11312_ _14176_/C _11311_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21779_/D sky130_fd_sc_hd__mux2_1
X_15080_ _15218_/A _15080_/B _15215_/B vssd1 vssd1 vccd1 vccd1 _15082_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_133_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12292_ _21725_/D hold156/X _11043_/X fanout6/X _12290_/Y vssd1 vssd1 vccd1 vccd1
+ _12292_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_105_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14031_ _14031_/A _14031_/B vssd1 vssd1 vccd1 vccd1 _14045_/A sky130_fd_sc_hd__xnor2_2
X_11243_ fanout59/X v0z[4] fanout19/X _11242_/X vssd1 vssd1 vccd1 vccd1 _11243_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11544__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18769__B _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11174_ _13155_/B _11173_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21741_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_98_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16483__A1 _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18770_ _18770_/A _18770_/B vssd1 vssd1 vccd1 vccd1 _18778_/A sky130_fd_sc_hd__xor2_1
X_15982_ _15983_/A _15983_/B vssd1 vssd1 vccd1 vccd1 _15982_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_100_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21359__A2 _13369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17721_ _17854_/B _19051_/C _18894_/B _18857_/B vssd1 vssd1 vccd1 vccd1 _17723_/B
+ sky130_fd_sc_hd__a22o_1
X_14933_ _14934_/A _14934_/B _14934_/C vssd1 vssd1 vccd1 vccd1 _14933_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12610__B _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17652_ _17652_/A _17652_/B _17652_/C vssd1 vssd1 vccd1 vccd1 _17652_/Y sky130_fd_sc_hd__nand3_4
X_14864_ _14865_/A _14865_/B _14865_/C _14865_/D vssd1 vssd1 vccd1 vccd1 _14868_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16603_ _16603_/A _16603_/B vssd1 vssd1 vccd1 vccd1 _16604_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_138_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13815_ fanout9/A _18689_/B vssd1 vssd1 vccd1 vccd1 _13815_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__20319__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14795_ _14784_/Y _14795_/B _14795_/C vssd1 vssd1 vccd1 vccd1 _14795_/X sky130_fd_sc_hd__and3b_1
X_17583_ _17579_/X _17581_/Y _17468_/Y _17470_/X vssd1 vssd1 vccd1 vccd1 _17584_/C
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__13722__A _13875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19322_ _19322_/A _19788_/B vssd1 vssd1 vccd1 vccd1 _19322_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13746_ _13746_/A _13746_/B vssd1 vssd1 vccd1 vccd1 _13756_/A sky130_fd_sc_hd__xnor2_1
X_16534_ _16534_/A _16534_/B _16534_/C vssd1 vssd1 vccd1 vccd1 _16537_/A sky130_fd_sc_hd__nand3_1
X_10958_ _10959_/B vssd1 vssd1 vccd1 vccd1 _10958_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_58_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14537__B _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19253_ _19252_/B _19252_/C _19252_/A vssd1 vssd1 vccd1 vccd1 _19254_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13677_ _13833_/A _13677_/B vssd1 vssd1 vccd1 vccd1 _13698_/A sky130_fd_sc_hd__or2_1
X_16465_ _17041_/A _17013_/D _17019_/C _16899_/B vssd1 vssd1 vccd1 vccd1 _16466_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10889_ hold216/A hold217/A vssd1 vssd1 vccd1 vccd1 _10899_/A sky130_fd_sc_hd__and2_1
XFILLER_0_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18204_ _18204_/A _18204_/B _18204_/C vssd1 vssd1 vccd1 vccd1 _18207_/A sky130_fd_sc_hd__nand3_1
X_15416_ _15417_/A _15417_/B vssd1 vssd1 vccd1 vccd1 _15560_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12628_ _12629_/A _12629_/B _12629_/C vssd1 vssd1 vccd1 vccd1 _12630_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_72_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16396_ _16396_/A _16396_/B vssd1 vssd1 vccd1 vccd1 _16398_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19184_ _19184_/A _19184_/B vssd1 vssd1 vccd1 vccd1 _19189_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__19488__A1 _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15347_ _15347_/A _15347_/B vssd1 vssd1 vccd1 vccd1 _15350_/A sky130_fd_sc_hd__xnor2_4
X_18135_ _19487_/A _19487_/B _19227_/C _19227_/D vssd1 vssd1 vccd1 vccd1 _18288_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13772__A2 _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ _13155_/B _12781_/D vssd1 vssd1 vccd1 vccd1 _12563_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15368__B _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15278_ _15279_/A _15279_/B vssd1 vssd1 vccd1 vccd1 _15419_/A sky130_fd_sc_hd__or2_1
XFILLER_0_112_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18066_ _18066_/A _18066_/B _18066_/C vssd1 vssd1 vccd1 vccd1 _18069_/A sky130_fd_sc_hd__nand3_1
Xhold106 hold106/A vssd1 vssd1 vccd1 vccd1 hold106/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 hold117/A vssd1 vssd1 vccd1 vccd1 hold117/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold128 hold128/A vssd1 vssd1 vccd1 vccd1 hold128/X sky130_fd_sc_hd__dlygate4sd3_1
X_14229_ _14228_/B _14228_/C _14228_/A vssd1 vssd1 vccd1 vccd1 _14230_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13524__A2 _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17017_ _17016_/B _17016_/C _17016_/A vssd1 vssd1 vccd1 vccd1 _17018_/C sky130_fd_sc_hd__a21bo_1
Xhold139 hold139/A vssd1 vssd1 vccd1 vccd1 hold139/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1170 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11535__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout608 _21718_/Q vssd1 vssd1 vccd1 vccd1 _11498_/A1 sky130_fd_sc_hd__buf_4
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18463__A2 _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout619 _21717_/Q vssd1 vssd1 vccd1 vccd1 _11027_/S sky130_fd_sc_hd__clkbuf_8
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20721__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13288__A1 _13875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18968_ _18967_/A _18967_/B _18967_/C vssd1 vssd1 vccd1 vccd1 _18969_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13288__B2 _13877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16199__B _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11299__B1 _11298_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17919_ _17919_/A _18047_/B _17919_/C vssd1 vssd1 vccd1 vccd1 _17921_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18899_ _19373_/B _19057_/D _18901_/C _18901_/D vssd1 vssd1 vccd1 vccd1 _18899_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19290__S _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20930_ _21842_/Q _21815_/Q _20930_/C _20930_/D vssd1 vssd1 vccd1 vccd1 _21048_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_135_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17974__A1 _17967_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16927__B _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20861_ _20991_/C _21296_/A _21283_/B _21305_/B vssd1 vssd1 vccd1 vccd1 _20985_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_135_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout165_A _16813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13460__A1 _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20792_ _21151_/A _20924_/A _21301_/A _21305_/A vssd1 vssd1 vccd1 vccd1 _20986_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12263__A2 _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout332_A _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12248__A _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17758__B _18008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21413_ _21720_/D _21027_/Y _21421_/S _21412_/Y vssd1 vssd1 vccd1 vccd1 _21413_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13763__A2 _14873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21344_ _21349_/A _17595_/Y _21421_/S _21343_/Y vssd1 vssd1 vccd1 vccd1 _21344_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14182__B _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21275_ _21275_/A _21275_/B vssd1 vssd1 vccd1 vccd1 _21277_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19692__C _19692_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11526__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21296__A _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20226_ _20224_/X _20226_/B vssd1 vssd1 vccd1 vccd1 _20372_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__17493__B _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20157_ _20157_/A _20157_/B vssd1 vssd1 vccd1 vccd1 _20159_/B sky130_fd_sc_hd__xor2_2
XANTENNA__14476__B1 _14635_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12711__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout78_A _21847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20088_ _20088_/A _20247_/D vssd1 vssd1 vccd1 vccd1 _20089_/B sky130_fd_sc_hd__nand2_1
XTAP_3502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16217__A1 _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_525 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21210__A1 _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21210__B2 _21311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ _12897_/C _12897_/D _13556_/A _12621_/C vssd1 vssd1 vccd1 vccd1 _11930_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__19954__A2 _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _12897_/C _12619_/A _13556_/A _12897_/D vssd1 vssd1 vccd1 vccd1 _11862_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_3579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13600_ _13600_/A _13600_/B vssd1 vssd1 vccd1 vccd1 _13602_/B sky130_fd_sc_hd__xor2_1
XTAP_2867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10812_ hold107/A hold104/A vssd1 vssd1 vccd1 vccd1 _10841_/B sky130_fd_sc_hd__or2_1
XANTENNA__17014__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14580_ _14580_/A _14580_/B vssd1 vssd1 vccd1 vccd1 _14583_/A sky130_fd_sc_hd__xor2_4
XTAP_2878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11792_ _11791_/A _11791_/C _11791_/B vssd1 vssd1 vccd1 vccd1 _11795_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14357__B _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13531_ _13528_/Y _13678_/A _13822_/B _16328_/B vssd1 vssd1 vccd1 vccd1 _13678_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_149_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16250_ _16250_/A _16250_/B vssd1 vssd1 vccd1 vccd1 _16253_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_125_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13462_ _13462_/A _13608_/B vssd1 vssd1 vccd1 vccd1 _13464_/B sky130_fd_sc_hd__or2_1
XFILLER_0_82_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12006__A2 _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15201_ _15201_/A _15201_/B vssd1 vssd1 vccd1 vccd1 _15203_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__16940__A2 _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12413_ _12413_/A _12413_/B vssd1 vssd1 vccd1 vccd1 _12414_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16181_ _16181_/A _16181_/B vssd1 vssd1 vccd1 vccd1 _16183_/A sky130_fd_sc_hd__xnor2_1
X_13393_ _13393_/A _13393_/B vssd1 vssd1 vccd1 vccd1 _13396_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15132_ _15129_/Y _15271_/A _15933_/C _16328_/A vssd1 vssd1 vccd1 vccd1 _15271_/B
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__12962__B1 _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12344_ _12444_/B _12897_/C _12897_/D _12877_/A vssd1 vssd1 vccd1 vccd1 _12345_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16153__B1 _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15063_ _15063_/A _15063_/B vssd1 vssd1 vccd1 vccd1 _15065_/B sky130_fd_sc_hd__xor2_1
XANTENNA__21029__B2 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19940_ _19942_/A _19942_/B _19942_/C vssd1 vssd1 vccd1 vccd1 _19941_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12275_ _12275_/A _12275_/B _12275_/C _12275_/D vssd1 vssd1 vccd1 vccd1 _12275_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_120_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11517__A1 _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14014_ _14131_/B _14012_/X _13886_/Y _13889_/Y vssd1 vssd1 vccd1 vccd1 _14015_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__11517__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11226_ _21718_/D t1x[0] v2z[0] _21724_/D _11225_/X vssd1 vssd1 vccd1 vccd1 _11226_/X
+ sky130_fd_sc_hd__a221o_2
X_19871_ _19972_/A _20394_/B _19872_/C _19972_/C vssd1 vssd1 vccd1 vccd1 _19871_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__15916__B _15916_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17102__C1 _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18822_ _18822_/A _18822_/B _18822_/C _18822_/D vssd1 vssd1 vccd1 vccd1 _18822_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11157_ hold278/X _11126_/A fanout45/X hold316/A vssd1 vssd1 vccd1 vccd1 _11157_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13436__B _13875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18753_ _18752_/B _18906_/B _18752_/A vssd1 vssd1 vccd1 vccd1 _18754_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15965_ _15965_/A _15965_/B vssd1 vssd1 vccd1 vccd1 _15966_/C sky130_fd_sc_hd__xnor2_1
X_11088_ _10988_/Y hold6/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21683_/D sky130_fd_sc_hd__mux2_1
X_17704_ _17704_/A _17704_/B vssd1 vssd1 vccd1 vccd1 _17830_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_136_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14916_ _14916_/A _14916_/B vssd1 vssd1 vccd1 vccd1 _14918_/B sky130_fd_sc_hd__and2_2
XANTENNA__13155__C _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18684_ _18529_/B _18684_/B vssd1 vssd1 vccd1 vccd1 _18686_/B sky130_fd_sc_hd__and2b_2
X_15896_ _16028_/A _15896_/B vssd1 vssd1 vccd1 vccd1 _15898_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_78_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17635_ _17718_/A _17633_/X _17513_/B _17514_/Y vssd1 vssd1 vccd1 vccd1 _17694_/B
+ sky130_fd_sc_hd__o211a_1
X_14847_ _14848_/A _16173_/B _14848_/B _14848_/C vssd1 vssd1 vccd1 vccd1 _14847_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19123__B _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14548__A _14548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15431__A2 _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17566_ _17455_/A _17455_/C _17455_/B vssd1 vssd1 vccd1 vccd1 _17567_/C sky130_fd_sc_hd__a21bo_1
X_14778_ _14778_/A _14778_/B vssd1 vssd1 vccd1 vccd1 _14780_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19305_ _19143_/A _19143_/C _19143_/B vssd1 vssd1 vccd1 vccd1 _19307_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_128_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16517_ _16514_/X _16517_/B vssd1 vssd1 vccd1 vccd1 _16674_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_46_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13729_ _13729_/A _13729_/B vssd1 vssd1 vccd1 vccd1 _13732_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_86_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17497_ _17498_/A _17498_/B vssd1 vssd1 vccd1 vccd1 _17497_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_129_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17184__A2 _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19236_ _19088_/A _19090_/B _19088_/B vssd1 vssd1 vccd1 vccd1 _19241_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_45_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16448_ _16917_/C _16447_/X _16446_/X vssd1 vssd1 vccd1 vccd1 _16449_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_116_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20285__A _20689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19167_ _18396_/Y _19164_/X _19165_/Y _19166_/X vssd1 vssd1 vccd1 vccd1 _19167_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16379_ _16379_/A _16379_/B vssd1 vssd1 vccd1 vccd1 _16436_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_41_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19330__B1 _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18118_ _18119_/A _18119_/B vssd1 vssd1 vccd1 vccd1 _18118_/X sky130_fd_sc_hd__or2_1
XFILLER_0_41_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15098__B _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19098_ _19097_/A _19097_/B _19097_/C vssd1 vssd1 vccd1 vccd1 _19099_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_42_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18049_ _18787_/B _19089_/B _18773_/B _18787_/A vssd1 vssd1 vccd1 vccd1 _18049_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_83_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11508__A1 _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11508__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21060_ _21171_/A hold264/A vssd1 vssd1 vccd1 vccd1 _21061_/B sky130_fd_sc_hd__nand2_1
Xfanout405 _21768_/Q vssd1 vssd1 vccd1 vccd1 _13155_/D sky130_fd_sc_hd__clkbuf_8
XANTENNA__13049__D _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout416 _21766_/Q vssd1 vssd1 vccd1 vccd1 _15217_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout427 _21763_/Q vssd1 vssd1 vccd1 vccd1 _12781_/D sky130_fd_sc_hd__buf_4
X_20011_ _19911_/A _19911_/C _19911_/B vssd1 vssd1 vccd1 vccd1 _20012_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__20243__A2 _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout438 _14712_/A vssd1 vssd1 vccd1 vccd1 _14713_/A sky130_fd_sc_hd__buf_4
XFILLER_0_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout449 _12269_/A vssd1 vssd1 vccd1 vccd1 _12458_/A sky130_fd_sc_hd__buf_4
XANTENNA__20170__D _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout282_A _21799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16938__A _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21962_ _21963_/CLK _21962_/D vssd1 vssd1 vccd1 vccd1 hold250/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20913_ _20913_/A _20914_/B vssd1 vssd1 vccd1 vccd1 _20913_/Y sky130_fd_sc_hd__nand2_1
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21893_ _21932_/CLK hold105/X vssd1 vssd1 vccd1 vccd1 hold104/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout547_A _21734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20844_ _20844_/A _20844_/B vssd1 vssd1 vccd1 vccd1 _20849_/A sky130_fd_sc_hd__xnor2_2
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout12 _11446_/S vssd1 vssd1 vccd1 vccd1 _11470_/S sky130_fd_sc_hd__buf_6
XFILLER_0_92_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13984__A2 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout23 _11126_/Y vssd1 vssd1 vccd1 vccd1 fanout23/X sky130_fd_sc_hd__buf_4
XFILLER_0_76_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout34 _21490_/S vssd1 vssd1 vccd1 vccd1 _21507_/S sky130_fd_sc_hd__clkbuf_8
X_20775_ _20774_/A _20774_/B _21056_/B vssd1 vssd1 vccd1 vccd1 _20776_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout45 _11126_/B vssd1 vssd1 vccd1 vccd1 fanout45/X sky130_fd_sc_hd__buf_4
XFILLER_0_64_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout56 _10798_/Y vssd1 vssd1 vccd1 vccd1 _21261_/B sky130_fd_sc_hd__buf_4
XFILLER_0_130_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout67 _19181_/B vssd1 vssd1 vccd1 vccd1 _20841_/B sky130_fd_sc_hd__buf_4
XFILLER_0_119_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout78 _21847_/Q vssd1 vssd1 vccd1 vccd1 _19199_/D sky130_fd_sc_hd__buf_4
XFILLER_0_134_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout89 _18894_/B vssd1 vssd1 vccd1 vccd1 _19221_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14193__A _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12622__A1_N _12621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15439__D _15439_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21327_ hold187/X _11551_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _21327_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_4_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14697__B1 _14698_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12060_ _12229_/A _12246_/C _12246_/D _12155_/B vssd1 vssd1 vccd1 vccd1 _12061_/B
+ sky130_fd_sc_hd__a22o_1
X_21258_ _21258_/A _21258_/B vssd1 vssd1 vccd1 vccd1 _21259_/B sky130_fd_sc_hd__nand2_1
X_11011_ mstream_o[85] hold52/X _11012_/S vssd1 vssd1 vccd1 vccd1 _21622_/D sky130_fd_sc_hd__mux2_1
XANTENNA__16438__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20209_ _20210_/A _20210_/B vssd1 vssd1 vccd1 vccd1 _20209_/X sky130_fd_sc_hd__and2_1
X_21189_ _21296_/A _21286_/B _21296_/B _21291_/A vssd1 vssd1 vccd1 vccd1 _21191_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__11983__C _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13256__B _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15174__D _15174_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15750_ _15586_/A _15586_/B _15584_/Y vssd1 vssd1 vccd1 vccd1 _15752_/B sky130_fd_sc_hd__o21a_1
X_12962_ _12839_/X _12844_/A _13394_/A _14155_/C vssd1 vssd1 vccd1 vccd1 _13244_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_3321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13672__A1 _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14701_ _15375_/A _16268_/B _14702_/C _14702_/D vssd1 vssd1 vccd1 vccd1 _14701_/X
+ sky130_fd_sc_hd__and4_1
X_11913_ _12261_/A _12877_/B _12751_/B _12269_/B vssd1 vssd1 vccd1 vccd1 _11914_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20463__A2_N _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15681_ _15682_/A _15682_/B _15682_/C vssd1 vssd1 vccd1 vccd1 _15683_/B sky130_fd_sc_hd__a21o_2
XTAP_3365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_310 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ _12761_/X _12763_/X _12891_/Y _12892_/X vssd1 vssd1 vccd1 vccd1 _12895_/A
+ sky130_fd_sc_hd__o211ai_2
XTAP_3376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_321 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11491__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_332 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17420_ _17420_/A _17420_/B vssd1 vssd1 vccd1 vccd1 _17423_/A sky130_fd_sc_hd__xnor2_2
XTAP_3398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14632_ _14632_/A _14632_/B vssd1 vssd1 vccd1 vccd1 _14640_/A sky130_fd_sc_hd__nand2_1
X_11844_ _12458_/A _12443_/A _12877_/B _12357_/C vssd1 vssd1 vccd1 vccd1 _11845_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14563_ _14563_/A _14563_/B vssd1 vssd1 vccd1 vccd1 _14576_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_83_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17351_ _17351_/A _17351_/B _17351_/C vssd1 vssd1 vccd1 vccd1 _17351_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_36_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11775_ _12297_/B _11776_/B _11776_/C _11776_/D vssd1 vssd1 vccd1 vccd1 _11775_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_56_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16302_ _16302_/A _16302_/B vssd1 vssd1 vccd1 vccd1 _16344_/A sky130_fd_sc_hd__or2_1
XFILLER_0_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12319__C _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13514_ fanout9/X _21361_/B vssd1 vssd1 vccd1 vccd1 _13514_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14494_ _14494_/A _14494_/B vssd1 vssd1 vccd1 vccd1 _14496_/B sky130_fd_sc_hd__xnor2_4
X_17282_ _17282_/A _17741_/B vssd1 vssd1 vccd1 vccd1 _17286_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19021_ _19021_/A _19021_/B vssd1 vssd1 vccd1 vccd1 _19024_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_153_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16233_ _16302_/A _16232_/C _16232_/A vssd1 vssd1 vccd1 vccd1 _16233_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_126_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13445_ _13445_/A _13445_/B vssd1 vssd1 vccd1 vccd1 _13447_/B sky130_fd_sc_hd__or2_1
XFILLER_0_36_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12616__A _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16164_ _16164_/A _16275_/B vssd1 vssd1 vccd1 vccd1 _16167_/A sky130_fd_sc_hd__or2_1
X_13376_ _13376_/A _13376_/B vssd1 vssd1 vccd1 vccd1 _13386_/A sky130_fd_sc_hd__or2_1
XFILLER_0_2_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15115_ _16092_/D _15788_/B _15115_/C _15115_/D vssd1 vssd1 vccd1 vccd1 _15116_/B
+ sky130_fd_sc_hd__and4_1
X_12327_ _12637_/A _13155_/C _12326_/D _12750_/A vssd1 vssd1 vccd1 vccd1 _12328_/B
+ sky130_fd_sc_hd__a22o_1
X_16095_ _16095_/A _16211_/A _16095_/C vssd1 vssd1 vccd1 vccd1 _16207_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_107_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15046_ _14883_/X _14887_/C _15044_/Y _15045_/X vssd1 vssd1 vccd1 vccd1 _15046_/Y
+ sky130_fd_sc_hd__o211ai_4
X_19923_ _19923_/A _19923_/B _19921_/Y _19922_/X vssd1 vssd1 vccd1 vccd1 _19925_/A
+ sky130_fd_sc_hd__or4bb_1
X_12258_ _12258_/A _12258_/B _12258_/C vssd1 vssd1 vccd1 vccd1 _12275_/A sky130_fd_sc_hd__and3_1
X_11209_ hold161/X fanout22/X _11208_/X vssd1 vssd1 vccd1 vccd1 _11209_/X sky130_fd_sc_hd__a21o_1
X_19854_ _20088_/A _20249_/B _19854_/C _19950_/A vssd1 vssd1 vccd1 vccd1 _19950_/B
+ sky130_fd_sc_hd__nand4_1
X_12189_ _12223_/A _12269_/C vssd1 vssd1 vccd1 vccd1 _12191_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12351__A _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18805_ _18805_/A _18805_/B _18805_/C vssd1 vssd1 vccd1 vccd1 _18807_/B sky130_fd_sc_hd__nand3_1
XANTENNA__17861__B _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19785_ _19785_/A _19785_/B vssd1 vssd1 vccd1 vccd1 _19786_/B sky130_fd_sc_hd__nand2_1
X_16997_ _16997_/A _16997_/B vssd1 vssd1 vccd1 vccd1 _16999_/C sky130_fd_sc_hd__nor2_1
X_18736_ _19373_/B _19057_/C _19057_/D _19051_/A vssd1 vssd1 vccd1 vccd1 _18741_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12501__D _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15948_ _15948_/A _15948_/B _15948_/C vssd1 vssd1 vccd1 vccd1 _15948_/Y sky130_fd_sc_hd__nor3_4
XFILLER_0_116_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18667_ _18663_/X _18665_/Y _18511_/B _18511_/Y vssd1 vssd1 vccd1 vccd1 _18669_/D
+ sky130_fd_sc_hd__o211a_1
X_15879_ _15876_/X _15877_/Y _15737_/B _15738_/Y vssd1 vssd1 vccd1 vccd1 _15879_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_116_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16196__C _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16601__A1 _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17618_ _17618_/A _17618_/B vssd1 vssd1 vccd1 vccd1 _17627_/A sky130_fd_sc_hd__or2_1
XANTENNA__16601__B2 _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18598_ _19531_/A _19240_/B _18598_/C _18598_/D vssd1 vssd1 vccd1 vccd1 _18598_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_59_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17549_ _17550_/A _17550_/B vssd1 vssd1 vccd1 vccd1 _17652_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_50_1122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20560_ _21169_/A _21046_/B _21278_/B _21056_/A vssd1 vssd1 vccd1 vccd1 _20564_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_132_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17739__D _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19219_ _19076_/A _19076_/B _19076_/C _19078_/X vssd1 vssd1 vccd1 vccd1 _19252_/A
+ sky130_fd_sc_hd__a31o_1
X_20491_ _20491_/A _20491_/B _20491_/C vssd1 vssd1 vccd1 vccd1 _20492_/A sky130_fd_sc_hd__or3_2
XFILLER_0_144_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20462__B _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21112_ _20993_/Y _20997_/A _21109_/Y _21110_/X vssd1 vssd1 vccd1 vccd1 _21112_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22092_ _22096_/CLK _22092_/D _11089_/A vssd1 vssd1 vccd1 vccd1 mstream_o[28] sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout497_A _21745_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21413__A1 _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout202 _21817_/Q vssd1 vssd1 vccd1 vccd1 _20242_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_100_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21043_ _21267_/A _21841_/Q _21278_/B _21818_/Q vssd1 vssd1 vccd1 vccd1 _21161_/A
+ sky130_fd_sc_hd__and4_1
Xfanout213 _21283_/A vssd1 vssd1 vccd1 vccd1 _21153_/B sky130_fd_sc_hd__buf_4
Xfanout224 _18640_/B vssd1 vssd1 vccd1 vccd1 _19906_/C sky130_fd_sc_hd__buf_4
Xfanout235 _21809_/Q vssd1 vssd1 vccd1 vccd1 _17924_/B sky130_fd_sc_hd__buf_4
Xfanout246 _21807_/Q vssd1 vssd1 vccd1 vccd1 _21261_/A sky130_fd_sc_hd__buf_2
XFILLER_0_5_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17668__A1_N _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout257 hold322/X vssd1 vssd1 vccd1 vccd1 _18166_/A sky130_fd_sc_hd__buf_8
Xfanout268 _17417_/A vssd1 vssd1 vccd1 vccd1 _17526_/B sky130_fd_sc_hd__clkbuf_8
Xfanout279 _21799_/Q vssd1 vssd1 vccd1 vccd1 _17520_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15572__A _21740_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18586__C _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21293__B _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17490__C _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21724__D _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21945_ _21945_/CLK _21945_/D vssd1 vssd1 vccd1 vccd1 hold117/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17396__A2 _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21876_ _21945_/CLK hold110/X vssd1 vssd1 vccd1 vccd1 hold109/A sky130_fd_sc_hd__dfxtp_1
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20827_ _20824_/X _20825_/Y _20659_/Y _20661_/Y vssd1 vssd1 vccd1 vccd1 _20827_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17499__A _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14916__A _14916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12090__B1 _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11560_ _11557_/X _11560_/B vssd1 vssd1 vccd1 vccd1 _11815_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_64_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20758_ _20755_/Y _20756_/X _20628_/A _20627_/X vssd1 vssd1 vccd1 vccd1 _20758_/Y
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__18896__A2 _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14635__B _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout7_A fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13709__A2 _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_806 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11491_ _11490_/X _18616_/D _11521_/S vssd1 vssd1 vccd1 vccd1 _21835_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20689_ _20689_/A _21169_/A _21278_/B _21256_/B vssd1 vssd1 vccd1 vccd1 _20808_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_52_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14354__C _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13230_ _13230_/A _13230_/B vssd1 vssd1 vccd1 vccd1 _13249_/A sky130_fd_sc_hd__or2_1
XFILLER_0_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20653__A _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12155__B _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12393__A1 _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13161_ _13298_/B _13160_/B _13160_/C vssd1 vssd1 vccd1 vccd1 _13162_/C sky130_fd_sc_hd__a21o_1
XANTENNA__17856__B1 _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12393__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12112_ _12112_/A _12112_/B vssd1 vssd1 vccd1 vccd1 _12115_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_103_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13092_ _14294_/D _13092_/B vssd1 vssd1 vccd1 vccd1 _21352_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__17384__D _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16920_ _16920_/A _16920_/B _16920_/C vssd1 vssd1 vccd1 vccd1 _16973_/A sky130_fd_sc_hd__nand3_1
X_12043_ _12043_/A _12043_/B _12043_/C vssd1 vssd1 vccd1 vccd1 _12050_/A sky130_fd_sc_hd__nand3_1
X_16851_ _16851_/A _16851_/B _16851_/C vssd1 vssd1 vccd1 vccd1 _16859_/A sky130_fd_sc_hd__nand3_2
XANTENNA__15095__B1 _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15634__A2 _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15802_ _15802_/A _15802_/B vssd1 vssd1 vccd1 vccd1 _15813_/A sky130_fd_sc_hd__or2_1
XFILLER_0_137_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19570_ _20394_/B _19866_/D _19874_/B _19972_/A vssd1 vssd1 vccd1 vccd1 _19575_/C
+ sky130_fd_sc_hd__a22o_1
X_16782_ _16783_/A _16783_/B _16783_/C vssd1 vssd1 vccd1 vccd1 _16789_/A sky130_fd_sc_hd__a21oi_2
X_13994_ _14306_/A _14138_/A _14477_/C _14635_/D _13839_/X vssd1 vssd1 vccd1 vccd1
+ _14002_/A sky130_fd_sc_hd__a41o_1
XFILLER_0_137_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18521_ _18521_/A _18521_/B _18521_/C _18521_/D vssd1 vssd1 vccd1 vccd1 _18521_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_73_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15733_ _15733_/A _15733_/B _15733_/C vssd1 vssd1 vccd1 vccd1 _15733_/X sky130_fd_sc_hd__or3_2
XTAP_3140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12945_ _12961_/B _12945_/B _12945_/C vssd1 vssd1 vccd1 vccd1 _13091_/A sky130_fd_sc_hd__nand3_4
XFILLER_0_133_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15632__D _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18452_ _18453_/A _18453_/B _18453_/C vssd1 vssd1 vccd1 vccd1 _18454_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_34_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15664_ _15665_/A _15665_/B vssd1 vssd1 vccd1 vccd1 _15862_/A sky130_fd_sc_hd__nand2b_1
XTAP_3195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12876_ _13858_/A _13012_/B vssd1 vssd1 vccd1 vccd1 _12880_/A sky130_fd_sc_hd__nand2_1
XANTENNA_140 v1z[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_151 v1z[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17403_ _17404_/A _17404_/B _17404_/C vssd1 vssd1 vccd1 vccd1 _17405_/B sky130_fd_sc_hd__a21oi_4
XANTENNA_162 v2z[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14615_ _15159_/D _14936_/D _15954_/D vssd1 vssd1 vccd1 vccd1 _14615_/X sky130_fd_sc_hd__and3_1
XFILLER_0_96_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_173 v2z[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_184 hold239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18383_ _18125_/Y _18128_/Y _18380_/Y _18381_/X vssd1 vssd1 vccd1 vccd1 _18385_/A
+ sky130_fd_sc_hd__a211o_1
X_11827_ _11794_/X _11824_/Y _11823_/Y _11823_/A vssd1 vssd1 vccd1 vccd1 _11830_/C
+ sky130_fd_sc_hd__o211ai_4
X_15595_ _15596_/B _15596_/A vssd1 vssd1 vccd1 vccd1 _15595_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__17139__A2 _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15441__A1_N _15439_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_195 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19533__B1 _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20547__B _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17334_ _17657_/A _17334_/B _17666_/A _17443_/D vssd1 vssd1 vccd1 vccd1 _17335_/B
+ sky130_fd_sc_hd__and4_1
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14546_ _14546_/A _14690_/A _14546_/C vssd1 vssd1 vccd1 vccd1 _14690_/B sky130_fd_sc_hd__nand3_2
X_11758_ _11758_/A _11758_/B _11758_/C vssd1 vssd1 vccd1 vccd1 _11784_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_28_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12620__A2 _13269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12991__D _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16463__D _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17265_ _17265_/A _17265_/B vssd1 vssd1 vccd1 vccd1 _17267_/B sky130_fd_sc_hd__xnor2_4
X_14477_ _15153_/B _15155_/C _14477_/C _14635_/D vssd1 vssd1 vccd1 vccd1 _14632_/A
+ sky130_fd_sc_hd__nand4_2
X_11689_ _14621_/D _12319_/C _12420_/D _12403_/A vssd1 vssd1 vccd1 vccd1 _11690_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19004_ hold97/X _19003_/X fanout4/X vssd1 vssd1 vccd1 vccd1 hold98/A sky130_fd_sc_hd__mux2_1
XFILLER_0_10_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16216_ _16323_/A vssd1 vssd1 vccd1 vccd1 _16218_/D sky130_fd_sc_hd__inv_2
XFILLER_0_144_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13428_ _13428_/A _13428_/B _13415_/Y vssd1 vssd1 vccd1 vccd1 _13428_/Y sky130_fd_sc_hd__nor3b_4
X_17196_ _17196_/A _17196_/B vssd1 vssd1 vccd1 vccd1 _17198_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__18639__A2 _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16147_ hold76/X _16146_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _21882_/D sky130_fd_sc_hd__mux2_1
X_13359_ _13218_/B _13218_/Y _13509_/B _13358_/X vssd1 vssd1 vccd1 vccd1 _13512_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_23_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21378__B _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17311__A2 _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18033__A _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16078_ _16078_/A _16078_/B _16078_/C vssd1 vssd1 vccd1 vccd1 _16079_/C sky130_fd_sc_hd__and3_1
XFILLER_0_87_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15029_ _15029_/A _15029_/B vssd1 vssd1 vccd1 vccd1 _15037_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17872__A _18008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19906_ _19906_/A _20146_/B _19906_/C _19906_/D vssd1 vssd1 vccd1 vccd1 _20001_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12512__C _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19837_ _19837_/A _19837_/B vssd1 vssd1 vccd1 vccd1 _19840_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19768_ _19768_/A _19768_/B vssd1 vssd1 vccd1 vccd1 _19769_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18719_ _18720_/A _18720_/B _18720_/C vssd1 vssd1 vccd1 vccd1 _18719_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__13624__B _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19699_ _19699_/A _19699_/B vssd1 vssd1 vccd1 vccd1 _19715_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21730_ _22020_/CLK _21730_/D vssd1 vssd1 vccd1 vccd1 _21730_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21661_ _21934_/CLK _21661_/D vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout245_A _21261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clk_i_A clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20612_ _20613_/A _20613_/B vssd1 vssd1 vccd1 vccd1 _20612_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19030__C _19030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21592_ _21888_/CLK _21592_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[55] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12611__A2 _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13997__D _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20543_ _20991_/C _21264_/A _20544_/C _20730_/A vssd1 vssd1 vccd1 vccd1 _20545_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14364__A2 _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20474_ _21199_/A _21283_/B _21305_/B _20838_/B vssd1 vssd1 vccd1 vccd1 _20478_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17302__A2 _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16510__B1 _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15717__D _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14621__D _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22075_ _22080_/CLK _22075_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[11] sky130_fd_sc_hd__dfrtp_4
X_21026_ _21138_/A _21026_/B vssd1 vssd1 vccd1 vccd1 _21027_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_156_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15077__B1 _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13815__A fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16829__C _17141_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout60_A _21407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11638__B1 _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10991_ mstream_o[65] hold72/X _21568_/S vssd1 vssd1 vccd1 vccd1 _21602_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12730_ _12730_/A _12730_/B vssd1 vssd1 vccd1 vccd1 _12731_/B sky130_fd_sc_hd__xor2_4
X_21928_ _21932_/CLK _21928_/D vssd1 vssd1 vccd1 vccd1 hold136/A sky130_fd_sc_hd__dfxtp_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16041__A2 _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10861__A1 _10860_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12661_ _13155_/B _12771_/C _21765_/Q _13018_/B vssd1 vssd1 vccd1 vccd1 _12661_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21859_ _21923_/CLK _21859_/D vssd1 vssd1 vccd1 vccd1 hold227/A sky130_fd_sc_hd__dfxtp_1
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19221__B _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18318__A1 _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18318__B2 _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14400_ _14224_/B _14226_/B _14397_/X _14399_/Y vssd1 vssd1 vccd1 vccd1 _14402_/A
+ sky130_fd_sc_hd__a211o_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _11612_/A _11612_/B vssd1 vssd1 vccd1 vccd1 _11897_/A sky130_fd_sc_hd__nor2_1
XANTENNA__17022__A _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15380_ _15380_/A _15380_/B vssd1 vssd1 vccd1 vccd1 _15382_/B sky130_fd_sc_hd__xor2_2
X_12592_ _12415_/X _12418_/Y _12589_/X _12590_/Y vssd1 vssd1 vccd1 vccd1 _12592_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14365__B _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14331_ _14331_/A _14331_/B _14331_/C vssd1 vssd1 vccd1 vccd1 _14333_/B sky130_fd_sc_hd__nand3_2
XANTENNA__20676__A2 _21040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11543_ _11089_/B t1y[31] t0x[31] _11543_/B2 vssd1 vssd1 vccd1 vccd1 _11543_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_52_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16861__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14084__C _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14262_ _14101_/B _14101_/Y _14260_/X _14261_/Y vssd1 vssd1 vccd1 vccd1 _14264_/B
+ sky130_fd_sc_hd__a211o_1
X_17050_ _17049_/B _17117_/A _17005_/Y _17008_/X vssd1 vssd1 vccd1 vccd1 _17050_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_68_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11474_ _11498_/A1 t1y[8] t0x[8] _11501_/B2 vssd1 vssd1 vccd1 vccd1 _11474_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_151_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16001_ _15826_/Y _15874_/X _15999_/Y _16000_/X vssd1 vssd1 vccd1 vccd1 _16001_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_122_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13213_ _13213_/A _13213_/B _13213_/C vssd1 vssd1 vccd1 vccd1 _13213_/Y sky130_fd_sc_hd__nand3_4
XANTENNA__20814__C _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14193_ _14365_/A _14367_/A _14516_/A _14365_/C vssd1 vssd1 vccd1 vccd1 _14362_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_151_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17395__C _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13144_ _13029_/B _13031_/A _13142_/X _13143_/Y vssd1 vssd1 vccd1 vccd1 _13230_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_21_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ _12931_/X _12934_/X _13072_/X _13073_/Y vssd1 vssd1 vccd1 vccd1 _13077_/B
+ sky130_fd_sc_hd__o211ai_1
X_17952_ _17953_/A _17953_/B _17953_/C vssd1 vssd1 vccd1 vccd1 _17952_/Y sky130_fd_sc_hd__nor3_2
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17057__A1 _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21418__S _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16903_ _16903_/A _16903_/B _16903_/C vssd1 vssd1 vccd1 vccd1 _16958_/A sky130_fd_sc_hd__nand3_1
X_12026_ _12077_/A _12077_/B vssd1 vssd1 vccd1 vccd1 _12029_/B sky130_fd_sc_hd__or2_1
XANTENNA__17057__B2 _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11877__B1 _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17883_ _17883_/A _17883_/B _17883_/C vssd1 vssd1 vccd1 vccd1 _17884_/A sky130_fd_sc_hd__and3_1
X_19622_ _19461_/A _19461_/B _19459_/Y vssd1 vssd1 vccd1 vccd1 _19624_/B sky130_fd_sc_hd__a21oi_1
X_16834_ _16836_/A _16836_/B vssd1 vssd1 vccd1 vccd1 _16834_/Y sky130_fd_sc_hd__nand2_1
X_19553_ _19395_/A _19395_/C _19395_/B vssd1 vssd1 vccd1 vccd1 _19554_/C sky130_fd_sc_hd__a21bo_1
X_16765_ _16765_/A _16765_/B vssd1 vssd1 vccd1 vccd1 _16838_/A sky130_fd_sc_hd__xor2_2
X_13977_ _13974_/Y _14142_/A _14312_/D _16409_/B vssd1 vssd1 vccd1 vccd1 _14142_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18504_ _18503_/A _18503_/B _18503_/C vssd1 vssd1 vccd1 vccd1 _18505_/C sky130_fd_sc_hd__a21o_1
X_15716_ _15719_/D vssd1 vssd1 vccd1 vccd1 _15716_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12928_ _12929_/A _12929_/B _12929_/C vssd1 vssd1 vccd1 vccd1 _12928_/Y sky130_fd_sc_hd__nor3_1
X_19484_ _19366_/A _19366_/B _19364_/Y vssd1 vssd1 vccd1 vccd1 _19526_/A sky130_fd_sc_hd__o21ba_1
X_16696_ _17096_/A _16917_/C _16444_/A _16442_/Y vssd1 vssd1 vccd1 vccd1 _16697_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_75_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18435_ _18435_/A _18588_/B vssd1 vssd1 vccd1 vccd1 _18438_/A sky130_fd_sc_hd__or2_1
X_15647_ _16151_/A _15647_/B vssd1 vssd1 vccd1 vccd1 _15648_/C sky130_fd_sc_hd__xnor2_1
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ _13858_/B _13269_/C _13269_/D _13860_/A vssd1 vssd1 vccd1 vccd1 _12860_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18028__A _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19506__B1 _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18366_ _18362_/X _18364_/Y _18215_/B _18215_/Y vssd1 vssd1 vccd1 vccd1 _18368_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15578_ _15578_/A _15578_/B vssd1 vssd1 vccd1 vccd1 _15582_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17317_ _17317_/A _17317_/B _17317_/C vssd1 vssd1 vccd1 vccd1 _17317_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_44_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14529_ _14526_/X _14527_/Y _14398_/Y _14402_/A vssd1 vssd1 vccd1 vccd1 _14530_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18297_ _18294_/Y _18442_/A _20317_/D _19240_/B vssd1 vssd1 vccd1 vccd1 _18442_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_3_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17248_ _17248_/A _17248_/B _17248_/C vssd1 vssd1 vccd1 vccd1 _17251_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_3_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17179_ _17741_/B _17387_/A _16543_/B _16541_/X vssd1 vssd1 vccd1 vccd1 _17188_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13619__B _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20190_ _20975_/D _20733_/C _20606_/D _20845_/D vssd1 vssd1 vccd1 vccd1 _20190_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__13857__A1 _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13857__B2 _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12242__C _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout195_A _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13872__A4 _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15553__C _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15963__A1_N _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13609__A1 _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout362_A _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19745__B1 _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20862__A2_N _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16559__B1 _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21713_ _22105_/CLK _21713_/D vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfxtp_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14034__A1 _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14034__B2 _21742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout627_A _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21644_ _21722_/CLK hold289/X fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[107]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12045__B1 _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_40 _11436_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21575_ mstream_o[38] _11057_/Y _21579_/S vssd1 vssd1 vccd1 vccd1 _22102_/D sky130_fd_sc_hd__mux2_1
XANTENNA_51 hold275/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17523__A2 _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_62 hold274/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_73 hold268/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20526_ _20397_/A _20396_/B _20650_/B vssd1 vssd1 vccd1 vccd1 _20526_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_133_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_84 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_95 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12136__D _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20457_ _20590_/D _21291_/B _20458_/C _20458_/D vssd1 vssd1 vccd1 vccd1 _20459_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13529__B _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11190_ hold302/X fanout51/X fanout47/X hold280/X vssd1 vssd1 vccd1 vccd1 _11190_/X
+ sky130_fd_sc_hd__a22o_1
X_20388_ _20774_/A _20774_/B _21256_/B _21258_/B vssd1 vssd1 vccd1 vccd1 _20559_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_24_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22058_ _22063_/CLK _22058_/D vssd1 vssd1 vccd1 vccd1 hold274/A sky130_fd_sc_hd__dfxtp_4
XFILLER_0_100_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13900_ _13901_/A _13901_/B _13901_/C vssd1 vssd1 vccd1 vccd1 _13900_/Y sky130_fd_sc_hd__a21oi_1
X_21009_ _21005_/X _21006_/Y _20826_/Y _20830_/B vssd1 vssd1 vccd1 vccd1 _21009_/X
+ sky130_fd_sc_hd__a211o_1
X_14880_ _14877_/X _14878_/Y _14699_/Y _14701_/X vssd1 vssd1 vccd1 vccd1 _14881_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11991__C _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13831_ _13831_/A _13831_/B vssd1 vssd1 vccd1 vccd1 _13833_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_97_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18539__B2 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16550_ _17197_/B _16550_/B vssd1 vssd1 vccd1 vccd1 _16552_/B sky130_fd_sc_hd__xnor2_1
X_13762_ _14848_/A _13913_/C _13622_/B _13620_/X vssd1 vssd1 vccd1 vccd1 _13767_/A
+ sky130_fd_sc_hd__a31o_1
X_10974_ _10972_/A _10971_/A _10971_/B vssd1 vssd1 vccd1 vccd1 _10978_/A sky130_fd_sc_hd__a21bo_2
XANTENNA__19200__A2 _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16575__B _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15501_ _15501_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _15907_/A sky130_fd_sc_hd__nor2_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12713_ hold203/X _12712_/X fanout3/X vssd1 vssd1 vccd1 vccd1 _21858_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14025__A1 _14659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16481_ _17041_/A _17019_/C _17123_/C _16899_/B vssd1 vssd1 vccd1 vccd1 _16482_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18493__D _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13693_ _13689_/A _13690_/X _13534_/A _13535_/Y vssd1 vssd1 vccd1 vccd1 _13693_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_84_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19495__A2_N _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18220_ _18220_/A _18220_/B _18220_/C _18220_/D vssd1 vssd1 vccd1 vccd1 _18220_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_66_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15432_ _15838_/D _15702_/D _15829_/C _15954_/D vssd1 vssd1 vccd1 vccd1 _15577_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_84_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12644_ _13013_/A _13155_/C _13155_/D _12877_/A vssd1 vssd1 vccd1 vccd1 _12645_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16970__B1 _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18151_ _18293_/B _18150_/C _18150_/A vssd1 vssd1 vccd1 vccd1 _18152_/C sky130_fd_sc_hd__o21ai_2
X_15363_ _15363_/A _15502_/B vssd1 vssd1 vccd1 vccd1 _15365_/B sky130_fd_sc_hd__xor2_1
X_12575_ _12575_/A _12575_/B _12575_/C vssd1 vssd1 vccd1 vccd1 _12578_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_0_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16591__A _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17102_ _17094_/B _17096_/X _17029_/A _17146_/D vssd1 vssd1 vccd1 vccd1 _17110_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_123_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14314_ _14312_/D _16406_/B _16374_/B _14133_/D vssd1 vssd1 vccd1 vccd1 _14315_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_18082_ _18082_/A _18082_/B _18082_/C vssd1 vssd1 vccd1 vccd1 _18082_/X sky130_fd_sc_hd__or3_2
X_11526_ _11544_/A1 t2x[25] v1z[25] fanout21/X _11525_/X vssd1 vssd1 vccd1 vccd1 _11526_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15294_ _15291_/Y _15292_/X _15147_/B _15146_/X vssd1 vssd1 vccd1 vccd1 _15295_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_123_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17033_ _17033_/A _17033_/B vssd1 vssd1 vccd1 vccd1 _17035_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_68_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14245_ _14245_/A _14245_/B vssd1 vssd1 vccd1 vccd1 _14255_/A sky130_fd_sc_hd__xor2_1
X_11457_ _21718_/D t2x[2] v1z[2] fanout18/X _11456_/X vssd1 vssd1 vccd1 vccd1 _11457_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_111_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14176_ _15435_/A _15153_/B _14176_/C vssd1 vssd1 vccd1 vccd1 _14176_/X sky130_fd_sc_hd__and3_1
XFILLER_0_22_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11388_ hold261/X fanout29/X _11387_/X vssd1 vssd1 vccd1 vccd1 _11388_/X sky130_fd_sc_hd__a21o_1
XANTENNA__20841__A _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15828__A2 _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13127_ _13127_/A _13127_/B vssd1 vssd1 vccd1 vccd1 _13142_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18949__C _19753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18984_ _19007_/B _18983_/B _18981_/X _18982_/Y vssd1 vssd1 vccd1 vccd1 _18984_/X
+ sky130_fd_sc_hd__a2bb2o_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ _12918_/A _12918_/C _12918_/B vssd1 vssd1 vccd1 vccd1 _13059_/C sky130_fd_sc_hd__a21bo_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17935_ _17935_/A _17935_/B _17935_/C vssd1 vssd1 vccd1 vccd1 _17937_/B sky130_fd_sc_hd__nand3_2
XANTENNA__18030__B _18030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20034__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12009_ _12009_/A _12009_/B vssd1 vssd1 vccd1 vccd1 _12011_/B sky130_fd_sc_hd__xor2_1
X_17866_ _17867_/B _17867_/A vssd1 vssd1 vccd1 vccd1 _17982_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__20585__A1 _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16817_ _17096_/A _17013_/C _16803_/X _16733_/X _16968_/C vssd1 vssd1 vccd1 vccd1
+ _16820_/A sky130_fd_sc_hd__a32o_1
X_19605_ _19604_/B _19729_/B _19604_/A vssd1 vssd1 vccd1 vccd1 _19606_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_75_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17797_ _17797_/A _17797_/B _17797_/C vssd1 vssd1 vccd1 vccd1 _17799_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_36_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19536_ _19686_/A _20419_/A _19538_/C _19538_/D vssd1 vssd1 vccd1 vccd1 _19536_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21534__A0 hold268/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16748_ _17096_/A _16968_/C _16736_/B _16734_/X vssd1 vssd1 vccd1 vccd1 _16751_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17202__A1 _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17202__B2 _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19467_ _19467_/A _19467_/B _19467_/C vssd1 vssd1 vccd1 vccd1 _19468_/B sky130_fd_sc_hd__nand3_1
X_16679_ _16652_/X _16677_/Y _16676_/Y _16676_/A vssd1 vssd1 vccd1 vccd1 _16682_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18950__A1 _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18418_ _18264_/X _18266_/Y _18415_/Y _18417_/X vssd1 vssd1 vccd1 vccd1 _18543_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_9_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19398_ _19398_/A _19398_/B _19398_/C vssd1 vssd1 vccd1 vccd1 _19400_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18349_ _19445_/A _19866_/D vssd1 vssd1 vccd1 vccd1 _18352_/A sky130_fd_sc_hd__and2_1
XFILLER_0_133_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20735__B _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21360_ hold190/X fanout40/X _21358_/Y _21359_/Y vssd1 vssd1 vccd1 vccd1 _21927_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11250__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11250__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20311_ _20462_/D _21291_/B _20312_/C _20312_/D vssd1 vssd1 vccd1 vccd1 _20313_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_25_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21291_ _21291_/A _21291_/B vssd1 vssd1 vccd1 vccd1 _21295_/A sky130_fd_sc_hd__nand2_1
XANTENNA_fanout110_A _19692_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout208_A _19753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18466__B1 _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20242_ _20774_/A _20774_/B _20242_/C _20242_/D vssd1 vssd1 vccd1 vccd1 _20428_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_40_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20173_ _20317_/D _20841_/B _20173_/C _20173_/D vssd1 vssd1 vccd1 vccd1 _20314_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__17763__C _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20025__B1 _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout577_A _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__A1 _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19966__B1 _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__B2 _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15452__B1 _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17992__A2 _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21525__A0 hold275/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11613__A _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14558__A2 _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout23_A _11126_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21627_ _21682_/CLK _21627_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[90] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15507__A1 _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17300__A _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11241__A1 _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12360_ _12359_/B _12359_/C _12359_/A vssd1 vssd1 vccd1 vccd1 _12362_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_145_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11241__B2 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21558_ mstream_o[21] hold26/X _21562_/S vssd1 vssd1 vccd1 vccd1 _22085_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_62_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15507__B2 _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11311_ fanout58/X v0z[21] fanout17/X _11310_/X vssd1 vssd1 vccd1 vccd1 _11311_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17657__D _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_15_clk_i _21806_/CLK vssd1 vssd1 vccd1 vccd1 _21817_/CLK sky130_fd_sc_hd__clkbuf_16
X_20509_ _20363_/A _20367_/A _20639_/B _20508_/X vssd1 vssd1 vccd1 vccd1 _20509_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_132_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12291_ _16363_/A _12291_/B vssd1 vssd1 vccd1 vccd1 fanout6/A sky130_fd_sc_hd__nor2_2
X_21489_ hold176/X sstream_i[66] _21489_/S vssd1 vssd1 vccd1 vccd1 _22016_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12444__A _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14030_ _14028_/X _14030_/B vssd1 vssd1 vccd1 vccd1 _14031_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_132_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11242_ _21718_/D t1x[4] v2z[4] _21724_/D _11241_/X vssd1 vssd1 vccd1 vccd1 _11242_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_28_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20264__B1 _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19227__A _19379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11173_ hold153/X fanout23/X _11172_/X vssd1 vssd1 vccd1 vccd1 _11173_/X sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_7_clk_i_A _21806_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18131__A _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16483__A2 _17141_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15981_ _15981_/A _15981_/B vssd1 vssd1 vccd1 vccd1 _15983_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11494__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17720_ _17854_/B _18857_/B _19051_/C _18894_/B vssd1 vssd1 vccd1 vccd1 _17720_/X
+ sky130_fd_sc_hd__and4_1
X_14932_ _14934_/A _14934_/B _14934_/C vssd1 vssd1 vccd1 vccd1 _14935_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__18797__A1_N _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17651_ _17652_/A _17652_/B _17652_/C vssd1 vssd1 vccd1 vccd1 _17651_/X sky130_fd_sc_hd__a21o_4
X_14863_ _14862_/B _14862_/C _14862_/A vssd1 vssd1 vccd1 vccd1 _14865_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_72_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16602_ _18166_/A _17666_/A _17443_/D _17434_/B vssd1 vssd1 vccd1 vccd1 _16603_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_98_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13814_ _13814_/A _13814_/B vssd1 vssd1 vccd1 vccd1 _18689_/B sky130_fd_sc_hd__xor2_4
X_17582_ _17468_/Y _17470_/X _17579_/X _17581_/Y vssd1 vssd1 vccd1 vccd1 _17584_/B
+ sky130_fd_sc_hd__a211o_1
X_14794_ _14793_/B _14793_/C _14793_/A vssd1 vssd1 vccd1 vccd1 _14795_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_98_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20319__B2 _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19321_ _19319_/X _19321_/B vssd1 vssd1 vccd1 vccd1 _19788_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_97_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16533_ _16532_/A _16532_/B _16532_/C vssd1 vssd1 vccd1 vccd1 _16534_/C sky130_fd_sc_hd__a21o_1
X_13745_ _14195_/A _14537_/A vssd1 vssd1 vccd1 vccd1 _13746_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13722__B _13877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10957_ _10957_/A _10957_/B vssd1 vssd1 vccd1 vccd1 _10959_/B sky130_fd_sc_hd__or2_2
XFILLER_0_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12619__A _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19252_ _19252_/A _19252_/B _19252_/C vssd1 vssd1 vccd1 vccd1 _19254_/A sky130_fd_sc_hd__and3_1
X_16464_ _17206_/B _17124_/C vssd1 vssd1 vccd1 vccd1 _16478_/A sky130_fd_sc_hd__nand2_1
X_13676_ _13676_/A _13676_/B vssd1 vssd1 vccd1 vccd1 _13677_/B sky130_fd_sc_hd__and2_1
XANTENNA__11480__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10888_ hold216/A hold217/A vssd1 vssd1 vccd1 vccd1 _10890_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_155_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18203_ _18498_/B _19866_/D _19874_/B _18652_/A vssd1 vssd1 vccd1 vccd1 _18204_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15415_ _15415_/A _15415_/B vssd1 vssd1 vccd1 vccd1 _15417_/B sky130_fd_sc_hd__xnor2_1
X_19183_ _19179_/C _19013_/X _19016_/A _19016_/B vssd1 vssd1 vccd1 vccd1 _19184_/B
+ sky130_fd_sc_hd__o2bb2a_2
X_12627_ _12627_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _12629_/C sky130_fd_sc_hd__xnor2_1
X_16395_ _16316_/A _16315_/A _16400_/A _16312_/B vssd1 vssd1 vccd1 vccd1 _16434_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18134_ _18134_/A _18134_/B vssd1 vssd1 vccd1 vccd1 _18143_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_5_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11232__A1 _11231_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15346_ _15346_/A _15346_/B vssd1 vssd1 vccd1 vccd1 _15347_/B sky130_fd_sc_hd__or2_2
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12558_ _12558_/A _12558_/B vssd1 vssd1 vccd1 vccd1 _12578_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_124_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11509_ _11508_/X _19227_/D _11521_/S vssd1 vssd1 vccd1 vccd1 _21841_/D sky130_fd_sc_hd__mux2_1
X_18065_ _18498_/B _19414_/C _19866_/D _18652_/A vssd1 vssd1 vccd1 vccd1 _18066_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15277_ _15277_/A _15406_/B vssd1 vssd1 vccd1 vccd1 _15279_/B sky130_fd_sc_hd__or2_2
Xhold107 hold107/A vssd1 vssd1 vccd1 vccd1 hold107/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12489_ _11907_/A _12387_/B _12708_/A vssd1 vssd1 vccd1 vccd1 _12490_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_112_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold118 hold118/A vssd1 vssd1 vccd1 vccd1 hold118/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_145_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold129 hold129/A vssd1 vssd1 vccd1 vccd1 hold129/X sky130_fd_sc_hd__dlygate4sd3_1
X_17016_ _17016_/A _17016_/B _17016_/C vssd1 vssd1 vccd1 vccd1 _17068_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_151_594 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14228_ _14228_/A _14228_/B _14228_/C vssd1 vssd1 vccd1 vccd1 _14230_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_21_250 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14159_ _14156_/Y _14157_/X _14020_/D _14021_/B vssd1 vssd1 vccd1 vccd1 _14160_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_1_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout609 _21718_/Q vssd1 vssd1 vccd1 vccd1 _11507_/A1 sky130_fd_sc_hd__buf_2
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20721__D _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13288__A2 _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18967_ _18967_/A _18967_/B _18967_/C vssd1 vssd1 vccd1 vccd1 _18969_/B sky130_fd_sc_hd__nand3_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13185__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17918_ _21087_/D _18789_/A _18047_/A _17917_/D vssd1 vssd1 vccd1 vccd1 _17919_/C
+ sky130_fd_sc_hd__a22o_1
X_18898_ _19382_/A _19230_/A _19240_/B _19057_/C vssd1 vssd1 vccd1 vccd1 _18901_/D
+ sky130_fd_sc_hd__nand4_1
X_17849_ _17850_/A _17850_/B vssd1 vssd1 vccd1 vccd1 _17990_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16496__A _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13913__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20860_ _20863_/D vssd1 vssd1 vccd1 vccd1 _20860_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_95_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13996__B1 _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19519_ _19519_/A _19519_/B vssd1 vssd1 vccd1 vccd1 _19521_/B sky130_fd_sc_hd__nor2_1
X_20791_ _20924_/A _21301_/A _21305_/A _21151_/A vssd1 vssd1 vccd1 vccd1 _20794_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13460__A2 _14212_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout158_A _21830_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11471__A1 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11471__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12248__B _21727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17758__C _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21412_ _21412_/A _21412_/B vssd1 vssd1 vccd1 vccd1 _21412_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__22066__RESET_B fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14463__B _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21343_ _21349_/A _21343_/B vssd1 vssd1 vccd1 vccd1 _21343_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_142_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16162__A1 _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20847__A1_N _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21274_ _21274_/A _21274_/B vssd1 vssd1 vccd1 vccd1 _21280_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19692__D _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20246__B1 _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13920__B1 _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15575__A _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20225_ _20224_/A _20224_/B _20224_/C vssd1 vssd1 vccd1 vccd1 _20226_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_12_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16465__A2 _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20156_ _20156_/A _20156_/B vssd1 vssd1 vccd1 vccd1 _20157_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__14476__A1 _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12711__B _21343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14476__B2 _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21630__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20087_ _20087_/A _20087_/B vssd1 vssd1 vccd1 vccd1 _20093_/A sky130_fd_sc_hd__nand2_1
XANTENNA__20549__A1 _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16217__A2 _21784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17414__A1 _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21210__A2 _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11860_ _12109_/C _12621_/C vssd1 vssd1 vccd1 vccd1 _11936_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10811_ hold107/A hold104/A vssd1 vssd1 vccd1 vccd1 _10843_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17014__B _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11791_ _11791_/A _11791_/B _11791_/C vssd1 vssd1 vccd1 vccd1 _11795_/A sky130_fd_sc_hd__nand3_4
XTAP_2879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20989_ _21296_/A _21286_/A _21283_/B _21305_/B vssd1 vssd1 vccd1 vccd1 _21096_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_67_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13530_ _13822_/B _16328_/B _13528_/Y _13678_/A vssd1 vssd1 vccd1 vccd1 _13530_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_83_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11462__A1 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11462__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13461_ _15217_/A _14212_/C _13461_/C _13461_/D vssd1 vssd1 vccd1 vccd1 _13608_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15200_ _15200_/A _15200_/B vssd1 vssd1 vccd1 vccd1 _15201_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_36_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12412_ _12413_/A _12413_/B vssd1 vssd1 vccd1 vccd1 _12412_/X sky130_fd_sc_hd__and2b_1
X_16180_ _16287_/A _16180_/B vssd1 vssd1 vccd1 vccd1 _16181_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13392_ _13393_/A _13393_/B vssd1 vssd1 vccd1 vccd1 _13392_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_51_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15131_ _15933_/C _16328_/A _15129_/Y _15271_/A vssd1 vssd1 vccd1 vccd1 _15133_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__16153__A1 _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12343_ _12444_/B _12877_/A _12897_/C _12897_/D vssd1 vssd1 vccd1 vccd1 _12343_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__16153__B2 _16391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21029__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15062_ _15063_/A _15063_/B vssd1 vssd1 vccd1 vccd1 _15203_/A sky130_fd_sc_hd__or2_1
X_12274_ _12258_/B _12258_/C _12258_/A vssd1 vssd1 vccd1 vccd1 _12275_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__12714__A1 _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14013_ _13886_/Y _13889_/Y _14131_/B _14012_/X vssd1 vssd1 vccd1 vccd1 _14015_/B
+ sky130_fd_sc_hd__a211o_1
X_11225_ _11122_/A t2y[0] t0y[0] _11123_/A vssd1 vssd1 vccd1 vccd1 _11225_/X sky130_fd_sc_hd__a22o_1
XANTENNA__17102__B1 _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19870_ _20394_/B _19872_/C _19972_/C _19972_/A vssd1 vssd1 vccd1 vccd1 _19874_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21718__RESET_B _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18821_ _18822_/A _18822_/B _18822_/C _18822_/D vssd1 vssd1 vccd1 vccd1 _18821_/Y
+ sky130_fd_sc_hd__nor4_2
X_11156_ _12751_/B _11155_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21735_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_156_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18752_ _18752_/A _18752_/B _18906_/B vssd1 vssd1 vccd1 vccd1 _18752_/X sky130_fd_sc_hd__and3_1
X_15964_ _15964_/A _15964_/B vssd1 vssd1 vccd1 vccd1 _15965_/B sky130_fd_sc_hd__nor2_1
X_11087_ _10984_/Y hold46/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21682_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13436__C _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17703_ _17703_/A _17703_/B vssd1 vssd1 vccd1 vccd1 _17704_/B sky130_fd_sc_hd__xnor2_4
X_14915_ _14608_/A _14757_/Y _14912_/Y _14603_/B _14756_/Y vssd1 vssd1 vccd1 vccd1
+ _14916_/B sky130_fd_sc_hd__a221oi_4
X_18683_ _18683_/A _18683_/B vssd1 vssd1 vccd1 vccd1 _18686_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11150__A0 _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15895_ _16027_/A _16380_/B vssd1 vssd1 vccd1 vccd1 _15896_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_136_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13155__D _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17634_ _17513_/B _17514_/Y _17718_/A _17633_/X vssd1 vssd1 vccd1 vccd1 _17718_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_72_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14846_ _14846_/A _14846_/B vssd1 vssd1 vccd1 vccd1 _14893_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_72_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19123__C _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17565_ _17564_/B _17564_/C _17564_/A vssd1 vssd1 vccd1 vccd1 _17567_/B sky130_fd_sc_hd__a21o_1
X_14777_ _14777_/A _14777_/B vssd1 vssd1 vccd1 vccd1 _14778_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_59_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11989_ _11989_/A _11989_/B _11989_/C vssd1 vssd1 vccd1 vccd1 _11996_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_128_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19304_ _19304_/A _19304_/B vssd1 vssd1 vccd1 vccd1 _19307_/A sky130_fd_sc_hd__xnor2_2
X_16516_ _16564_/B _16513_/X _16507_/X _16668_/A vssd1 vssd1 vccd1 vccd1 _16517_/B
+ sky130_fd_sc_hd__a211o_1
X_13728_ _13729_/A _13729_/B vssd1 vssd1 vccd1 vccd1 _13883_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_105_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11453__A1 _21718_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17496_ _17388_/A _17388_/B _17386_/A vssd1 vssd1 vccd1 vccd1 _17498_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__11453__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19235_ _19235_/A _19235_/B vssd1 vssd1 vccd1 vccd1 _19243_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_129_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16447_ _16813_/A _17029_/B _16968_/C vssd1 vssd1 vccd1 vccd1 _16447_/X sky130_fd_sc_hd__and3_1
XFILLER_0_27_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13659_ _13656_/Y _13657_/X _13504_/X _13508_/A vssd1 vssd1 vccd1 vccd1 _13660_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_128_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20285__B _20562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19166_ _19000_/A _19000_/B _18836_/Y _18838_/Y vssd1 vssd1 vccd1 vccd1 _19166_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16378_ _16378_/A _16378_/B vssd1 vssd1 vccd1 vccd1 _16379_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18117_ _18117_/A _18117_/B vssd1 vssd1 vccd1 vccd1 _18119_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__19330__B2 _19650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15329_ _15177_/B _15179_/B _15327_/Y _15328_/X vssd1 vssd1 vccd1 vccd1 _15332_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_53_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19097_ _19097_/A _19097_/B _19097_/C vssd1 vssd1 vccd1 vccd1 _19099_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_152_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18048_ _17928_/A _17927_/B _17927_/A vssd1 vssd1 vccd1 vccd1 _18055_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout406 _15514_/B vssd1 vssd1 vccd1 vccd1 _15373_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20010_ _20154_/A _20009_/C _20009_/A vssd1 vssd1 vccd1 vccd1 _20012_/B sky130_fd_sc_hd__a21o_1
XANTENNA__17644__A1 _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout417 _12897_/D vssd1 vssd1 vccd1 vccd1 _12155_/B sky130_fd_sc_hd__buf_4
XANTENNA__18202__C _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout428 _14716_/A vssd1 vssd1 vccd1 vccd1 _14848_/A sky130_fd_sc_hd__buf_4
XANTENNA__14458__A1 _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout439 _21761_/Q vssd1 vssd1 vccd1 vccd1 _14712_/A sky130_fd_sc_hd__buf_4
X_19999_ _19999_/A _19999_/B vssd1 vssd1 vccd1 vccd1 _20000_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16938__B _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21961_ _21963_/CLK _21961_/D vssd1 vssd1 vccd1 vccd1 hold318/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11141__A0 _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout275_A _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20912_ _20912_/A _20912_/B vssd1 vssd1 vccd1 vccd1 _20914_/B sky130_fd_sc_hd__xor2_4
X_21892_ _21926_/CLK _21892_/D vssd1 vssd1 vccd1 vccd1 hold80/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20843_ _20843_/A _20843_/B vssd1 vssd1 vccd1 vccd1 _20844_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_7_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20590__A_N _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11444__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout13 wire16/A vssd1 vssd1 vccd1 vccd1 _11446_/S sky130_fd_sc_hd__buf_6
X_20774_ _20774_/A _20774_/B _21056_/B vssd1 vssd1 vccd1 vccd1 _20776_/A sky130_fd_sc_hd__and3_1
Xfanout24 _11260_/S vssd1 vssd1 vccd1 vccd1 _11195_/S sky130_fd_sc_hd__clkbuf_8
Xfanout35 _21490_/S vssd1 vssd1 vccd1 vccd1 _21510_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20476__A _21261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout46 fanout49/X vssd1 vssd1 vccd1 vccd1 _11126_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout57 _10797_/Y vssd1 vssd1 vccd1 vccd1 _16374_/B sky130_fd_sc_hd__buf_4
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout68 hold325/X vssd1 vssd1 vccd1 vccd1 _19181_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_130_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout79 _20606_/D vssd1 vssd1 vccd1 vccd1 _21305_/B sky130_fd_sc_hd__buf_4
XFILLER_0_134_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14193__B _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21326_ _11550_/A _21324_/Y _21325_/X vssd1 vssd1 vccd1 vccd1 _21326_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_130_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14697__A1 _21768_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14697__B2 _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21257_ _21257_/A _21257_/B vssd1 vssd1 vccd1 vccd1 _21260_/A sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout90_A _21844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11010_ mstream_o[84] hold14/X _11012_/S vssd1 vssd1 vccd1 vccd1 _21621_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18112__C _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20208_ _20208_/A _20208_/B vssd1 vssd1 vccd1 vccd1 _20210_/B sky130_fd_sc_hd__xnor2_1
X_21188_ _21188_/A _21188_/B vssd1 vssd1 vccd1 vccd1 _21230_/A sky130_fd_sc_hd__or2_2
XFILLER_0_25_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11983__D _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20139_ _20139_/A _20275_/B _20140_/B vssd1 vssd1 vccd1 vccd1 _20343_/A sky130_fd_sc_hd__or3b_1
XTAP_3300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11132__A0 _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ _12961_/A _12961_/B vssd1 vssd1 vccd1 vccd1 _13088_/A sky130_fd_sc_hd__nand2_2
XTAP_3311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14700_ _15375_/A _16268_/B _14702_/C _14702_/D vssd1 vssd1 vccd1 vccd1 _14700_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11912_ _12268_/A _12637_/B vssd1 vssd1 vccd1 vccd1 _11914_/B sky130_fd_sc_hd__and2_1
X_15680_ _15680_/A _15680_/B vssd1 vssd1 vccd1 vccd1 _15682_/C sky130_fd_sc_hd__xnor2_1
XTAP_3355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_300 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ _13010_/B _12891_/C _12891_/A vssd1 vssd1 vccd1 vccd1 _12892_/X sky130_fd_sc_hd__a21o_1
XTAP_3366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_311 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_322 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_333 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14631_ _14512_/A _14511_/B _14509_/X vssd1 vssd1 vccd1 vccd1 _14631_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _12268_/A _12751_/B vssd1 vssd1 vccd1 vccd1 _11845_/B sky130_fd_sc_hd__and2_1
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_620 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11435__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17350_ _17351_/A _17351_/B _17351_/C vssd1 vssd1 vccd1 vccd1 _17350_/X sky130_fd_sc_hd__and3_1
X_14562_ _14560_/X _14562_/B vssd1 vssd1 vccd1 vccd1 _14563_/B sky130_fd_sc_hd__and2b_1
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ _11752_/X _11754_/Y _11772_/A _11772_/Y vssd1 vssd1 vccd1 vccd1 _11776_/D
+ sky130_fd_sc_hd__o211a_2
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16301_ _16301_/A _16301_/B vssd1 vssd1 vccd1 vccd1 _16345_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_95_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13513_ _13513_/A _13518_/D vssd1 vssd1 vccd1 vccd1 _21361_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_27_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17281_ _17281_/A _17281_/B vssd1 vssd1 vccd1 vccd1 _17288_/A sky130_fd_sc_hd__or2_1
XANTENNA__12319__D _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14384__A _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14493_ _14494_/B _14494_/A vssd1 vssd1 vccd1 vccd1 _14611_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_126_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19020_ _19021_/A _19021_/B vssd1 vssd1 vccd1 vccd1 _19190_/B sky130_fd_sc_hd__nor2_1
X_16232_ _16232_/A _16302_/A _16232_/C vssd1 vssd1 vccd1 vccd1 _16302_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_67_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13444_ _13444_/A _13444_/B vssd1 vssd1 vccd1 vccd1 _13447_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_24_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12616__B _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16163_ _16273_/A _16414_/B _16163_/C _16163_/D vssd1 vssd1 vccd1 vccd1 _16275_/B
+ sky130_fd_sc_hd__and4_1
X_13375_ _13266_/A _13265_/B _13265_/A vssd1 vssd1 vccd1 vccd1 _13388_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_24_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15114_ _16092_/D _15788_/B _15115_/C _15115_/D vssd1 vssd1 vccd1 vccd1 _15116_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__14137__B1 _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12326_ _12637_/A _12750_/A _13155_/C _12326_/D vssd1 vssd1 vccd1 vccd1 _12326_/X
+ sky130_fd_sc_hd__and4_1
X_16094_ _16211_/A _16095_/C _16095_/A vssd1 vssd1 vccd1 vccd1 _16096_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_121_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15045_ _15044_/B _15044_/C _15044_/A vssd1 vssd1 vccd1 vccd1 _15045_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19922_ _19919_/X _19920_/Y _19712_/Y _19714_/X vssd1 vssd1 vccd1 vccd1 _19922_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_107_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12257_ _12256_/A _12256_/B _12256_/C vssd1 vssd1 vccd1 vccd1 _12258_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11208_ hold220/X fanout51/X fanout48/X hold238/A vssd1 vssd1 vccd1 vccd1 _11208_/X
+ sky130_fd_sc_hd__a22o_1
X_12188_ _12199_/A _12188_/B vssd1 vssd1 vccd1 vccd1 _12191_/A sky130_fd_sc_hd__nor2_1
X_19853_ _19432_/A _20249_/B _19854_/C _19950_/A vssd1 vssd1 vccd1 vccd1 _19855_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12351__B _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18804_ _18653_/A _18653_/B _18653_/C vssd1 vssd1 vccd1 vccd1 _18805_/C sky130_fd_sc_hd__a21bo_1
X_11139_ hold249/A _11126_/A fanout45/X hold165/X vssd1 vssd1 vccd1 vccd1 _11139_/X
+ sky130_fd_sc_hd__a22o_1
X_16996_ _17041_/A _17493_/A _18859_/A _16899_/B vssd1 vssd1 vccd1 vccd1 _16997_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__17861__C _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19784_ _19785_/A _19785_/B vssd1 vssd1 vccd1 vccd1 _19796_/A sky130_fd_sc_hd__or2_1
X_15947_ _15944_/Y _15945_/X _15816_/B _15817_/Y vssd1 vssd1 vccd1 vccd1 _15948_/C
+ sky130_fd_sc_hd__o211a_1
X_18735_ _18735_/A _18735_/B vssd1 vssd1 vccd1 vccd1 _18745_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__14559__A _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18666_ _18511_/B _18511_/Y _18663_/X _18665_/Y vssd1 vssd1 vccd1 vccd1 _18669_/C
+ sky130_fd_sc_hd__a211oi_4
X_15878_ _15737_/B _15738_/Y _15876_/X _15877_/Y vssd1 vssd1 vccd1 vccd1 _15878_/Y
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__16601__A2 _17666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16196__D _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14829_ _15808_/C _16404_/A _14830_/C _15029_/A vssd1 vssd1 vccd1 vccd1 _14831_/B
+ sky130_fd_sc_hd__a22o_1
X_17617_ _17617_/A _17617_/B vssd1 vssd1 vccd1 vccd1 _17630_/A sky130_fd_sc_hd__xor2_2
X_18597_ _19531_/A _19240_/B _18598_/C _18598_/D vssd1 vssd1 vccd1 vccd1 _18597_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_54_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11426__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17548_ _17548_/A _17548_/B vssd1 vssd1 vccd1 vccd1 _17550_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17479_ _17479_/A _17479_/B vssd1 vssd1 vccd1 vccd1 _17593_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_73_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19218_ _19218_/A _19218_/B vssd1 vssd1 vccd1 vccd1 _19308_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_144_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20490_ _20487_/Y _20488_/X _20342_/X _20344_/X vssd1 vssd1 vccd1 vccd1 _20491_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19149_ _19148_/B _19148_/C _19148_/A vssd1 vssd1 vccd1 vccd1 _19149_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12245__C _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21111_ _20993_/Y _20997_/A _21109_/Y _21110_/X vssd1 vssd1 vccd1 vccd1 _21111_/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__20462__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19067__B1 _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22091_ _22105_/CLK _22091_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[27] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21042_ _21841_/Q _21278_/B _21818_/Q _21267_/A vssd1 vssd1 vccd1 vccd1 _21046_/C
+ sky130_fd_sc_hd__a22o_1
Xfanout203 _21817_/Q vssd1 vssd1 vccd1 vccd1 _19872_/C sky130_fd_sc_hd__buf_4
Xfanout214 hold332/X vssd1 vssd1 vccd1 vccd1 _21283_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_34_clk_i_A clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout392_A _15892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout225 _20270_/C vssd1 vssd1 vccd1 vccd1 _18640_/B sky130_fd_sc_hd__buf_4
Xfanout236 _20991_/C vssd1 vssd1 vccd1 vccd1 _21291_/A sky130_fd_sc_hd__buf_4
Xfanout247 _21807_/Q vssd1 vssd1 vccd1 vccd1 _17915_/A sky130_fd_sc_hd__buf_4
Xfanout258 _21803_/Q vssd1 vssd1 vccd1 vccd1 _17434_/B sky130_fd_sc_hd__clkbuf_8
Xfanout269 _19051_/A vssd1 vssd1 vccd1 vccd1 _20462_/D sky130_fd_sc_hd__buf_4
XANTENNA__18586__D _19060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11114__A0 _10946_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17490__D _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21944_ _21945_/CLK _21944_/D vssd1 vssd1 vccd1 vccd1 hold124/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19790__A1 _19169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21875_ _21939_/CLK _21875_/D vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19060__A _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11417__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20826_ _20659_/Y _20661_/Y _20824_/X _20825_/Y vssd1 vssd1 vccd1 vccd1 _20826_/Y
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__17499__B _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19995__A _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20757_ _20628_/A _20627_/X _20755_/Y _20756_/X vssd1 vssd1 vccd1 vccd1 _20757_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_134_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15564__C1 _15386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11490_ _11493_/A1 t2x[13] v1z[13] fanout20/X _11489_/X vssd1 vssd1 vccd1 vccd1 _11490_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20688_ _20691_/D vssd1 vssd1 vccd1 vccd1 _20688_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_45_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21101__A1 _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18404__A _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12155__C _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20653__B _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13590__A1 _13875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17856__A1 _18851_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13160_ _13298_/B _13160_/B _13160_/C vssd1 vssd1 vccd1 vccd1 _13287_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_62_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17856__B2 _17854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14651__B _14652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12111_ _12112_/B _12112_/A vssd1 vssd1 vccd1 vccd1 _12120_/B sky130_fd_sc_hd__and2b_1
X_21309_ _21309_/A _21309_/B vssd1 vssd1 vccd1 vccd1 _21310_/B sky130_fd_sc_hd__xnor2_1
X_13091_ _13091_/A _13091_/B vssd1 vssd1 vccd1 vccd1 _13518_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12452__A _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12042_ _11986_/A _11986_/C _11986_/B vssd1 vssd1 vccd1 vccd1 _12043_/C sky130_fd_sc_hd__a21o_1
Xhold290 hold290/A vssd1 vssd1 vccd1 vccd1 hold290/X sky130_fd_sc_hd__buf_4
XANTENNA__11353__B1 _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15763__A _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16850_ _16855_/A _16850_/B vssd1 vssd1 vccd1 vccd1 _16851_/C sky130_fd_sc_hd__and2_1
XANTENNA__15095__A1 _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15801_ _15986_/B _15801_/B vssd1 vssd1 vccd1 vccd1 _15816_/A sky130_fd_sc_hd__and2_1
XANTENNA__15095__B2 _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16831__A2 _17141_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16781_ _16781_/A _16781_/B vssd1 vssd1 vccd1 vccd1 _16783_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__11105__A0 _10881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13993_ _13871_/A _13870_/B _13868_/X vssd1 vssd1 vccd1 vccd1 _13993_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18520_ _18521_/A _18521_/B _18521_/C _18521_/D vssd1 vssd1 vccd1 vccd1 _18520_/Y
+ sky130_fd_sc_hd__nor4_1
X_15732_ _15733_/A _15733_/B _15733_/C vssd1 vssd1 vccd1 vccd1 _15732_/Y sky130_fd_sc_hd__nor3_1
XTAP_3130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12944_ _12818_/A _12818_/C _12818_/B vssd1 vssd1 vccd1 vccd1 _12945_/C sky130_fd_sc_hd__o21bai_2
XTAP_3141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16044__B1 _21753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18451_ _18451_/A _18451_/B vssd1 vssd1 vccd1 vccd1 _18453_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_38_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15663_ _15663_/A _15663_/B vssd1 vssd1 vccd1 vccd1 _15665_/B sky130_fd_sc_hd__or2_1
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_130 v1z[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12875_ _12778_/A _12777_/B _12775_/X vssd1 vssd1 vccd1 vccd1 _12891_/A sky130_fd_sc_hd__a21o_1
XTAP_3196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_141 v1z[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17402_ _17402_/A _17402_/B vssd1 vssd1 vccd1 vccd1 _17404_/C sky130_fd_sc_hd__xnor2_2
XANTENNA_152 v1z[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14614_ _15159_/D _15829_/C _15954_/D _14936_/D vssd1 vssd1 vccd1 vccd1 _14614_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11408__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18382_ _18125_/Y _18128_/Y _18380_/Y _18381_/X vssd1 vssd1 vccd1 vccd1 _18382_/Y
+ sky130_fd_sc_hd__a211oi_2
XANTENNA_163 v2z[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11826_ _11830_/B vssd1 vssd1 vccd1 vccd1 _11826_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_68_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15594_ _15594_/A _15713_/B vssd1 vssd1 vccd1 vccd1 _15596_/B sky130_fd_sc_hd__or2_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_174 v2z[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_185 hold239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_196 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19533__A1 _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17333_ _17657_/A _17666_/A _17443_/D _17334_/B vssd1 vssd1 vccd1 vccd1 _17335_/A
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__19533__B2 _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20547__C _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14545_ _14542_/Y _14543_/X _14391_/D _14393_/B vssd1 vssd1 vccd1 vccd1 _14546_/C
+ sky130_fd_sc_hd__o211ai_2
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ _12261_/A _13157_/A _13017_/A _12269_/B vssd1 vssd1 vccd1 vccd1 _11758_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17544__B1 _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17264_ _17264_/A _17264_/B vssd1 vssd1 vccd1 vccd1 _17265_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_153_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14476_ _15153_/B _14477_/C _14635_/D _15155_/C vssd1 vssd1 vccd1 vccd1 _14479_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11688_ _14621_/D _12319_/C _12420_/D _12403_/A vssd1 vssd1 vccd1 vccd1 _11688_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_125_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19003_ hold191/A fanout7/X _14126_/X _11550_/B _19002_/Y vssd1 vssd1 vccd1 vccd1
+ _19003_/X sky130_fd_sc_hd__a221o_1
XANTENNA__12908__A1 _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16215_ _16328_/A _16326_/A _16396_/B _16418_/B vssd1 vssd1 vccd1 vccd1 _16323_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_148_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_829 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13427_ _13427_/A _13427_/B _13427_/C vssd1 vssd1 vccd1 vccd1 _13428_/B sky130_fd_sc_hd__and3_1
XFILLER_0_36_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17195_ _17196_/A _17196_/B vssd1 vssd1 vccd1 vccd1 _17195_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_24_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18314__A _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1203 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16146_ _16363_/A hold77/X _10972_/Y fanout5/X _16145_/Y vssd1 vssd1 vccd1 vccd1
+ _16146_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_11_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13358_ _13509_/A _13357_/C _13357_/A vssd1 vssd1 vccd1 vccd1 _13358_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18033__B _19379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13458__A _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12309_ _12310_/A _12310_/B vssd1 vssd1 vccd1 vccd1 _12309_/Y sky130_fd_sc_hd__nor2_1
X_16077_ _16078_/A _16078_/B _16078_/C vssd1 vssd1 vccd1 vccd1 _16077_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_80_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13289_ _13875_/B _14024_/B _14384_/A _14212_/B vssd1 vssd1 vccd1 vccd1 _13290_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_20_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15028_ _15028_/A _15028_/B vssd1 vssd1 vccd1 vccd1 _15044_/A sky130_fd_sc_hd__xnor2_2
X_19905_ _20146_/B _19906_/C _19906_/D _19906_/A vssd1 vssd1 vccd1 vccd1 _19908_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17872__B _18010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11344__A0 _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15673__A _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12512__D _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19836_ _19833_/X _19834_/Y _19671_/X _19673_/Y vssd1 vssd1 vccd1 vccd1 _19837_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_120_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19767_ _19768_/B _19768_/A vssd1 vssd1 vccd1 vccd1 _19767_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_127_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16979_ _16973_/A _16973_/B _16973_/C vssd1 vssd1 vccd1 vccd1 _16980_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_39_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11706__A _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18718_ _18718_/A _18718_/B vssd1 vssd1 vccd1 vccd1 _18720_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19698_ _19696_/X _19698_/B vssd1 vssd1 vccd1 vccd1 _19699_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_91_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18649_ _18649_/A _18649_/B vssd1 vssd1 vccd1 vccd1 _18658_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_8_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13921__A _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21660_ _21934_/CLK _21660_/D vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20611_ _20611_/A _20611_/B vssd1 vssd1 vccd1 vccd1 _20613_/B sky130_fd_sc_hd__xnor2_1
X_21591_ _21888_/CLK _21591_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[54] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_145_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_1084 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19030__D _21847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout238_A _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20542_ _21296_/A _21286_/A _21151_/A _21301_/A vssd1 vssd1 vccd1 vccd1 _20730_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_116_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20473_ _20473_/A _20473_/B vssd1 vssd1 vccd1 vccd1 _20481_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_104_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout405_A _21768_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16510__A1 _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16510__B2 _16743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22074_ _22080_/CLK _22074_/D fanout639/X vssd1 vssd1 vccd1 vccd1 mstream_o[10] sky130_fd_sc_hd__dfrtp_4
XANTENNA__11335__B1 _11334_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21025_ _21138_/B _21025_/B vssd1 vssd1 vccd1 vccd1 _21027_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20477__A2_N _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15077__A1 _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13815__B _18689_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16829__D _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18894__A _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11638__A1 _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11616__A _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11638__B2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10990_ mstream_o[64] hold59/X _10992_/S vssd1 vssd1 vccd1 vccd1 _21601_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_97_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21927_ _21932_/CLK _21927_/D vssd1 vssd1 vccd1 vccd1 hold190/A sky130_fd_sc_hd__dfxtp_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21570__A1 _11045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ _14195_/A _13018_/B _21765_/Q vssd1 vssd1 vccd1 vccd1 _12660_/X sky130_fd_sc_hd__and3_1
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19221__C _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21858_ _21926_/CLK _21858_/D vssd1 vssd1 vccd1 vccd1 hold203/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18318__A2 _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11611_ _11601_/X _11609_/X _11610_/Y _11833_/A vssd1 vssd1 vccd1 vccd1 _11833_/B
+ sky130_fd_sc_hd__o211ai_4
X_20809_ _20910_/A hold264/A _20656_/A _20654_/B vssd1 vssd1 vccd1 vccd1 _20817_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17022__B _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14772__A1_N _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12591_ _12415_/X _12418_/Y _12589_/X _12590_/Y vssd1 vssd1 vccd1 vccd1 _12591_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_26_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21789_ _21789_/CLK _21789_/D vssd1 vssd1 vccd1 vccd1 hold319/A sky130_fd_sc_hd__dfxtp_4
XFILLER_0_19_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14365__C _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14330_ _14329_/B _14474_/B _14329_/A vssd1 vssd1 vccd1 vccd1 _14331_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_93_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11542_ _11541_/X _19185_/B _11545_/S vssd1 vssd1 vccd1 vccd1 _21852_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_65_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14261_ _14260_/B _14260_/C _14260_/A vssd1 vssd1 vccd1 vccd1 _14261_/Y sky130_fd_sc_hd__a21oi_2
X_11473_ _11472_/X _18787_/B _11521_/S vssd1 vssd1 vccd1 vccd1 _21829_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14662__A _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16000_ _15999_/A _15999_/B _15999_/C _15999_/D vssd1 vssd1 vccd1 vccd1 _16000_/X
+ sky130_fd_sc_hd__o22a_1
X_13212_ _13209_/X _13210_/Y _13072_/B _13071_/Y vssd1 vssd1 vccd1 vccd1 _13213_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_21_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14192_ _21743_/Q _14516_/A _14365_/C _14367_/A vssd1 vssd1 vccd1 vccd1 _14195_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17395__D _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11497__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13143_ _13142_/B _13142_/C _13142_/A vssd1 vssd1 vccd1 vccd1 _13143_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_108_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13074_ _12931_/X _12934_/X _13072_/X _13073_/Y vssd1 vssd1 vccd1 vccd1 _13074_/X
+ sky130_fd_sc_hd__o211a_1
X_17951_ _17948_/X _17949_/Y _17810_/B _17809_/Y vssd1 vssd1 vccd1 vccd1 _17953_/C
+ sky130_fd_sc_hd__a211oi_2
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17057__A2 _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16902_ _16823_/X _16891_/Y _16890_/Y _16890_/A vssd1 vssd1 vccd1 vccd1 _16903_/C
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__18254__A1 _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12025_ _12029_/A _12025_/B vssd1 vssd1 vccd1 vccd1 _12077_/B sky130_fd_sc_hd__nand2_1
X_17882_ _17881_/A _17881_/B _17881_/C vssd1 vssd1 vccd1 vccd1 _17883_/C sky130_fd_sc_hd__a21o_1
XANTENNA__18254__B2 _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11877__A1 _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12910__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11877__B2 _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16265__B1 _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19621_ _19621_/A _19621_/B vssd1 vssd1 vccd1 vccd1 _19624_/A sky130_fd_sc_hd__xor2_1
X_16833_ _16833_/A _16898_/A vssd1 vssd1 vccd1 vccd1 _16836_/B sky130_fd_sc_hd__or2_1
XFILLER_0_75_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14815__B2 _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16764_ _16765_/A _16765_/B vssd1 vssd1 vccd1 vccd1 _16764_/X sky130_fd_sc_hd__and2_1
X_19552_ _19551_/B _19551_/C _19551_/A vssd1 vssd1 vccd1 vccd1 _19554_/B sky130_fd_sc_hd__a21o_1
X_13976_ _13682_/C _16409_/B _13974_/Y _14142_/A vssd1 vssd1 vccd1 vccd1 _13980_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16106__A2_N _21784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15715_ _15717_/B _15717_/C _15976_/D _16084_/A vssd1 vssd1 vccd1 vccd1 _15719_/D
+ sky130_fd_sc_hd__a22o_1
X_18503_ _18503_/A _18503_/B _18503_/C vssd1 vssd1 vccd1 vccd1 _18505_/B sky130_fd_sc_hd__nand3_1
X_12927_ _12923_/X _12925_/Y _12798_/B _12798_/Y vssd1 vssd1 vccd1 vccd1 _12929_/C
+ sky130_fd_sc_hd__o211a_1
X_16695_ _16694_/A _16694_/C _16694_/B vssd1 vssd1 vccd1 vccd1 _16698_/B sky130_fd_sc_hd__a21o_1
X_19483_ _19483_/A _19483_/B vssd1 vssd1 vccd1 vccd1 _19626_/A sky130_fd_sc_hd__or2_1
XFILLER_0_38_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15646_ _16036_/A _15647_/B vssd1 vssd1 vccd1 vccd1 _15782_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_115_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18434_ _18431_/Y _18588_/A _19487_/A _19382_/B vssd1 vssd1 vccd1 vccd1 _18588_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_87_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12858_ _13858_/B _13860_/A _12858_/C _13269_/D vssd1 vssd1 vccd1 vccd1 _12989_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_69_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19506__A1 _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18028__B _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19506__B2 _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18365_ _18215_/B _18215_/Y _18362_/X _18364_/Y vssd1 vssd1 vccd1 vccd1 _18368_/C
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__12054__A1 _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11809_ _12458_/A _12444_/B _12443_/A _12357_/C vssd1 vssd1 vccd1 vccd1 _11810_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_145_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15577_ _15577_/A _15577_/B vssd1 vssd1 vccd1 vccd1 _15578_/B sky130_fd_sc_hd__nor2_2
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12789_ _12676_/A _12676_/C _12676_/B vssd1 vssd1 vccd1 vccd1 _12790_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_84_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17316_ _17317_/A _17317_/B _17317_/C vssd1 vssd1 vccd1 vccd1 _17316_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14528_ _14398_/Y _14402_/A _14526_/X _14527_/Y vssd1 vssd1 vccd1 vccd1 _14530_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18296_ _20317_/D _19240_/B _18294_/Y _18442_/A vssd1 vssd1 vccd1 vccd1 _18296_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17247_ _16617_/A _16617_/C _16617_/B vssd1 vssd1 vccd1 vccd1 _17248_/C sky130_fd_sc_hd__a21bo_1
X_14459_ _14621_/D _15698_/B vssd1 vssd1 vccd1 vccd1 _14460_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_4_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14572__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17178_ _17178_/A _17178_/B vssd1 vssd1 vccd1 vccd1 _17196_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_141_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16129_ _16128_/A _16128_/B _16128_/C vssd1 vssd1 vccd1 vccd1 _16129_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_109_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19690__B1 _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18698__B _19181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13857__A2 _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12242__D _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19819_ _19699_/A _19698_/B _19696_/X vssd1 vssd1 vccd1 vccd1 _19830_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13609__A2 _14873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout188_A _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19603__A _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19745__A1 _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19745__B2 _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16559__A1 _16813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16559__B2 _16743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17123__A _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21712_ _22105_/CLK _21712_/D vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14034__A2 _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21643_ _21722_/CLK hold300/X fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[106]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_fanout522_A _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21304__A1 _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12267__A _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18257__A2_N _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_30 _11343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21574_ mstream_o[37] _11055_/Y _21579_/S vssd1 vssd1 vccd1 vccd1 _22101_/D sky130_fd_sc_hd__mux2_1
XANTENNA_41 _11445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_52 hold275/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_63 hold274/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20525_ _20249_/A _21056_/B _20396_/B vssd1 vssd1 vccd1 vccd1 _20657_/A sky130_fd_sc_hd__a21oi_1
XANTENNA_74 hold277/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_85 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_96 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20456_ _20588_/A vssd1 vssd1 vccd1 vccd1 _20458_/D sky130_fd_sc_hd__inv_2
XFILLER_0_127_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20387_ _20774_/B _21256_/B _21258_/B _20774_/A vssd1 vssd1 vccd1 vccd1 _20390_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13529__C _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11308__A0 _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22057_ _22063_/CLK _22057_/D vssd1 vssd1 vccd1 vccd1 hold288/A sky130_fd_sc_hd__dfxtp_4
X_21008_ _21008_/A vssd1 vssd1 vccd1 vccd1 _21008_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11991__D _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13830_ _13831_/A _13831_/B vssd1 vssd1 vccd1 vccd1 _13992_/B sky130_fd_sc_hd__or2_1
XFILLER_0_138_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18539__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13761_ _14557_/A _14557_/B _14218_/B _14391_/B _13614_/B vssd1 vssd1 vccd1 vccd1
+ _13770_/A sky130_fd_sc_hd__a41o_1
X_10973_ mstream_o[60] _10972_/Y _11005_/S vssd1 vssd1 vccd1 vccd1 _21597_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_134_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15500_ hold79/X _15499_/X fanout4/X vssd1 vssd1 vccd1 vccd1 _21877_/D sky130_fd_sc_hd__mux2_1
X_12712_ _21725_/D hold60/X _11053_/X fanout6/X _12711_/Y vssd1 vssd1 vccd1 vccd1
+ _12712_/X sky130_fd_sc_hd__a221o_1
X_16480_ _17206_/B _17141_/C vssd1 vssd1 vccd1 vccd1 _16758_/A sky130_fd_sc_hd__nand2_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13692_ _13534_/A _13535_/Y _13689_/A _13690_/X vssd1 vssd1 vccd1 vccd1 _13692_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA_clkbuf_leaf_3_clk_i_A _21822_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15431_ _14813_/A _15829_/C _15954_/D _15702_/D vssd1 vssd1 vccd1 vccd1 _15435_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17968__A _17969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12643_ _13013_/A _12877_/A _13155_/C _13155_/D vssd1 vssd1 vccd1 vccd1 _12643_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_109_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18150_ _18150_/A _18293_/B _18150_/C vssd1 vssd1 vccd1 vccd1 _18304_/A sky130_fd_sc_hd__or3_4
XFILLER_0_65_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15362_ _15362_/A _15362_/B vssd1 vssd1 vccd1 vccd1 _15502_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_108_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12574_ _12465_/A _12465_/C _12465_/B vssd1 vssd1 vccd1 vccd1 _12575_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__20394__A _21831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17101_ _17101_/A _17101_/B _17101_/C vssd1 vssd1 vccd1 vccd1 _17106_/A sky130_fd_sc_hd__and3_1
XANTENNA__16591__B _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14313_ _14315_/A vssd1 vssd1 vccd1 vccd1 _14471_/A sky130_fd_sc_hd__inv_2
XFILLER_0_0_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18081_ _18082_/A _18082_/B _18082_/C vssd1 vssd1 vccd1 vccd1 _18081_/Y sky130_fd_sc_hd__nor3_1
X_11525_ _11089_/B t1y[25] t0x[25] _11223_/A vssd1 vssd1 vccd1 vccd1 _11525_/X sky130_fd_sc_hd__a22o_1
X_15293_ _15147_/B _15146_/X _15291_/Y _15292_/X vssd1 vssd1 vccd1 vccd1 _15295_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_123_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12905__A _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17032_ _16989_/C _17146_/D _16990_/A _16988_/Y vssd1 vssd1 vccd1 vccd1 _17033_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14244_ _14848_/A _15098_/B vssd1 vssd1 vccd1 vccd1 _14245_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_123_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11456_ _11123_/A t1y[2] t0x[2] _21724_/D vssd1 vssd1 vccd1 vccd1 _11456_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_145_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18799__A _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14175_ _15435_/A _14176_/C _15112_/D _15153_/B vssd1 vssd1 vccd1 vccd1 _14175_/X
+ sky130_fd_sc_hd__a22o_1
X_11387_ _11124_/A hold244/X fanout45/X hold211/X vssd1 vssd1 vccd1 vccd1 _11387_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20841__B _20841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12343__C _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13126_ _13126_/A _13126_/B vssd1 vssd1 vccd1 vccd1 _13127_/B sky130_fd_sc_hd__nor2_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18983_ _19007_/B _18983_/B _18981_/X _18982_/Y vssd1 vssd1 vccd1 vccd1 _18983_/X
+ sky130_fd_sc_hd__or4bb_4
XANTENNA__18949__D _19751_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ _13056_/B _13056_/C _13056_/A vssd1 vssd1 vccd1 vccd1 _13059_/B sky130_fd_sc_hd__a21o_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17934_ _17794_/A _17794_/C _17794_/B vssd1 vssd1 vccd1 vccd1 _17935_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__18030__C _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12008_ _12899_/B _12268_/B _12007_/B _12004_/X vssd1 vssd1 vccd1 vccd1 _12009_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__20034__B2 _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17865_ _17865_/A _17865_/B vssd1 vssd1 vccd1 vccd1 _17867_/B sky130_fd_sc_hd__nor2_1
X_19604_ _19604_/A _19604_/B _19729_/B vssd1 vssd1 vccd1 vccd1 _19606_/B sky130_fd_sc_hd__nand3_1
X_16816_ _16816_/A _16816_/B vssd1 vssd1 vccd1 vccd1 _16822_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_108_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17796_ _17673_/A _17673_/C _17673_/B vssd1 vssd1 vccd1 vccd1 _17797_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_152_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19535_ _19535_/A _19535_/B _19692_/C _20416_/B vssd1 vssd1 vccd1 vccd1 _19538_/D
+ sky130_fd_sc_hd__nand4_2
X_13959_ _13960_/A _13960_/B vssd1 vssd1 vccd1 vccd1 _14290_/A sky130_fd_sc_hd__and2b_1
X_16747_ _21830_/Q _17019_/C _16746_/B _16743_/X vssd1 vssd1 vccd1 vccd1 _16753_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_76_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17202__A2 _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16678_ _16676_/A _16676_/Y _16677_/Y _16652_/X vssd1 vssd1 vccd1 vccd1 _16682_/A
+ sky130_fd_sc_hd__a211oi_4
X_19466_ _19467_/A _19467_/B _19467_/C vssd1 vssd1 vccd1 vccd1 _19468_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_29_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18950__A2 _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18417_ _18413_/A _18414_/X _18260_/X _18262_/Y vssd1 vssd1 vccd1 vccd1 _18417_/X
+ sky130_fd_sc_hd__o211a_1
X_15629_ hold263/X _15628_/X fanout4/X vssd1 vssd1 vccd1 vccd1 _21878_/D sky130_fd_sc_hd__mux2_1
X_19397_ _19243_/A _19243_/C _19243_/B vssd1 vssd1 vccd1 vccd1 _19398_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18348_ _18348_/A _18348_/B vssd1 vssd1 vccd1 vccd1 _18357_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20735__C _21261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18279_ _18873_/A _18849_/A _18732_/C _19221_/C vssd1 vssd1 vccd1 vccd1 _18281_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15829__C _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20310_ _20460_/A vssd1 vssd1 vccd1 vccd1 _20312_/D sky130_fd_sc_hd__inv_2
XFILLER_0_142_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21290_ _21290_/A _21290_/B vssd1 vssd1 vccd1 vccd1 _21298_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12534__B _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20241_ _20774_/B _20242_/C _20242_/D _20774_/A vssd1 vssd1 vccd1 vccd1 _20244_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18466__A1 _19092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout103_A _19691_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18466__B2 _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19663__B1 _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20172_ _20026_/B _20841_/B _20173_/C _20173_/D vssd1 vssd1 vccd1 vccd1 _20176_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__17763__D _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20432__A1_N _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20025__A1 _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19966__A1 _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12502__A2 _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20025__B2 _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19966__B2 _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout472_A _15091_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19333__A _19493_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12266__A1 _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14477__A _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15072__S fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12018__A1 _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11613__B _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13531__D _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21626_ _21682_/CLK _21626_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[89] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17300__B _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15507__A2 _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21557_ mstream_o[20] hold64/X _21562_/S vssd1 vssd1 vccd1 vccd1 _22084_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11310_ _11224_/A t1x[21] v2z[21] _11223_/A _11309_/X vssd1 vssd1 vccd1 vccd1 _11310_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_105_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20508_ _20639_/A _20506_/X _20324_/Y _20327_/Y vssd1 vssd1 vccd1 vccd1 _20508_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_22_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12290_ fanout9/X _17173_/B vssd1 vssd1 vccd1 vccd1 _12290_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_132_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21488_ hold197/X sstream_i[65] _21489_/S vssd1 vssd1 vccd1 vccd1 _22015_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_50_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12444__B _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14191__A1 _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11241_ _11122_/A t2y[4] t0y[4] _11123_/A vssd1 vssd1 vccd1 vccd1 _11241_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_31_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14191__B2 _14212_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20439_ _20440_/A _20440_/B _20440_/C vssd1 vssd1 vccd1 vccd1 _20441_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_132_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20264__A1 _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20264__B2 _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11172_ hold265/X _11126_/A fanout47/X hold269/A vssd1 vssd1 vccd1 vccd1 _11172_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18131__B _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13556__A _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15980_ _15981_/B _15981_/A vssd1 vssd1 vccd1 vccd1 _15980_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_98_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14931_ _14771_/A _14771_/B _14769_/B vssd1 vssd1 vccd1 vccd1 _14934_/C sky130_fd_sc_hd__o21ai_2
XANTENNA__18149__A2_N _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14862_ _14862_/A _14862_/B _14862_/C vssd1 vssd1 vccd1 vccd1 _14865_/C sky130_fd_sc_hd__nand3_1
X_17650_ _17650_/A _17650_/B vssd1 vssd1 vccd1 vccd1 _17652_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13813_ _13813_/A _13813_/B vssd1 vssd1 vccd1 vccd1 _13814_/B sky130_fd_sc_hd__xnor2_2
X_16601_ _18166_/A _17666_/A _17443_/D _17434_/B vssd1 vssd1 vccd1 vccd1 _16603_/A
+ sky130_fd_sc_hd__a22oi_2
X_17581_ _17602_/B _17580_/B _17580_/C _17580_/D vssd1 vssd1 vccd1 vccd1 _17581_/Y
+ sky130_fd_sc_hd__a22oi_4
X_14793_ _14793_/A _14793_/B _14793_/C vssd1 vssd1 vccd1 vccd1 _14795_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_86_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16532_ _16532_/A _16532_/B _16532_/C vssd1 vssd1 vccd1 vccd1 _16534_/B sky130_fd_sc_hd__nand3_2
X_19320_ _19320_/A _19320_/B _19320_/C vssd1 vssd1 vccd1 vccd1 _19321_/B sky130_fd_sc_hd__or3_1
X_13744_ _13744_/A _13744_/B vssd1 vssd1 vccd1 vccd1 _13746_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13722__C _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10956_ hold208/A hold226/A vssd1 vssd1 vccd1 vccd1 _10957_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_156_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12619__B _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16463_ _17041_/A _16899_/B _17013_/D _17019_/C vssd1 vssd1 vccd1 vccd1 _16463_/X
+ sky130_fd_sc_hd__and4_1
X_19251_ _19248_/X _19249_/Y _19103_/B _19105_/A vssd1 vssd1 vccd1 vccd1 _19252_/C
+ sky130_fd_sc_hd__o211ai_2
X_13675_ _13676_/A _13676_/B vssd1 vssd1 vccd1 vccd1 _13833_/A sky130_fd_sc_hd__nor2_1
X_10887_ mstream_o[48] _10886_/Y _10992_/S vssd1 vssd1 vccd1 vccd1 _21585_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_155_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15414_ _15415_/B _15415_/A vssd1 vssd1 vccd1 vccd1 _15560_/A sky130_fd_sc_hd__nand2b_1
X_18202_ _18652_/A _18498_/B _19866_/D _19874_/B vssd1 vssd1 vccd1 vccd1 _18204_/B
+ sky130_fd_sc_hd__nand4_2
X_19182_ _19182_/A _19182_/B vssd1 vssd1 vccd1 vccd1 _19184_/A sky130_fd_sc_hd__xnor2_4
X_12626_ _12627_/A _12627_/B vssd1 vssd1 vccd1 vccd1 _12743_/B sky130_fd_sc_hd__nand2_1
X_16394_ _16394_/A _16394_/B vssd1 vssd1 vccd1 vccd1 _16435_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_66_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18133_ _19185_/D _19223_/B vssd1 vssd1 vccd1 vccd1 _18134_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15345_ _15345_/A _15345_/B vssd1 vssd1 vccd1 vccd1 _15347_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_65_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ _12558_/A _12558_/B vssd1 vssd1 vccd1 vccd1 _12653_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_136_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11508_ _11224_/A t2x[19] v1z[19] fanout21/X _11507_/X vssd1 vssd1 vccd1 vccd1 _11508_/X
+ sky130_fd_sc_hd__a221o_1
X_18064_ _18652_/A _18498_/B _19414_/C _19866_/D vssd1 vssd1 vccd1 vccd1 _18066_/B
+ sky130_fd_sc_hd__nand4_2
X_15276_ _15273_/Y _15406_/A _15808_/C _16424_/A vssd1 vssd1 vccd1 vccd1 _15406_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_112_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12488_ _12825_/A _12488_/B vssd1 vssd1 vccd1 vccd1 _12708_/B sky130_fd_sc_hd__nand2_2
Xhold108 hold108/A vssd1 vssd1 vccd1 vccd1 hold108/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17015_ _17141_/A _17013_/C _17013_/D _17141_/B vssd1 vssd1 vccd1 vccd1 _17016_/C
+ sky130_fd_sc_hd__a22o_1
X_14227_ _14226_/B _14226_/C _14226_/A vssd1 vssd1 vccd1 vccd1 _14228_/C sky130_fd_sc_hd__a21o_1
Xhold119 hold119/A vssd1 vssd1 vccd1 vccd1 hold119/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11439_ hold245/A fanout28/X _11438_/X vssd1 vssd1 vccd1 vccd1 _11439_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_0_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16459__B1 _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14158_ _14020_/D _14021_/B _14156_/Y _14157_/X vssd1 vssd1 vccd1 vccd1 _14160_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19648__A1_N _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13109_ _13109_/A _13109_/B vssd1 vssd1 vccd1 vccd1 _13111_/B sky130_fd_sc_hd__xnor2_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14089_ _14089_/A hold313/A hold319/A vssd1 vssd1 vccd1 vccd1 _14090_/C sky130_fd_sc_hd__and3_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18966_ _18802_/A _18802_/B _18802_/C vssd1 vssd1 vccd1 vccd1 _18967_/C sky130_fd_sc_hd__a21bo_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13185__B _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17917_ _21087_/D _18789_/A _18047_/A _17917_/D vssd1 vssd1 vccd1 vccd1 _18047_/B
+ sky130_fd_sc_hd__nand4_2
X_18897_ _19686_/B _19529_/B _19240_/B _19057_/C vssd1 vssd1 vccd1 vccd1 _18897_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17848_ _18127_/B _17848_/B vssd1 vssd1 vccd1 vccd1 _17850_/B sky130_fd_sc_hd__nor2_1
XANTENNA__15434__A1 _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16496__B _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13913__B _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17779_ _17915_/A _18787_/A _18787_/B _17657_/A vssd1 vssd1 vccd1 vccd1 _17780_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13996__A1 _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19518_ _19676_/B _19518_/B vssd1 vssd1 vccd1 vccd1 _19521_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_53_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13996__B2 _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20790_ _20790_/A _20790_/B vssd1 vssd1 vccd1 vccd1 _20830_/A sky130_fd_sc_hd__or2_1
XFILLER_0_14_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19449_ _19449_/A _19449_/B vssd1 vssd1 vccd1 vccd1 _19452_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_14_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18136__B1 _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21411_ hold117/X fanout40/X _21410_/X vssd1 vssd1 vccd1 vccd1 _21945_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout220_A _18789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout318_A _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14463__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21342_ hold125/X _21381_/B _21341_/X vssd1 vssd1 vccd1 vccd1 _21921_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_103_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16162__A2 _14698_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21273_ _21256_/A _21278_/B _21155_/X _21156_/X _21258_/B vssd1 vssd1 vccd1 vccd1
+ _21274_/B sky130_fd_sc_hd__a32o_1
XFILLER_0_102_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14760__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20246__A1 _21832_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20246__B2 _21831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13920__A1 _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20224_ _20224_/A _20224_/B _20224_/C vssd1 vssd1 vccd1 vccd1 _20224_/X sky130_fd_sc_hd__and3_1
XANTENNA__13920__B2 _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15575__B _21787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20155_ _20156_/A _20156_/B vssd1 vssd1 vccd1 vccd1 _20155_/X sky130_fd_sc_hd__and2b_1
XANTENNA__14476__A2 _14477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20086_ hold50/X _20085_/X fanout4/X vssd1 vssd1 vccd1 vccd1 _21907_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_85_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20549__A2 _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15591__A _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17414__A2 _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ _10810_/A _10810_/B vssd1 vssd1 vccd1 vccd1 _11061_/A sky130_fd_sc_hd__nand2_2
XTAP_2858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11790_ _11764_/A _11764_/B _11764_/C vssd1 vssd1 vccd1 vccd1 _11791_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20988_ _20991_/D vssd1 vssd1 vccd1 vccd1 _20988_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_156_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15131__A2_N _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_29_clk_i_A clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13460_ _15217_/A _14212_/C _13461_/C _13461_/D vssd1 vssd1 vccd1 vccd1 _13462_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_48_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12849__A2_N _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12411_ _12307_/A _12307_/B _12305_/X vssd1 vssd1 vccd1 vccd1 _12413_/B sky130_fd_sc_hd__a21bo_1
X_21609_ _21934_/CLK _21609_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[72] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_91_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13391_ _13243_/A _13243_/B _13241_/X vssd1 vssd1 vccd1 vccd1 _13393_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15130_ _16173_/A _16284_/A _16326_/A _16418_/A vssd1 vssd1 vccd1 vccd1 _15271_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_23_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12342_ _12642_/A _12899_/B vssd1 vssd1 vccd1 vccd1 _12346_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17965__B _17966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10973__A1 _10972_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15766__A _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15061_ _14901_/A _14901_/B _14899_/Y vssd1 vssd1 vccd1 vccd1 _15063_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_65_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19238__A _19692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12273_ _12259_/Y _12271_/A _12271_/B _12267_/Y _12267_/C vssd1 vssd1 vccd1 vccd1
+ _12275_/C sky130_fd_sc_hd__o311a_1
X_14012_ _14284_/A _14011_/B _14131_/A _14011_/D vssd1 vssd1 vccd1 vccd1 _14012_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__13911__A1 _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ _11224_/A _11555_/B vssd1 vssd1 vccd1 vccd1 _11224_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__12714__A2 _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13911__B2 _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15916__D _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18820_ _18817_/X _18818_/X _18669_/C _18668_/Y vssd1 vssd1 vccd1 vccd1 _18822_/D
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__12190__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11155_ hold199/X fanout23/X _11154_/X vssd1 vssd1 vccd1 vccd1 _11155_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12621__C _12621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18751_ _19529_/B _19240_/B _18751_/C _18906_/A vssd1 vssd1 vccd1 vccd1 _18906_/B
+ sky130_fd_sc_hd__nand4_2
X_15963_ _14508_/A _21788_/Q _10797_/Y _14813_/A vssd1 vssd1 vccd1 vccd1 _15964_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_11086_ _10978_/Y hold41/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21681_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_41_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13436__D _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17702_ _17703_/A _17703_/B vssd1 vssd1 vccd1 vccd1 _17702_/X sky130_fd_sc_hd__or2_1
X_14914_ _14295_/A _14295_/B _14295_/C _14913_/X vssd1 vssd1 vccd1 vccd1 _14916_/A
+ sky130_fd_sc_hd__a31o_1
X_15894_ _15894_/A _15894_/B vssd1 vssd1 vccd1 vccd1 _16028_/A sky130_fd_sc_hd__nor2_2
X_18682_ _18682_/A _18682_/B vssd1 vssd1 vccd1 vccd1 _18683_/B sky130_fd_sc_hd__nor2_2
X_17633_ _17630_/Y _17631_/X _17535_/X _17538_/Y vssd1 vssd1 vccd1 vccd1 _17633_/X
+ sky130_fd_sc_hd__o211a_1
X_14845_ _14844_/B _14844_/C _14844_/A vssd1 vssd1 vccd1 vccd1 _14846_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14776_ _14774_/D _15838_/B _16374_/B _14621_/D vssd1 vssd1 vccd1 vccd1 _14777_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_86_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17564_ _17564_/A _17564_/B _17564_/C vssd1 vssd1 vccd1 vccd1 _17567_/A sky130_fd_sc_hd__nand3_2
X_11988_ _11914_/A _11914_/C _11914_/B vssd1 vssd1 vccd1 vccd1 _11989_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19303_ _19303_/A _19303_/B vssd1 vssd1 vccd1 vccd1 _19304_/B sky130_fd_sc_hd__xnor2_2
X_13727_ _13883_/A _13727_/B vssd1 vssd1 vccd1 vccd1 _13729_/B sky130_fd_sc_hd__and2_1
X_16515_ _16989_/C _17013_/C _16446_/X _16447_/X _16917_/C vssd1 vssd1 vccd1 vccd1
+ _16674_/A sky130_fd_sc_hd__a32o_1
X_10939_ _10940_/A _10940_/B _10938_/Y vssd1 vssd1 vccd1 vccd1 _10945_/B sky130_fd_sc_hd__o21bai_2
X_17495_ _17614_/B _17495_/B vssd1 vssd1 vccd1 vccd1 _17498_/A sky130_fd_sc_hd__or2_1
XFILLER_0_6_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18317__A _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14927__B1 _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19234_ _19234_/A _19234_/B vssd1 vssd1 vccd1 vccd1 _19248_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13658_ _13504_/X _13508_/A _13656_/Y _13657_/X vssd1 vssd1 vccd1 vccd1 _13813_/A
+ sky130_fd_sc_hd__a211o_2
X_16446_ _17029_/A _16917_/C _16968_/C _17029_/B vssd1 vssd1 vccd1 vccd1 _16446_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20285__C _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12609_ _13682_/C _13258_/C _13258_/D _13822_/B vssd1 vssd1 vccd1 vccd1 _12610_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_144_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16377_ _16377_/A _16377_/B vssd1 vssd1 vccd1 vccd1 _16378_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_121_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19165_ _18999_/A _18835_/Y _18997_/Y vssd1 vssd1 vccd1 vccd1 _19165_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13589_ _21742_/Q _14195_/A _14384_/A _14212_/B vssd1 vssd1 vccd1 vccd1 _13591_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_42_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15328_ _15328_/A _15328_/B _15328_/C vssd1 vssd1 vccd1 vccd1 _15328_/X sky130_fd_sc_hd__and3_1
XFILLER_0_124_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18116_ _18114_/Y _18116_/B vssd1 vssd1 vccd1 vccd1 _18117_/B sky130_fd_sc_hd__and2b_1
XANTENNA__19330__A2 _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19096_ _18936_/A _18936_/B _18936_/C vssd1 vssd1 vccd1 vccd1 _19097_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15259_ _15259_/A _15451_/B vssd1 vssd1 vccd1 vccd1 _15270_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_83_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18047_ _18047_/A _18047_/B vssd1 vssd1 vccd1 vccd1 _18057_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15395__B _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11913__B1 _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout407 _21768_/Q vssd1 vssd1 vccd1 vccd1 _15514_/B sky130_fd_sc_hd__buf_6
XFILLER_0_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout418 _21765_/Q vssd1 vssd1 vccd1 vccd1 _12897_/D sky130_fd_sc_hd__clkbuf_8
XANTENNA__18202__D _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout429 _21763_/Q vssd1 vssd1 vccd1 vccd1 _14716_/A sky130_fd_sc_hd__buf_4
X_19998_ _19997_/A _20138_/B _19997_/C vssd1 vssd1 vccd1 vccd1 _19999_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_10_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18949_ _19439_/A _19951_/A _19753_/B _19751_/C vssd1 vssd1 vccd1 vccd1 _19106_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__13666__B1 _10852_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16938__C _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21960_ _21963_/CLK _21960_/D vssd1 vssd1 vccd1 vccd1 hold278/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_119_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20911_ _20911_/A _20911_/B vssd1 vssd1 vccd1 vccd1 _20912_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_94_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk_i _21806_/CLK vssd1 vssd1 vccd1 vccd1 _21821_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21891_ _21923_/CLK _21891_/D vssd1 vssd1 vccd1 vccd1 hold229/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout170_A _21828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14938__A2_N _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout268_A _17417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13969__A1 _12291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20842_ _20842_/A _20971_/B vssd1 vssd1 vccd1 vccd1 _20844_/A sky130_fd_sc_hd__or2_2
XFILLER_0_77_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20773_ _20658_/A _20912_/A _20651_/B vssd1 vssd1 vccd1 vccd1 _20786_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout14 wire16/X vssd1 vssd1 vccd1 vccd1 _11521_/S sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout435_A _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout25 _11284_/S vssd1 vssd1 vccd1 vccd1 _11260_/S sky130_fd_sc_hd__buf_6
Xfanout36 _21490_/S vssd1 vssd1 vccd1 vccd1 _21528_/S sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_30_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20476__B _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout47 fanout49/X vssd1 vssd1 vccd1 vccd1 fanout47/X sky130_fd_sc_hd__buf_4
XFILLER_0_147_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_29_clk_i clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21932_/CLK sky130_fd_sc_hd__clkbuf_16
Xfanout58 fanout59/X vssd1 vssd1 vccd1 vccd1 fanout58/X sky130_fd_sc_hd__buf_4
XFILLER_0_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout69 _20838_/D vssd1 vssd1 vccd1 vccd1 _21296_/B sky130_fd_sc_hd__buf_4
XFILLER_0_130_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout602_A _11459_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14193__C _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15343__B1 _15151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21325_ _11550_/B _16437_/Y fanout8/X vssd1 vssd1 vccd1 vccd1 _21325_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_5_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14697__A2 _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21416__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21256_ _21256_/A _21256_/B vssd1 vssd1 vccd1 vccd1 _21257_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12722__B _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18897__A _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20207_ _20208_/B _20208_/A vssd1 vssd1 vccd1 vccd1 _20207_/X sky130_fd_sc_hd__and2b_1
XANTENNA__18112__D _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21187_ _21231_/A vssd1 vssd1 vccd1 vccd1 _21187_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11380__A1 _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout83_A _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15807__A1_N _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20138_ _20138_/A _20138_/B vssd1 vssd1 vccd1 vccd1 _20140_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_102_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17306__A _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20069_ _20069_/A _20069_/B vssd1 vssd1 vccd1 vccd1 _20070_/B sky130_fd_sc_hd__xnor2_1
X_12960_ _12600_/A _12956_/X _12957_/Y _12959_/X vssd1 vssd1 vccd1 vccd1 _14294_/D
+ sky130_fd_sc_hd__a31o_4
XTAP_3301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11911_ _12458_/A _12357_/C _12877_/B _12751_/B vssd1 vssd1 vccd1 vccd1 _11914_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_3334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18060__A2 _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ _12891_/A _13010_/B _12891_/C vssd1 vssd1 vccd1 vccd1 _12891_/Y sky130_fd_sc_hd__nand3_2
XTAP_3356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_301 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_312 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14630_ _14630_/A _14630_/B vssd1 vssd1 vccd1 vccd1 _14650_/A sky130_fd_sc_hd__or2_2
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_323 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ _12458_/A _12357_/C _12443_/A _12877_/B vssd1 vssd1 vccd1 vccd1 _11845_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_135_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_334 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14561_ _14560_/B _14724_/B _14560_/A vssd1 vssd1 vccd1 vccd1 _14562_/B sky130_fd_sc_hd__a21o_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18899__A1 _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19240__B _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11773_ _11772_/A _11772_/Y _11752_/X _11754_/Y vssd1 vssd1 vccd1 vccd1 _11776_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_71_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14665__A _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18137__A _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16300_ _16300_/A _16300_/B vssd1 vssd1 vccd1 vccd1 _16301_/B sky130_fd_sc_hd__nor2_1
X_13512_ _13512_/A _13520_/A vssd1 vssd1 vccd1 vccd1 _13518_/D sky130_fd_sc_hd__xnor2_4
XANTENNA__17020__B1 _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17280_ _17490_/A _17282_/A _17739_/C _17739_/D _17186_/B vssd1 vssd1 vccd1 vccd1
+ _17290_/A sky130_fd_sc_hd__a41o_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14492_ _14492_/A _14492_/B vssd1 vssd1 vccd1 vccd1 _14494_/B sky130_fd_sc_hd__xnor2_4
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14384__B _15892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16231_ _16228_/X _16229_/Y _16113_/Y _16115_/Y vssd1 vssd1 vccd1 vccd1 _16232_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_138_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13443_ _13443_/A _13443_/B vssd1 vssd1 vccd1 vccd1 _13444_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12396__B1 _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16162_ _16273_/A _14698_/D _16163_/C _16163_/D vssd1 vssd1 vccd1 vccd1 _16164_/A
+ sky130_fd_sc_hd__a22oi_1
X_13374_ _13240_/A _13239_/B _13237_/Y vssd1 vssd1 vccd1 vccd1 _13390_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_140_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15113_ _15113_/A vssd1 vssd1 vccd1 vccd1 _15115_/D sky130_fd_sc_hd__inv_2
XANTENNA__14137__A1 _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12325_ _12639_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _12329_/A sky130_fd_sc_hd__nand2_1
X_16093_ _16092_/D _21788_/Q _16374_/B _14508_/A vssd1 vssd1 vccd1 vccd1 _16095_/C
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14137__B2 _14463_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21407__A0 _15888_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15044_ _15044_/A _15044_/B _15044_/C vssd1 vssd1 vccd1 vccd1 _15044_/Y sky130_fd_sc_hd__nand3_2
X_19921_ _19712_/Y _19714_/X _19919_/X _19920_/Y vssd1 vssd1 vccd1 vccd1 _19921_/Y
+ sky130_fd_sc_hd__o211ai_4
X_12256_ _12256_/A _12256_/B _12256_/C vssd1 vssd1 vccd1 vccd1 _12258_/B sky130_fd_sc_hd__or3_1
XFILLER_0_107_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11207_ _15370_/B _11206_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21752_/D sky130_fd_sc_hd__mux2_1
X_19852_ _19951_/A _19951_/B _20247_/C _20247_/D vssd1 vssd1 vccd1 vccd1 _19950_/A
+ sky130_fd_sc_hd__nand4_2
X_12187_ _12267_/A _12246_/C _12246_/D _12242_/B vssd1 vssd1 vccd1 vccd1 _12188_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__11371__A1 _17063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15637__A1 _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18803_ _18802_/B _18802_/C _18802_/A vssd1 vssd1 vccd1 vccd1 _18805_/B sky130_fd_sc_hd__a21o_1
X_11138_ _12246_/C _11137_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21729_/D sky130_fd_sc_hd__mux2_1
X_19783_ _19631_/A _19630_/B _19628_/Y vssd1 vssd1 vccd1 vccd1 _19785_/B sky130_fd_sc_hd__a21oi_1
X_16995_ _16994_/A _16994_/Y _16946_/X _16965_/Y vssd1 vssd1 vccd1 vccd1 _17002_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17861__D _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18734_ _19487_/B _19053_/B vssd1 vssd1 vccd1 vccd1 _18735_/B sky130_fd_sc_hd__nand2_1
X_15946_ _15816_/B _15817_/Y _15944_/Y _15945_/X vssd1 vssd1 vccd1 vccd1 _15948_/B
+ sky130_fd_sc_hd__a211oi_4
X_11069_ _10860_/Y hold55/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21664_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_92_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18665_ _18664_/B _18664_/C _18664_/A vssd1 vssd1 vccd1 vccd1 _18665_/Y sky130_fd_sc_hd__a21oi_2
X_15877_ _15874_/X _15875_/Y _15741_/A _15740_/Y vssd1 vssd1 vccd1 vccd1 _15877_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_116_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17616_ _17616_/A _17616_/B vssd1 vssd1 vccd1 vccd1 _17617_/B sky130_fd_sc_hd__xor2_4
XANTENNA__19339__A2_N _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14828_ _16173_/A _14828_/B _16409_/A _16328_/A vssd1 vssd1 vccd1 vccd1 _15029_/A
+ sky130_fd_sc_hd__nand4_2
X_18596_ _19686_/B _19529_/B _19068_/C _19238_/C vssd1 vssd1 vccd1 vccd1 _18598_/D
+ sky130_fd_sc_hd__nand4_1
XTAP_3890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17547_ _17548_/A _17548_/B vssd1 vssd1 vccd1 vccd1 _17652_/A sky130_fd_sc_hd__nand2b_2
X_14759_ _14759_/A _14911_/B vssd1 vssd1 vccd1 vccd1 _19636_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__13820__B1 _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17478_ _17478_/A _17478_/B vssd1 vssd1 vccd1 vccd1 _17593_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_50_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19217_ _19218_/A _19218_/B vssd1 vssd1 vccd1 vccd1 _19327_/B sky130_fd_sc_hd__and2b_1
X_16429_ _16429_/A _16429_/B vssd1 vssd1 vccd1 vccd1 _16430_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11711__B _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19148_ _19148_/A _19148_/B _19148_/C vssd1 vssd1 vccd1 vccd1 _19148_/X sky130_fd_sc_hd__and3_1
XFILLER_0_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14128__A1 _12291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12245__D _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19079_ _19078_/B _19078_/C _19078_/A vssd1 vssd1 vccd1 vccd1 _19079_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_41_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21110_ _21110_/A _21110_/B _21110_/C vssd1 vssd1 vccd1 vccd1 _21110_/X sky130_fd_sc_hd__and3_1
XANTENNA__19067__A1 _19692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20462__D _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22090_ _22105_/CLK _22090_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[26] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_10_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21041_ _21041_/A _21209_/B vssd1 vssd1 vccd1 vccd1 _21052_/A sky130_fd_sc_hd__or2_1
Xfanout204 _21817_/Q vssd1 vssd1 vccd1 vccd1 _21278_/B sky130_fd_sc_hd__buf_4
XFILLER_0_10_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout215 _19868_/B vssd1 vssd1 vccd1 vccd1 _19262_/C sky130_fd_sc_hd__clkbuf_8
XANTENNA__15628__A1 _12291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout226 _20270_/C vssd1 vssd1 vccd1 vccd1 _21286_/A sky130_fd_sc_hd__buf_4
XANTENNA__11362__A1 _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12261__C _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout237 _21809_/Q vssd1 vssd1 vccd1 vccd1 _20991_/C sky130_fd_sc_hd__buf_2
XFILLER_0_22_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout248 _19379_/B vssd1 vssd1 vccd1 vccd1 _19686_/A sky130_fd_sc_hd__buf_4
Xfanout259 _19230_/A vssd1 vssd1 vccd1 vccd1 _19529_/B sky130_fd_sc_hd__buf_4
XANTENNA_fanout385_A _21773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17126__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16030__A _16031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15572__C _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18578__B1 _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21943_ _21945_/CLK _21943_/D vssd1 vssd1 vccd1 vccd1 hold112/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout552_A _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21874_ _21906_/CLK _21874_/D vssd1 vssd1 vccd1 vccd1 hold205/A sky130_fd_sc_hd__dfxtp_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20825_ _20824_/B _20824_/C _20824_/A vssd1 vssd1 vccd1 vccd1 _20825_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_38_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19060__B _19060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12090__A2 _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19995__B _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20756_ _20755_/A _20755_/B _20755_/C _20755_/D vssd1 vssd1 vccd1 vccd1 _20756_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14635__D _14635_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15564__B1 _15381_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20687_ _21169_/A _21278_/B _21256_/B _21056_/A vssd1 vssd1 vccd1 vccd1 _20691_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21101__A2 _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18404__B _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13829__A _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12155__D _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13590__A2 _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17856__A2 _19051_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12733__A _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12110_ _12110_/A _12153_/A vssd1 vssd1 vccd1 vccd1 _12112_/B sky130_fd_sc_hd__nor2_1
X_21308_ _21308_/A _21308_/B vssd1 vssd1 vccd1 vccd1 _21309_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__19058__A1 _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13090_ _13091_/A _13091_/B vssd1 vssd1 vccd1 vccd1 _13092_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_130_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12452__B _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12041_ _12040_/B _12040_/C _12040_/A vssd1 vssd1 vccd1 vccd1 _12043_/B sky130_fd_sc_hd__a21bo_1
Xhold280 hold280/A vssd1 vssd1 vccd1 vccd1 hold280/X sky130_fd_sc_hd__dlygate4sd3_1
X_21239_ _21240_/A _21240_/B vssd1 vssd1 vccd1 vccd1 _21239_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold291 hold291/A vssd1 vssd1 vccd1 vccd1 hold291/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11353__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15800_ _15800_/A _15800_/B vssd1 vssd1 vccd1 vccd1 _15801_/B sky130_fd_sc_hd__nand2_1
X_13992_ _13992_/A _13992_/B _13992_/C vssd1 vssd1 vccd1 vccd1 _14011_/B sky130_fd_sc_hd__and3_1
X_16780_ _16712_/Y _16777_/X _16776_/X _16756_/Y vssd1 vssd1 vccd1 vccd1 _16785_/B
+ sky130_fd_sc_hd__a211o_1
X_15731_ _15728_/X _15729_/Y _15599_/Y _15601_/Y vssd1 vssd1 vccd1 vccd1 _15733_/C
+ sky130_fd_sc_hd__a211oi_2
XTAP_3120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12943_ _12961_/A _12942_/C _12942_/A vssd1 vssd1 vccd1 vccd1 _12945_/B sky130_fd_sc_hd__a21o_1
XTAP_3131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16044__A1 _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16044__B2 _16380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18450_ _18451_/A _18451_/B vssd1 vssd1 vccd1 vccd1 _18606_/B sky130_fd_sc_hd__nand2_1
X_15662_ _15662_/A _15796_/B vssd1 vssd1 vccd1 vccd1 _15665_/A sky130_fd_sc_hd__or2_1
XTAP_3175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_120 v0z[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12874_ _12971_/A _12872_/Y _12744_/B _12744_/Y vssd1 vssd1 vccd1 vccd1 _12934_/B
+ sky130_fd_sc_hd__a211o_1
XTAP_3186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_131 v1z[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17401_ _17402_/A _17402_/B vssd1 vssd1 vccd1 vccd1 _17512_/B sky130_fd_sc_hd__nand2_1
XANTENNA_142 v1z[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14613_ _14531_/A _14531_/B _14530_/A vssd1 vssd1 vccd1 vccd1 _14652_/A sky130_fd_sc_hd__a21o_2
XANTENNA_153 v1z[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11825_ _11823_/A _11823_/Y _11824_/Y _11794_/X vssd1 vssd1 vccd1 vccd1 _11830_/B
+ sky130_fd_sc_hd__a211o_2
X_15593_ _15713_/A _15978_/B _16092_/D _15593_/D vssd1 vssd1 vccd1 vccd1 _15713_/B
+ sky130_fd_sc_hd__and4b_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18381_ _18377_/X _18379_/Y _18230_/B _18230_/Y vssd1 vssd1 vccd1 vccd1 _18381_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA_164 v2z[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_175 v2z[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_186 hold239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14310__A1_N _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14544_ _14391_/D _14393_/B _14542_/Y _14543_/X vssd1 vssd1 vccd1 vccd1 _14690_/A
+ sky130_fd_sc_hd__a211o_2
XANTENNA_197 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17332_ _18166_/A _18058_/A vssd1 vssd1 vccd1 vccd1 _17336_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19533__A2 _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11756_ _12268_/A _12444_/B vssd1 vssd1 vccd1 vccd1 _11758_/B sky130_fd_sc_hd__and2_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20547__D _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17544__A1 _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17544__B2 _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14475_ _15153_/B _15788_/B _14347_/X _14348_/X _13858_/C vssd1 vssd1 vccd1 vccd1
+ _14480_/A sky130_fd_sc_hd__a32o_1
X_17263_ _17363_/B _17261_/X _16684_/Y _16686_/X vssd1 vssd1 vccd1 vccd1 _17264_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_43_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11687_ _13012_/B _12511_/A vssd1 vssd1 vccd1 vccd1 _11691_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19002_ _20770_/B _21373_/B vssd1 vssd1 vccd1 vccd1 _19002_/Y sky130_fd_sc_hd__nor2_1
X_16214_ _16326_/A _16396_/B _16418_/B _16328_/A vssd1 vssd1 vccd1 vccd1 _16218_/C
+ sky130_fd_sc_hd__a22o_1
X_13426_ _13427_/A _13427_/B _13427_/C vssd1 vssd1 vccd1 vccd1 _13428_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_24_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17194_ _17194_/A _17194_/B vssd1 vssd1 vccd1 vccd1 _17196_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18314__B _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16145_ fanout9/A _21412_/B vssd1 vssd1 vccd1 vccd1 _16145_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_12_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13357_ _13357_/A _13509_/A _13357_/C vssd1 vssd1 vccd1 vccd1 _13509_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_12_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1215 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18033__C _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12308_ _11667_/A _11665_/A _11666_/A vssd1 vssd1 vccd1 vccd1 _12310_/B sky130_fd_sc_hd__o21ai_2
X_16076_ _16078_/A _16078_/B _16078_/C vssd1 vssd1 vccd1 vccd1 _16079_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__13458__B _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13288_ _13875_/B _14384_/A _14212_/B _13877_/A vssd1 vssd1 vccd1 vccd1 _13290_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15027_ _15025_/X _15027_/B vssd1 vssd1 vccd1 vccd1 _15028_/B sky130_fd_sc_hd__nand2b_1
X_19904_ _20103_/A _19906_/D _19745_/X _19746_/X _19866_/C vssd1 vssd1 vccd1 vccd1
+ _19909_/A sky130_fd_sc_hd__a32o_1
X_12239_ _12235_/X _12238_/X _12207_/X _12210_/Y vssd1 vssd1 vccd1 vccd1 _12239_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11344__A1 _11343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17872__C _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15592__A2_N _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19835_ _19671_/X _19673_/Y _19833_/X _19834_/Y vssd1 vssd1 vccd1 vccd1 _19837_/A
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15673__B _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19766_ _19613_/A _19613_/B _19611_/Y vssd1 vssd1 vccd1 vccd1 _19768_/B sky130_fd_sc_hd__a21oi_2
X_16978_ _16978_/A _16983_/B vssd1 vssd1 vccd1 vccd1 _16980_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_78_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18717_ _18718_/A _18718_/B vssd1 vssd1 vccd1 vccd1 _18717_/Y sky130_fd_sc_hd__nand2_1
X_15929_ _15931_/B _16369_/B _16177_/B _15931_/A vssd1 vssd1 vccd1 vccd1 _15933_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19697_ _19693_/X _19695_/Y _19534_/X _19537_/X vssd1 vssd1 vccd1 vccd1 _19698_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18648_ _19874_/B _18647_/X _18646_/X vssd1 vssd1 vccd1 vccd1 _18649_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_94_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13921__B _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18579_ _19487_/A _19487_/B _18732_/C _18894_/B vssd1 vssd1 vccd1 vccd1 _18581_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_52_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20610_ _20611_/B _20611_/A vssd1 vssd1 vccd1 vccd1 _20610_/Y sky130_fd_sc_hd__nand2b_1
X_21590_ _21888_/CLK _21590_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[53] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_35_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14349__A1 _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11280__A0 _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20541_ _21286_/A _21151_/A _21301_/A _21296_/A vssd1 vssd1 vccd1 vccd1 _20544_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout133_A _19087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20472_ _20472_/A _20472_/B vssd1 vssd1 vccd1 vccd1 _20483_/A sky130_fd_sc_hd__or2_1
XFILLER_0_132_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout300_A _21795_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16510__A2 _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22073_ _22080_/CLK _22073_/D fanout639/X vssd1 vssd1 vccd1 vccd1 mstream_o[9] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_61_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11335__A1 _21407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21024_ _21135_/B _21022_/X _20892_/A _20894_/X vssd1 vssd1 vccd1 vccd1 _21025_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_22_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15077__A2 _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11099__A0 _11063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18894__B _18894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11616__B _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11638__A2 _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21926_ _21926_/CLK _21926_/D vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfxtp_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout46_A fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21857_ _21923_/CLK hold75/X vssd1 vssd1 vccd1 vccd1 hold74/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11610_ _11610_/A _11610_/B _11610_/C vssd1 vssd1 vccd1 vccd1 _11610_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20808_ _20808_/A _20808_/B vssd1 vssd1 vccd1 vccd1 _20819_/A sky130_fd_sc_hd__or2_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ _12587_/X _12588_/X _12479_/C _12479_/Y vssd1 vssd1 vccd1 vccd1 _12590_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21788_ _21788_/CLK _21788_/D vssd1 vssd1 vccd1 vccd1 _21788_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_108_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14365__D _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11271__B1 _11270_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11541_ _11544_/A1 t2x[30] v1z[30] fanout21/X _11540_/X vssd1 vssd1 vccd1 vccd1 _11541_/X
+ sky130_fd_sc_hd__a221o_1
X_20739_ _20740_/A _20740_/B vssd1 vssd1 vccd1 vccd1 _20739_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_19_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14260_ _14260_/A _14260_/B _14260_/C vssd1 vssd1 vccd1 vccd1 _14260_/X sky130_fd_sc_hd__and3_1
XFILLER_0_52_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13380__A2_N _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11472_ _11502_/A1 t2x[7] v1z[7] fanout18/X _11471_/X vssd1 vssd1 vccd1 vccd1 _11472_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14662__B _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13211_ _13072_/B _13071_/Y _13209_/X _13210_/Y vssd1 vssd1 vccd1 vccd1 _13213_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__13559__A _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14191_ _14212_/B _14365_/D _14054_/X _14055_/X _14212_/C vssd1 vssd1 vccd1 vccd1
+ _14196_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_116_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13142_ _13142_/A _13142_/B _13142_/C vssd1 vssd1 vccd1 vccd1 _13142_/X sky130_fd_sc_hd__and3_2
XFILLER_0_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15774__A _16031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13073_ _13072_/B _13072_/C _13072_/A vssd1 vssd1 vccd1 vccd1 _13073_/Y sky130_fd_sc_hd__o21ai_2
X_17950_ _17810_/B _17809_/Y _17948_/X _17949_/Y vssd1 vssd1 vccd1 vccd1 _17953_/B
+ sky130_fd_sc_hd__o211a_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21389__A2 _21390_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16901_ _16901_/A _16952_/A vssd1 vssd1 vccd1 vccd1 _16903_/B sky130_fd_sc_hd__xor2_1
X_12024_ _11941_/X _12012_/Y _12011_/Y _12011_/A vssd1 vssd1 vccd1 vccd1 _12025_/B
+ sky130_fd_sc_hd__o211ai_1
X_17881_ _17881_/A _17881_/B _17881_/C vssd1 vssd1 vccd1 vccd1 _17883_/B sky130_fd_sc_hd__nand3_2
XANTENNA__18254__A2 _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11877__A2 _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16265__A1 _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12910__B _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16265__B2 _16391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13294__A _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19620_ _19620_/A _19620_/B vssd1 vssd1 vccd1 vccd1 _19621_/B sky130_fd_sc_hd__xor2_2
X_16832_ _16833_/A _16832_/B _17206_/B _17146_/D vssd1 vssd1 vccd1 vccd1 _16898_/A
+ sky130_fd_sc_hd__and4b_1
Xfanout590 _11224_/A vssd1 vssd1 vccd1 vccd1 _11544_/A1 sky130_fd_sc_hd__buf_4
X_19551_ _19551_/A _19551_/B _19551_/C vssd1 vssd1 vccd1 vccd1 _19554_/A sky130_fd_sc_hd__nand3_1
X_16763_ _17206_/B _17277_/A _16762_/B _16759_/X vssd1 vssd1 vccd1 vccd1 _16765_/B
+ sky130_fd_sc_hd__a31o_1
X_13975_ _14138_/A _13975_/B _16328_/B _16399_/B vssd1 vssd1 vccd1 vccd1 _14142_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_88_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18502_ _18352_/A _18352_/C _18352_/B vssd1 vssd1 vccd1 vccd1 _18503_/C sky130_fd_sc_hd__a21bo_1
X_15714_ _15714_/A _15714_/B vssd1 vssd1 vccd1 vccd1 _15722_/A sky130_fd_sc_hd__nand2_1
X_12926_ _12798_/B _12798_/Y _12923_/X _12925_/Y vssd1 vssd1 vccd1 vccd1 _12929_/B
+ sky130_fd_sc_hd__a211oi_4
X_19482_ _19343_/A _19343_/B _19346_/A vssd1 vssd1 vccd1 vccd1 _19631_/A sky130_fd_sc_hd__a21o_1
X_16694_ _16694_/A _16694_/B _16694_/C vssd1 vssd1 vccd1 vccd1 _16698_/A sky130_fd_sc_hd__nand3_1
XANTENNA__18962__B1 _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18433_ _19487_/A _19382_/B _18431_/Y _18588_/A vssd1 vssd1 vccd1 vccd1 _18435_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_15645_ _15645_/A _15645_/B vssd1 vssd1 vccd1 vccd1 _15647_/B sky130_fd_sc_hd__xnor2_1
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ _13858_/B _15768_/A _12752_/X _12751_/X _13152_/C vssd1 vssd1 vccd1 vccd1
+ _12862_/A sky130_fd_sc_hd__a32o_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19506__A2 _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18364_ _18363_/B _18363_/C _18363_/A vssd1 vssd1 vccd1 vccd1 _18364_/Y sky130_fd_sc_hd__a21oi_2
X_11808_ _12268_/A _12877_/B vssd1 vssd1 vccd1 vccd1 _11810_/B sky130_fd_sc_hd__and2_1
XFILLER_0_139_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15576_ _15576_/A _15700_/B vssd1 vssd1 vccd1 vccd1 _15578_/A sky130_fd_sc_hd__or2_2
X_12788_ _12787_/B _12787_/C _12787_/A vssd1 vssd1 vccd1 vccd1 _12790_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12054__A2 _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12357__B _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17315_ _17315_/A _17315_/B vssd1 vssd1 vccd1 vccd1 _17317_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14527_ _14526_/B _14526_/C _14526_/A vssd1 vssd1 vccd1 vccd1 _14527_/Y sky130_fd_sc_hd__a21oi_1
X_11739_ _12784_/A _13017_/A vssd1 vssd1 vccd1 vccd1 _11741_/B sky130_fd_sc_hd__and2_1
XFILLER_0_56_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18295_ _19373_/B _19051_/A _19068_/C _19238_/C vssd1 vssd1 vccd1 vccd1 _18442_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17246_ _17245_/B _17245_/C _17245_/A vssd1 vssd1 vccd1 vccd1 _17248_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_142_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14458_ _16084_/C _14457_/X _14456_/X vssd1 vssd1 vccd1 vccd1 _14460_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_25_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13409_ _13409_/A _13409_/B vssd1 vssd1 vccd1 vccd1 _13410_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_40_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14389_ _15373_/A _15373_/B _16418_/A _16268_/B vssd1 vssd1 vccd1 vccd1 _14391_/D
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17177_ _16553_/A _16553_/B _16551_/Y vssd1 vssd1 vccd1 vccd1 _17265_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_113_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11565__A1 _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16128_ _16128_/A _16128_/B _16128_/C vssd1 vssd1 vccd1 vccd1 _16128_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_110_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19690__B2 _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14503__A1 _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18698__C _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16059_ _16173_/A _16284_/A _16177_/B _16286_/B vssd1 vssd1 vccd1 vccd1 _16171_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__14503__B2 _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11317__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11317__B2 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16499__B _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19818_ _19818_/A _19818_/B vssd1 vssd1 vccd1 vccd1 _19840_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19749_ _19749_/A _19749_/B vssd1 vssd1 vccd1 vccd1 _19756_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_155_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19745__A2 _19868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16559__A2 _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21711_ _22105_/CLK _21711_/D vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_63_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17123__B _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout250_A _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout348_A hold241/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21642_ _21722_/CLK _21642_/D fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[105]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__12045__A2 _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21304__A2 _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12267__B _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_20 _11339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21573_ mstream_o[36] _11053_/X _21579_/S vssd1 vssd1 vccd1 vccd1 _22100_/D sky130_fd_sc_hd__mux2_1
XANTENNA_31 _11343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout515_A _13018_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_42 _11445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_53 hold275/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20524_ _20528_/A _20686_/B vssd1 vssd1 vccd1 vccd1 _20529_/A sky130_fd_sc_hd__or2_1
XFILLER_0_145_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_64 hold274/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_75 hold277/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_86 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_97 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13379__A _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20455_ _20845_/D _20721_/D _21286_/B _21296_/B vssd1 vssd1 vccd1 vccd1 _20588_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__20047__A1_N _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21624__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_1265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20386_ _20386_/A _20386_/B vssd1 vssd1 vccd1 vccd1 _20913_/A sky130_fd_sc_hd__or2_4
XFILLER_0_28_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11308__A1 _11307_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22056_ _22063_/CLK _22056_/D vssd1 vssd1 vccd1 vccd1 hold299/A sky130_fd_sc_hd__dfxtp_4
X_21007_ _20826_/Y _20830_/B _21005_/X _21006_/Y vssd1 vssd1 vccd1 vccd1 _21008_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__17444__B1 _17443_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13760_ _13757_/X _13758_/Y _13599_/Y _13601_/X vssd1 vssd1 vccd1 vccd1 _13795_/B
+ sky130_fd_sc_hd__o211a_1
X_10972_ _10972_/A _10972_/B vssd1 vssd1 vccd1 vccd1 _10972_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_69_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21909_ _21942_/CLK _21909_/D vssd1 vssd1 vccd1 vccd1 hold101/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12711_ fanout9/X _21343_/B vssd1 vssd1 vccd1 vccd1 _12711_/Y sky130_fd_sc_hd__nor2_1
X_13691_ _13534_/A _13535_/Y _13689_/A _13690_/X vssd1 vssd1 vccd1 vccd1 _13691_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_97_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15430_ _15334_/B _15430_/B vssd1 vssd1 vccd1 vccd1 _15473_/A sky130_fd_sc_hd__nand2b_2
X_12642_ _12642_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _12646_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11244__A0 _12242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15361_ _15361_/A _15361_/B vssd1 vssd1 vccd1 vccd1 _15362_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12573_ _12572_/B _12572_/C _12572_/A vssd1 vssd1 vccd1 vccd1 _12575_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_93_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20394__B _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17100_ _17099_/B _17099_/C _17099_/A vssd1 vssd1 vccd1 vccd1 _17101_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_110_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14312_ _14133_/D _16406_/B _16314_/D _14312_/D vssd1 vssd1 vccd1 vccd1 _14315_/A
+ sky130_fd_sc_hd__and4b_2
X_11524_ _11523_/X _19199_/C _11545_/S vssd1 vssd1 vccd1 vccd1 _21846_/D sky130_fd_sc_hd__mux2_1
X_15292_ _15292_/A _15292_/B vssd1 vssd1 vccd1 vccd1 _15292_/X sky130_fd_sc_hd__or2_1
XFILLER_0_124_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18080_ _18076_/X _18078_/Y _17943_/B _17943_/Y vssd1 vssd1 vccd1 vccd1 _18082_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_135_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12905__B _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14243_ _14557_/D _14242_/X _14241_/X vssd1 vssd1 vccd1 vccd1 _14245_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__13289__A _13875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17031_ _17096_/A _17145_/B _17021_/B _17019_/X vssd1 vssd1 vccd1 vccd1 _17035_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_150_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11455_ _11454_/X _17557_/B _11470_/S vssd1 vssd1 vccd1 vccd1 _21823_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_40_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14174_ _14045_/B _14174_/B vssd1 vssd1 vccd1 vccd1 _14208_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_22_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11386_ _11385_/X _17223_/A _11401_/S vssd1 vssd1 vccd1 vccd1 _21800_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_150_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16486__A1 _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13125_ _13124_/A _13124_/B _13124_/C vssd1 vssd1 vccd1 vccd1 _13126_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__16486__B2 _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12343__D _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18982_ _18979_/Y _18980_/X _18815_/X _18817_/X vssd1 vssd1 vccd1 vccd1 _18982_/Y
+ sky130_fd_sc_hd__o211ai_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ _13056_/A _13056_/B _13056_/C vssd1 vssd1 vccd1 vccd1 _13059_/A sky130_fd_sc_hd__nand3_2
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17933_ _17932_/B _17932_/C _17932_/A vssd1 vssd1 vccd1 vccd1 _17935_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_84_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17435__B1 _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12007_ _12004_/X _12007_/B vssd1 vssd1 vccd1 vccd1 _12055_/B sky130_fd_sc_hd__and2b_1
XANTENNA__18030__D _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17864_ _17864_/A _17864_/B vssd1 vssd1 vccd1 vccd1 _17867_/A sky130_fd_sc_hd__xnor2_2
X_19603_ _20088_/A _19872_/C _19603_/C _19729_/A vssd1 vssd1 vccd1 vccd1 _19729_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_75_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16815_ _16989_/C _17123_/C _16815_/C _16815_/D vssd1 vssd1 vccd1 vccd1 _16816_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_89_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17795_ _17794_/B _17794_/C _17794_/A vssd1 vssd1 vccd1 vccd1 _17797_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_75_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14848__A _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17224__A _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19534_ _19535_/A _19695_/A _20416_/A _19691_/D vssd1 vssd1 vccd1 vccd1 _19534_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_152_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13272__A2_N _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16746_ _16743_/X _16746_/B vssd1 vssd1 vccd1 vccd1 _16818_/B sky130_fd_sc_hd__and2b_1
X_13958_ _13958_/A _13958_/B vssd1 vssd1 vccd1 vccd1 _13960_/B sky130_fd_sc_hd__nor2_2
XANTENNA__17738__A1 _18010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17738__B2 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12909_ _12909_/A _12909_/B vssd1 vssd1 vccd1 vccd1 _12918_/A sky130_fd_sc_hd__xor2_2
X_19465_ _19465_/A _19465_/B vssd1 vssd1 vccd1 vccd1 _19467_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16677_ _16653_/A _16653_/B _16653_/C vssd1 vssd1 vccd1 vccd1 _16677_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_29_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13889_ _13730_/Y _13733_/X _13886_/Y _13887_/X vssd1 vssd1 vccd1 vccd1 _13889_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_119_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18416_ _18260_/X _18262_/Y _18413_/A _18414_/X vssd1 vssd1 vccd1 vccd1 _18416_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15628_ _12291_/B _15626_/Y _15627_/X vssd1 vssd1 vccd1 vccd1 _15628_/X sky130_fd_sc_hd__a21o_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19396_ _19395_/B _19395_/C _19395_/A vssd1 vssd1 vccd1 vccd1 _19398_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_146_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11235__B1 _11234_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18347_ _18345_/X _18347_/B vssd1 vssd1 vccd1 vccd1 _18348_/B sky130_fd_sc_hd__and2b_1
X_15559_ _15560_/A _15560_/B _15560_/C vssd1 vssd1 vccd1 vccd1 _15561_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_514 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1066 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15398__B _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18278_ _18873_/A _18732_/C _19221_/C _18849_/A vssd1 vssd1 vccd1 vccd1 _18281_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15829__D _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17894__A _18030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17229_ _17229_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17231_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11538__B2 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12534__C _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20240_ _20386_/A _20240_/B vssd1 vssd1 vccd1 vccd1 _20256_/A sky130_fd_sc_hd__or2_1
XANTENNA__18466__A2 _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19663__A1 _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19663__B2 _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13927__A _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20171_ _20314_/A vssd1 vssd1 vccd1 vccd1 _20173_/D sky130_fd_sc_hd__inv_2
XFILLER_0_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12550__B _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout298_A _17063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20025__A2 _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19966__A2 _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19333__B _20841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout465_A _21753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12266__A2 _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14477__B _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_308 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout632_A _21776_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16401__A1 _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16401__B2 _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12018__A2 _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21289__A1 _21293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21625_ _21682_/CLK _21625_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[88] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21556_ mstream_o[19] hold144/X _21562_/S vssd1 vssd1 vccd1 vccd1 _22083_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_62_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_262 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17300__C _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12725__B _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14715__A1 _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20507_ _20324_/Y _20327_/Y _20639_/A _20506_/X vssd1 vssd1 vccd1 vccd1 _20639_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_105_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21487_ hold200/X sstream_i[64] _21489_/S vssd1 vssd1 vccd1 vccd1 _22014_/D sky130_fd_sc_hd__mux2_1
XANTENNA__11529__B2 fanout21/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12444__C _12771_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11240_ _12267_/A _11239_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21761_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14191__A2 _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20438_ _20438_/A _20438_/B vssd1 vssd1 vccd1 vccd1 _20440_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17665__B1 _17924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20264__A2 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13837__A _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11171_ _13157_/A _11170_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21740_/D sky130_fd_sc_hd__mux2_1
X_20369_ _20370_/A _20370_/B vssd1 vssd1 vccd1 vccd1 _20513_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_30_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19227__C _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18131__C _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13556__B _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_25_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13151__B1 _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22039_ _22049_/CLK _22039_/D vssd1 vssd1 vccd1 vccd1 hold228/A sky130_fd_sc_hd__dfxtp_1
X_14930_ _15159_/D _15698_/B _14930_/C _14930_/D vssd1 vssd1 vccd1 vccd1 _14934_/B
+ sky130_fd_sc_hd__nand4_2
X_14861_ _14860_/B _14976_/B _14860_/A vssd1 vssd1 vccd1 vccd1 _14862_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_98_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16600_ _18058_/A _17433_/A vssd1 vssd1 vccd1 vccd1 _16604_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_138_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13812_ _13962_/A _13812_/B vssd1 vssd1 vccd1 vccd1 _13813_/B sky130_fd_sc_hd__nand2_2
X_17580_ _17602_/B _17580_/B _17580_/C _17580_/D vssd1 vssd1 vccd1 vccd1 _17580_/Y
+ sky130_fd_sc_hd__nand4_1
X_14792_ _14791_/B _14946_/B _14791_/A vssd1 vssd1 vccd1 vccd1 _14793_/C sky130_fd_sc_hd__a21o_1
X_16531_ _16531_/A _16531_/B vssd1 vssd1 vccd1 vccd1 _16532_/C sky130_fd_sc_hd__xnor2_1
X_13743_ _13743_/A vssd1 vssd1 vccd1 vccd1 _13744_/B sky130_fd_sc_hd__inv_2
X_10955_ hold208/A hold226/A vssd1 vssd1 vccd1 vccd1 _10957_/A sky130_fd_sc_hd__and2_1
XFILLER_0_98_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13722__D _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16883__A _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19250_ _19103_/B _19105_/A _19248_/X _19249_/Y vssd1 vssd1 vccd1 vccd1 _19252_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12619__C _13269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16462_ _16462_/A _16462_/B vssd1 vssd1 vccd1 vccd1 _16468_/A sky130_fd_sc_hd__xor2_1
X_13674_ _13674_/A _13674_/B vssd1 vssd1 vccd1 vccd1 _13676_/B sky130_fd_sc_hd__xnor2_1
X_10886_ _10886_/A _10886_/B vssd1 vssd1 vccd1 vccd1 _10886_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_38_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18201_ _19445_/A _19414_/C vssd1 vssd1 vccd1 vccd1 _18204_/A sky130_fd_sc_hd__and2_1
XFILLER_0_66_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15413_ _15413_/A _15547_/B vssd1 vssd1 vccd1 vccd1 _15415_/B sky130_fd_sc_hd__or2_1
XFILLER_0_156_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19181_ _19337_/D _19181_/B vssd1 vssd1 vccd1 vccd1 _19182_/B sky130_fd_sc_hd__nand2_2
X_12625_ _12743_/A _12625_/B vssd1 vssd1 vccd1 vccd1 _12627_/B sky130_fd_sc_hd__and2_1
X_16393_ _16393_/A _16393_/B vssd1 vssd1 vccd1 vccd1 _16394_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18132_ _18732_/C _18131_/X _18130_/X vssd1 vssd1 vccd1 vccd1 _18134_/A sky130_fd_sc_hd__a21bo_1
X_15344_ _15345_/B _15345_/A vssd1 vssd1 vccd1 vccd1 _15344_/X sky130_fd_sc_hd__and2b_1
X_12556_ _12556_/A _12556_/B vssd1 vssd1 vccd1 vccd1 _12558_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_109_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16107__B _21784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11507_ _11507_/A1 t1y[19] t0x[19] _11507_/B2 vssd1 vssd1 vccd1 vccd1 _11507_/X sky130_fd_sc_hd__a22o_1
X_18063_ _19445_/A _19262_/C vssd1 vssd1 vccd1 vccd1 _18066_/A sky130_fd_sc_hd__and2_1
XFILLER_0_41_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15275_ _15933_/C _16424_/A _15273_/Y _15406_/A vssd1 vssd1 vccd1 vccd1 _15277_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_123_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12487_ _12484_/X _12485_/Y _12381_/Y _12383_/Y vssd1 vssd1 vccd1 vccd1 _12488_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_79_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold109 hold109/A vssd1 vssd1 vccd1 vccd1 hold109/X sky130_fd_sc_hd__dlygate4sd3_1
X_17014_ _17145_/A _17019_/C vssd1 vssd1 vccd1 vccd1 _17016_/B sky130_fd_sc_hd__and2_1
X_14226_ _14226_/A _14226_/B _14226_/C vssd1 vssd1 vccd1 vccd1 _14228_/B sky130_fd_sc_hd__nand3_2
X_11438_ _11447_/A1 hold214/A fanout48/X hold181/A vssd1 vssd1 vccd1 vccd1 _11438_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14157_ _14306_/A _16328_/B _14157_/C _14157_/D vssd1 vssd1 vccd1 vccd1 _14157_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_42_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11369_ _11124_/A hold255/X fanout45/X hold139/X vssd1 vssd1 vccd1 vccd1 _11369_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ _13244_/A _13250_/B vssd1 vssd1 vccd1 vccd1 _13109_/B sky130_fd_sc_hd__nor2_1
X_14088_ _14089_/A hold313/A hold319/A vssd1 vssd1 vccd1 vccd1 _14090_/B sky130_fd_sc_hd__a21oi_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18965_ _18964_/B _18964_/C _18964_/A vssd1 vssd1 vccd1 vccd1 _18967_/B sky130_fd_sc_hd__o21ai_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ _13169_/B _13038_/C _13038_/A vssd1 vssd1 vccd1 vccd1 _13040_/C sky130_fd_sc_hd__a21o_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17916_ _17915_/A _18787_/B _17915_/D _18787_/A vssd1 vssd1 vccd1 vccd1 _17917_/D
+ sky130_fd_sc_hd__a22o_1
X_18896_ _19686_/B _19240_/B _19057_/C _19230_/A vssd1 vssd1 vccd1 vccd1 _18901_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17847_ _17847_/A _17847_/B _17847_/C vssd1 vssd1 vccd1 vccd1 _17848_/B sky130_fd_sc_hd__and3_1
XFILLER_0_117_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15434__A2 _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13913__C _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17778_ _17915_/A _21087_/D _18787_/A _18787_/B vssd1 vssd1 vccd1 vccd1 _17913_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_117_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18908__B1 _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19187__A1_N _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19517_ _19676_/A _19515_/Y _19356_/B _19358_/B vssd1 vssd1 vccd1 vccd1 _19518_/B
+ sky130_fd_sc_hd__o211ai_1
X_16729_ _16691_/A _16691_/C _16691_/B vssd1 vssd1 vccd1 vccd1 _16730_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13996__A2 _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19448_ _19448_/A _19448_/B vssd1 vssd1 vccd1 vccd1 _19449_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_53_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19379_ _19535_/B _19379_/B _20416_/A _20416_/B vssd1 vssd1 vccd1 vccd1 _19382_/D
+ sky130_fd_sc_hd__nand4_1
XANTENNA__18136__A1 _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18136__B2 _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21410_ _21412_/A _20906_/Y _21421_/S _21409_/Y vssd1 vssd1 vccd1 vccd1 _21410_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11730__A _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14463__D _14463_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17895__B1 _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21341_ _21349_/A _17484_/X _21421_/S _21340_/Y vssd1 vssd1 vccd1 vccd1 _21341_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout213_A _21283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21272_ _21241_/B _21243_/B _21239_/Y vssd1 vssd1 vccd1 vccd1 _21274_/A sky130_fd_sc_hd__a21o_1
XANTENNA__14760__B _19636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20223_ _20221_/X _20223_/B vssd1 vssd1 vccd1 vccd1 _20224_/C sky130_fd_sc_hd__nand2b_1
XANTENNA__20246__A2 _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13920__A2 _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17129__A _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_274 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20154_ _20154_/A _20154_/B vssd1 vssd1 vccd1 vccd1 _20156_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout582_A _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20085_ hold38/X fanout8/X _20084_/X vssd1 vssd1 vccd1 vccd1 _20085_/X sky130_fd_sc_hd__a21bo_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold258_A hold258/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20987_ _21286_/A _21283_/B _21305_/B _21296_/A vssd1 vssd1 vccd1 vccd1 _20991_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12410_ _12410_/A _12410_/B vssd1 vssd1 vccd1 vccd1 _12413_/A sky130_fd_sc_hd__xnor2_1
X_21608_ _21934_/CLK _21608_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[71] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13390_ _13390_/A _13390_/B vssd1 vssd1 vccd1 vccd1 _13393_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_152_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12341_ _11723_/A _11722_/A _11722_/B vssd1 vssd1 vccd1 vccd1 _12348_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_145_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21539_ mstream_o[2] hold85/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22066_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_50_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15060_ _15060_/A _15060_/B vssd1 vssd1 vccd1 vccd1 _15063_/A sky130_fd_sc_hd__xnor2_1
X_12272_ _12267_/Y _12271_/Y _12259_/Y vssd1 vssd1 vccd1 vccd1 _12275_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__15766__B _15892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19238__B _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14011_ _14284_/A _14011_/B _14131_/A _14011_/D vssd1 vssd1 vccd1 vccd1 _14131_/B
+ sky130_fd_sc_hd__nor4_2
X_11223_ _11223_/A _21723_/D vssd1 vssd1 vccd1 vccd1 _11555_/B sky130_fd_sc_hd__or2_4
XANTENNA__17638__B1 _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13911__A2 _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11154_ hold314/X _11126_/A fanout45/X hold308/A vssd1 vssd1 vccd1 vccd1 _11154_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12190__B _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15782__A _15907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18750_ _19529_/B _20148_/C _18751_/C _18906_/A vssd1 vssd1 vccd1 vccd1 _18752_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18796__C _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12621__D _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15962_ _15964_/A vssd1 vssd1 vccd1 vccd1 _16100_/A sky130_fd_sc_hd__inv_2
X_11085_ _10972_/Y hold44/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21680_/D sky130_fd_sc_hd__mux2_1
XANTENNA__21198__B1 _21853_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17701_ _17584_/A _17584_/C _17584_/B vssd1 vssd1 vccd1 vccd1 _17703_/B sky130_fd_sc_hd__a21boi_4
X_14913_ _14913_/A _14913_/B _14913_/C _14445_/A vssd1 vssd1 vccd1 vccd1 _14913_/X
+ sky130_fd_sc_hd__or4b_1
X_18681_ _18678_/X _18679_/X _18525_/C _18525_/Y vssd1 vssd1 vccd1 vccd1 _18682_/B
+ sky130_fd_sc_hd__a211oi_1
X_15893_ _15892_/A _15632_/B _16027_/B vssd1 vssd1 vccd1 vccd1 _15894_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__14398__A _14398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17632_ _17535_/X _17538_/Y _17630_/Y _17631_/X vssd1 vssd1 vccd1 vccd1 _17718_/A
+ sky130_fd_sc_hd__a211oi_4
X_14844_ _14844_/A _14844_/B _14844_/C vssd1 vssd1 vccd1 vccd1 _14846_/A sky130_fd_sc_hd__and3_1
X_17563_ _17562_/A _17562_/B _17562_/C vssd1 vssd1 vccd1 vccd1 _17564_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_59_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14775_ _14777_/A vssd1 vssd1 vccd1 vccd1 _14944_/A sky130_fd_sc_hd__inv_2
X_11987_ _11986_/B _11986_/C _11986_/A vssd1 vssd1 vccd1 vccd1 _11989_/B sky130_fd_sc_hd__a21bo_1
X_19302_ _19303_/A _19303_/B vssd1 vssd1 vccd1 vccd1 _19302_/X sky130_fd_sc_hd__and2b_1
X_16514_ _16507_/X _16668_/A _16564_/B _16513_/X vssd1 vssd1 vccd1 vccd1 _16514_/X
+ sky130_fd_sc_hd__o211a_1
X_13726_ _13723_/Y _13724_/X _13591_/D _13592_/B vssd1 vssd1 vccd1 vccd1 _13727_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__17502__A _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10938_ _10938_/A _10945_/A vssd1 vssd1 vccd1 vccd1 _10938_/Y sky130_fd_sc_hd__nand2_1
X_17494_ _17493_/A _21256_/A _17493_/C _17493_/D vssd1 vssd1 vccd1 vccd1 _17495_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__21370__B1 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18317__B _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19233_ _19231_/X _19233_/B vssd1 vssd1 vccd1 vccd1 _19234_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__14927__A1 _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16445_ _16989_/C _17013_/C vssd1 vssd1 vccd1 vccd1 _16449_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16627__A2_N _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14927__B2 _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10869_ hold140/A hold97/A vssd1 vssd1 vccd1 vccd1 _10871_/A sky130_fd_sc_hd__nor2_1
X_13657_ _13656_/B _13656_/C _13656_/A vssd1 vssd1 vccd1 vccd1 _13657_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_38_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11550__A _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19164_ _19000_/A _19000_/B _18839_/A _18839_/B _18836_/Y vssd1 vssd1 vccd1 vccd1
+ _19164_/X sky130_fd_sc_hd__o2111a_1
XFILLER_0_27_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20285__D _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12608_ _12728_/A vssd1 vssd1 vccd1 vccd1 _12610_/C sky130_fd_sc_hd__inv_2
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16376_ _16376_/A _16376_/B vssd1 vssd1 vccd1 vccd1 _16378_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13588_ _14367_/A _14384_/A _14212_/B _14195_/A vssd1 vssd1 vccd1 vccd1 _13591_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18115_ _18253_/B _18114_/C _18114_/A vssd1 vssd1 vccd1 vccd1 _18116_/B sky130_fd_sc_hd__o21ai_1
X_15327_ _15328_/A _15328_/B _15328_/C vssd1 vssd1 vccd1 vccd1 _15327_/Y sky130_fd_sc_hd__a21oi_4
X_19095_ _19095_/A _19095_/B _19095_/C vssd1 vssd1 vccd1 vccd1 _19097_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12539_ _12540_/A _12540_/B vssd1 vssd1 vccd1 vccd1 _12539_/X sky130_fd_sc_hd__and2_2
XFILLER_0_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18046_ _18046_/A _18046_/B vssd1 vssd1 vccd1 vccd1 _18082_/A sky130_fd_sc_hd__nand2_1
X_15258_ _16087_/A _15913_/B _15258_/C _15451_/A vssd1 vssd1 vccd1 vccd1 _15451_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14209_ _14209_/A _14209_/B vssd1 vssd1 vccd1 vccd1 _14228_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15189_ _14962_/Y _14965_/X _15346_/A _15188_/X vssd1 vssd1 vccd1 vccd1 _15346_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_10_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout408 _14698_/A vssd1 vssd1 vccd1 vccd1 _12020_/A sky130_fd_sc_hd__buf_4
Xfanout419 _15076_/B vssd1 vssd1 vccd1 vccd1 _14557_/B sky130_fd_sc_hd__clkbuf_8
X_19997_ _19997_/A _20138_/B _19997_/C vssd1 vssd1 vccd1 vccd1 _19999_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_10_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13666__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18948_ _19951_/A _19753_/B _19751_/C _19439_/A vssd1 vssd1 vccd1 vccd1 _18951_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13666__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16938__D _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18879_ _18878_/B _18878_/C _18867_/Y vssd1 vssd1 vccd1 vccd1 _18879_/Y sky130_fd_sc_hd__a21boi_2
XANTENNA__20103__A _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20910_ _20910_/A _21056_/B vssd1 vssd1 vccd1 vccd1 _20911_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_55_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21890_ _21926_/CLK _21890_/D vssd1 vssd1 vccd1 vccd1 hold215/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20841_ _20975_/D _20841_/B _20841_/C _20841_/D vssd1 vssd1 vccd1 vccd1 _20971_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__13969__A2 _13967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout163_A _17324_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20772_ hold226/X _20771_/X fanout2/X vssd1 vssd1 vccd1 vccd1 _21912_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout15 wire16/X vssd1 vssd1 vccd1 vccd1 _11545_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout26 _11348_/S vssd1 vssd1 vccd1 vccd1 _11284_/S sky130_fd_sc_hd__buf_8
XFILLER_0_119_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout37 _21490_/S vssd1 vssd1 vccd1 vccd1 _21536_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20476__C _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout48 fanout49/X vssd1 vssd1 vccd1 vccd1 fanout48/X sky130_fd_sc_hd__buf_4
XFILLER_0_64_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout330_A _21787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18109__A1 _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout59 _10791_/Y vssd1 vssd1 vccd1 vccd1 fanout59/X sky130_fd_sc_hd__buf_4
XFILLER_0_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout428_A _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14193__D _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21324_ _21324_/A _21324_/B vssd1 vssd1 vccd1 vccd1 _21324_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__15343__A1 _15192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21416__A1 _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21255_ _21255_/A _21255_/B vssd1 vssd1 vccd1 vccd1 _21257_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12291__A _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12722__C _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18897__B _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20206_ _20206_/A _20206_/B vssd1 vssd1 vccd1 vccd1 _20208_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21186_ _21186_/A _21186_/B vssd1 vssd1 vccd1 vccd1 _21231_/A sky130_fd_sc_hd__and2_1
XFILLER_0_25_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20137_ _20139_/A _20275_/B vssd1 vssd1 vccd1 vccd1 _20140_/A sky130_fd_sc_hd__or2_1
XFILLER_0_99_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout76_A _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17306__B _20249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20068_ _20069_/A _20069_/B vssd1 vssd1 vccd1 vccd1 _20068_/X sky130_fd_sc_hd__and2b_1
XTAP_3302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11910_ _11905_/A _11905_/B _11900_/A vssd1 vssd1 vccd1 vccd1 _11910_/X sky130_fd_sc_hd__o21ba_1
XTAP_3335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19802__A _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14606__B1 _10892_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12890_ _13010_/A _12889_/C _12889_/A vssd1 vssd1 vccd1 vccd1 _12891_/C sky130_fd_sc_hd__a21o_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_302 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_313 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_324 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ _11840_/A _11840_/B _11834_/A vssd1 vssd1 vccd1 vccd1 _11841_/Y sky130_fd_sc_hd__o21bai_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_335 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14560_ _14560_/A _14560_/B _14724_/B vssd1 vssd1 vccd1 vccd1 _14560_/X sky130_fd_sc_hd__and3_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11772_ _11772_/A _11772_/B _11772_/C vssd1 vssd1 vccd1 vccd1 _11772_/Y sky130_fd_sc_hd__nand3_2
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17020__A1 _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18137__B _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13511_ _13511_/A _13511_/B vssd1 vssd1 vccd1 vccd1 _13520_/A sky130_fd_sc_hd__xor2_4
XANTENNA__17020__B2 _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17041__B _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14491_ _14491_/A _14491_/B vssd1 vssd1 vccd1 vccd1 _14492_/B sky130_fd_sc_hd__xnor2_4
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15031__B1 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16230_ _16113_/Y _16115_/Y _16228_/X _16229_/Y vssd1 vssd1 vccd1 vccd1 _16302_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14384__C _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13442_ _14365_/A _15514_/A _15514_/B _14365_/D vssd1 vssd1 vccd1 vccd1 _13443_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_36_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12396__A1 _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13593__B1 _14212_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12396__B2 _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16161_ _16275_/A vssd1 vssd1 vccd1 vccd1 _16163_/D sky130_fd_sc_hd__inv_2
XFILLER_0_141_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13373_ _13373_/A _13373_/B vssd1 vssd1 vccd1 vccd1 _13398_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15112_ _16084_/A _16087_/A _15653_/C _15112_/D vssd1 vssd1 vccd1 vccd1 _15113_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_121_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14137__A2 _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12324_ _12401_/B _12324_/B vssd1 vssd1 vccd1 vccd1 _12334_/A sky130_fd_sc_hd__nor2_1
X_16092_ _14508_/A _21788_/Q hold319/A _16092_/D vssd1 vssd1 vccd1 vccd1 _16211_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_133_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15043_ _15044_/A _15044_/B _15044_/C vssd1 vssd1 vccd1 vccd1 _15043_/X sky130_fd_sc_hd__and3_1
XFILLER_0_50_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12255_ _12259_/A _12254_/B _12250_/X vssd1 vssd1 vccd1 vccd1 _12256_/C sky130_fd_sc_hd__a21oi_1
X_19920_ _19917_/X _19918_/Y _19759_/Y _19763_/C vssd1 vssd1 vccd1 vccd1 _19920_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_142_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11206_ hold178/X fanout22/X _11205_/X vssd1 vssd1 vccd1 vccd1 _11206_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_43_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18284__B1 _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19851_ _19951_/B _20247_/C _20247_/D _19951_/A vssd1 vssd1 vccd1 vccd1 _19854_/C
+ sky130_fd_sc_hd__a22o_1
X_12186_ _12267_/A _12242_/B _12246_/C _12246_/D vssd1 vssd1 vccd1 vccd1 _12199_/A
+ sky130_fd_sc_hd__and4_1
X_18802_ _18802_/A _18802_/B _18802_/C vssd1 vssd1 vccd1 vccd1 _18805_/A sky130_fd_sc_hd__nand3_1
X_11137_ hold196/X fanout23/X _11136_/X vssd1 vssd1 vccd1 vccd1 _11137_/X sky130_fd_sc_hd__a21o_1
X_19782_ _19782_/A _19782_/B vssd1 vssd1 vccd1 vccd1 _19785_/A sky130_fd_sc_hd__xnor2_1
X_16994_ _16994_/A _16994_/B _16994_/C vssd1 vssd1 vccd1 vccd1 _16994_/Y sky130_fd_sc_hd__nor3_2
XANTENNA__20813__A2_N _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18733_ _18733_/A _18733_/B vssd1 vssd1 vccd1 vccd1 _18735_/A sky130_fd_sc_hd__nor2_1
X_15945_ _15942_/A _15943_/Y _15776_/A _15777_/Y vssd1 vssd1 vccd1 vccd1 _15945_/X
+ sky130_fd_sc_hd__o211a_1
X_11068_ _10852_/X hold27/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21663_/D sky130_fd_sc_hd__mux2_1
X_18664_ _18664_/A _18664_/B _18664_/C vssd1 vssd1 vccd1 vccd1 _18664_/Y sky130_fd_sc_hd__nand3_1
X_15876_ _15741_/A _15740_/Y _15874_/X _15875_/Y vssd1 vssd1 vccd1 vccd1 _15876_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_118_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17615_ _17616_/A _17616_/B vssd1 vssd1 vccd1 vccd1 _17715_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_149_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14827_ _15931_/B _16409_/A _16328_/A _15931_/A vssd1 vssd1 vccd1 vccd1 _14830_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10882__A1 _10881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18595_ _19686_/B _19068_/C _19238_/C _19529_/B vssd1 vssd1 vccd1 vccd1 _18598_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17232__A _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17546_ _17546_/A _17546_/B vssd1 vssd1 vccd1 vccd1 _17548_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_47_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14758_ _14758_/A _14758_/B vssd1 vssd1 vccd1 vccd1 _14911_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_86_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13820__A1 _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13820__B2 _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13709_ _13864_/B _14354_/C _14663_/D _13867_/A vssd1 vssd1 vccd1 vccd1 _13709_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_128_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17477_ _17478_/A _17478_/B vssd1 vssd1 vccd1 vccd1 _17705_/A sky130_fd_sc_hd__nand2_1
X_14689_ _14689_/A _14689_/B vssd1 vssd1 vccd1 vccd1 _14743_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_11_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19216_ _19216_/A _19216_/B vssd1 vssd1 vccd1 vccd1 _19218_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16428_ _16173_/A _16284_/A _10794_/Y _16027_/B vssd1 vssd1 vccd1 vccd1 _16429_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11711__C _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19147_ _19143_/X _19144_/Y _18981_/X _18983_/X vssd1 vssd1 vccd1 vccd1 _19148_/C
+ sky130_fd_sc_hd__o211ai_2
X_16359_ _16359_/A _16359_/B vssd1 vssd1 vccd1 vccd1 _16360_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_14_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18063__A _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14128__A2 _14126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19078_ _19078_/A _19078_/B _19078_/C vssd1 vssd1 vccd1 vccd1 _19078_/X sky130_fd_sc_hd__and3_1
XFILLER_0_2_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18029_ _19823_/A _18767_/B _18616_/D _18030_/B vssd1 vssd1 vccd1 vccd1 _18031_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19067__A2 _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21040_ _21040_/A _21264_/A _21040_/C _21040_/D vssd1 vssd1 vccd1 vccd1 _21209_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_22_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout205 _19751_/C vssd1 vssd1 vccd1 vccd1 _19874_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_1_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout216 _21040_/A vssd1 vssd1 vccd1 vccd1 _19868_/B sky130_fd_sc_hd__buf_4
XANTENNA__15628__A2 _15626_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12261__D _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout227 hold324/X vssd1 vssd1 vccd1 vccd1 _20270_/C sky130_fd_sc_hd__clkbuf_8
Xfanout238 _17915_/D vssd1 vssd1 vccd1 vccd1 _19089_/B sky130_fd_sc_hd__buf_4
Xfanout249 _20583_/A vssd1 vssd1 vccd1 vccd1 _19379_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__17126__B _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout280_A _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15572__D _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18578__A1 _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout378_A _16284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18578__B2 _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21942_ _21942_/CLK _21942_/D vssd1 vssd1 vccd1 vccd1 hold185/A sky130_fd_sc_hd__dfxtp_1
X_21873_ _21938_/CLK hold103/X vssd1 vssd1 vccd1 vccd1 hold102/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1047 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout545_A _21734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20824_ _20824_/A _20824_/B _20824_/C vssd1 vssd1 vccd1 vccd1 _20824_/X sky130_fd_sc_hd__and3_2
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20755_ _20755_/A _20755_/B _20755_/C _20755_/D vssd1 vssd1 vccd1 vccd1 _20755_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_135_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18750__A1 _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16761__B1 _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20686_ _20686_/A _20686_/B vssd1 vssd1 vccd1 vccd1 _20694_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_17_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18404__C _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20653__D _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13829__B _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12733__B _13554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21307_ _21307_/A _21307_/B vssd1 vssd1 vccd1 vccd1 _21308_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19058__A2 _19060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12040_ _12040_/A _12040_/B _12040_/C vssd1 vssd1 vccd1 vccd1 _12093_/A sky130_fd_sc_hd__nand3_1
Xhold270 hold270/A vssd1 vssd1 vccd1 vccd1 hold270/X sky130_fd_sc_hd__dlygate4sd3_1
X_21238_ _21238_/A _21238_/B vssd1 vssd1 vccd1 vccd1 _21240_/B sky130_fd_sc_hd__and2_1
Xhold281 hold281/A vssd1 vssd1 vccd1 vccd1 hold281/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 hold312/A vssd1 vssd1 vccd1 vccd1 hold292/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11353__A2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21169_ _21169_/A _21169_/B vssd1 vssd1 vccd1 vccd1 _21171_/D sky130_fd_sc_hd__nand2_1
XANTENNA__14827__B1 _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13991_ _13992_/A _13992_/B _13992_/C vssd1 vssd1 vccd1 vccd1 _14284_/A sky130_fd_sc_hd__a21oi_4
X_15730_ _15599_/Y _15601_/Y _15728_/X _15729_/Y vssd1 vssd1 vccd1 vccd1 _15733_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_3110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12942_ _12942_/A _12961_/A _12942_/C vssd1 vssd1 vccd1 vccd1 _12961_/B sky130_fd_sc_hd__nand3_4
XTAP_3132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16044__A2 _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15661_ _16369_/A _16326_/A _15661_/C _15661_/D vssd1 vssd1 vccd1 vccd1 _15796_/B
+ sky130_fd_sc_hd__and4_1
XTAP_3165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_110 sstream_i[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12873_ _12744_/B _12744_/Y _12971_/A _12872_/Y vssd1 vssd1 vccd1 vccd1 _12971_/B
+ sky130_fd_sc_hd__o211ai_4
XTAP_3176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14676__A _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_121 v0z[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17400_ _17400_/A _17400_/B vssd1 vssd1 vccd1 vccd1 _17402_/B sky130_fd_sc_hd__xor2_2
XANTENNA_132 v1z[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14612_ _14492_/A _14492_/B _14490_/Y vssd1 vssd1 vccd1 vccd1 _14654_/A sky130_fd_sc_hd__o21ba_2
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_143 v1z[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17052__A _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18380_ _18230_/B _18230_/Y _18377_/X _18379_/Y vssd1 vssd1 vccd1 vccd1 _18380_/Y
+ sky130_fd_sc_hd__a211oi_4
X_11824_ _11795_/A _11795_/B _11795_/C vssd1 vssd1 vccd1 vccd1 _11824_/Y sky130_fd_sc_hd__a21oi_2
X_15592_ _15695_/A _15978_/B _15590_/Y _15713_/A vssd1 vssd1 vccd1 vccd1 _15594_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__21325__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_154 v2z[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_165 v2z[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_176 v2z[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_187 hold239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17331_ _17331_/A _17331_/B vssd1 vssd1 vccd1 vccd1 _17351_/A sky130_fd_sc_hd__xor2_2
X_14543_ _15375_/A _16418_/A _14543_/C _14543_/D vssd1 vssd1 vccd1 vccd1 _14543_/X
+ sky130_fd_sc_hd__and4_2
XANTENNA_198 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ _12261_/A _12269_/B _13157_/A _13017_/A vssd1 vssd1 vccd1 vccd1 _11758_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17544__A2 _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17262_ _16684_/Y _16686_/X _17363_/B _17261_/X vssd1 vssd1 vccd1 vccd1 _17264_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_37_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14474_ _14474_/A _14474_/B vssd1 vssd1 vccd1 vccd1 _14482_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11686_ _11685_/B _11685_/C _11685_/A vssd1 vssd1 vccd1 vccd1 _11701_/A sky130_fd_sc_hd__a21bo_1
X_19001_ _19001_/A _19001_/B vssd1 vssd1 vccd1 vccd1 _21373_/B sky130_fd_sc_hd__xnor2_4
X_16213_ _16213_/A _16213_/B vssd1 vssd1 vccd1 vccd1 _16221_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13425_ _13425_/A _13425_/B vssd1 vssd1 vccd1 vccd1 _13427_/C sky130_fd_sc_hd__xnor2_2
X_17193_ _17387_/A _20797_/A _17194_/A vssd1 vssd1 vccd1 vccd1 _17193_/X sky130_fd_sc_hd__and3_1
XFILLER_0_23_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15300__A _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16144_ _16144_/A _16144_/B vssd1 vssd1 vccd1 vccd1 _21412_/B sky130_fd_sc_hd__xnor2_2
X_13356_ _13352_/X _13354_/Y _13213_/B _13213_/Y vssd1 vssd1 vccd1 vccd1 _13357_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_10_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk_i _21806_/CLK vssd1 vssd1 vccd1 vccd1 _22063_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12307_ _12307_/A _12307_/B vssd1 vssd1 vccd1 vccd1 _12310_/A sky130_fd_sc_hd__xnor2_2
X_16075_ _16075_/A _16075_/B vssd1 vssd1 vccd1 vccd1 _16078_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_121_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18033__D _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13458__C _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13287_ _13287_/A _13287_/B vssd1 vssd1 vccd1 vccd1 _13306_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_87_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15026_ _15023_/X _15024_/Y _14816_/X _14819_/X vssd1 vssd1 vccd1 vccd1 _15027_/B
+ sky130_fd_sc_hd__a211o_1
X_19903_ _19903_/A _19903_/B vssd1 vssd1 vccd1 vccd1 _19911_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15954__B _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12238_ _12238_/A _12238_/B _12238_/C vssd1 vssd1 vccd1 vccd1 _12238_/X sky130_fd_sc_hd__and3_1
XANTENNA__17872__D _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12169_ _12168_/A _12167_/Y _12124_/X _12132_/Y vssd1 vssd1 vccd1 vccd1 _12169_/X
+ sky130_fd_sc_hd__o211a_1
X_19834_ _19830_/X _19831_/Y _19669_/B _19671_/B vssd1 vssd1 vccd1 vccd1 _19834_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__15673__C _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_28_clk_i clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21926_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__18009__B1 _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16977_ _16974_/Y _16983_/A _17096_/A _17124_/C vssd1 vssd1 vccd1 vccd1 _16983_/B
+ sky130_fd_sc_hd__and4bb_1
X_19765_ _19763_/X _19765_/B vssd1 vssd1 vccd1 vccd1 _19768_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_36_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15928_ _16027_/A _16177_/B _15769_/A _15767_/B vssd1 vssd1 vccd1 vccd1 _15936_/A
+ sky130_fd_sc_hd__a31o_1
X_18716_ _18716_/A _18716_/B vssd1 vssd1 vccd1 vccd1 _18718_/B sky130_fd_sc_hd__and2_1
X_19696_ _19534_/X _19537_/X _19693_/X _19695_/Y vssd1 vssd1 vccd1 vccd1 _19696_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11706__C _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18647_ _19587_/A _19587_/B _19866_/D vssd1 vssd1 vccd1 vccd1 _18647_/X sky130_fd_sc_hd__and3_1
X_15859_ _15859_/A _15859_/B vssd1 vssd1 vccd1 vccd1 _15860_/B sky130_fd_sc_hd__or2_1
XANTENNA__18058__A _18058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18578_ _19487_/A _18732_/C _19221_/C _19487_/B vssd1 vssd1 vccd1 vccd1 _18581_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13921__C _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17529_ _17529_/A _17529_/B vssd1 vssd1 vccd1 vccd1 _17532_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20540_ _20540_/A _20712_/A vssd1 vssd1 vccd1 vccd1 _20578_/A sky130_fd_sc_hd__or2_1
XFILLER_0_145_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20471_ _20471_/A _20471_/B vssd1 vssd1 vccd1 vccd1 _20491_/A sky130_fd_sc_hd__or2_1
XANTENNA__11032__A1 hold299/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15210__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20770__B _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22072_ _22080_/CLK _22072_/D fanout639/X vssd1 vssd1 vccd1 vccd1 mstream_o[8] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_1160 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout495_A _21745_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13665__A fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21023_ _20892_/A _20894_/X _21135_/B _21022_/X vssd1 vssd1 vccd1 vccd1 _21138_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_22_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11616__C _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21925_ _21932_/CLK _21925_/D vssd1 vssd1 vccd1 vccd1 hold155/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17303__C _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21856_ _21888_/CLK hold114/X vssd1 vssd1 vccd1 vccd1 hold113/A sky130_fd_sc_hd__dfxtp_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout39_A fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20807_ _20999_/B _20807_/B vssd1 vssd1 vccd1 vccd1 _20824_/A sky130_fd_sc_hd__and2_1
X_21787_ _21788_/CLK _21787_/D vssd1 vssd1 vccd1 vccd1 _21787_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11540_ _11089_/B t1y[30] t0x[30] _11543_/B2 vssd1 vssd1 vccd1 vccd1 _11540_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20738_ _20738_/A _20738_/B vssd1 vssd1 vccd1 vccd1 _20740_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout5_A fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19323__A2_N fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ _11123_/A t1y[7] t0x[7] _21724_/D vssd1 vssd1 vccd1 vccd1 _11471_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_34_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20669_ _21286_/A _21151_/A _20924_/A _21301_/A vssd1 vssd1 vccd1 vccd1 _20858_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_18_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11023__A1 hold258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13210_ _13230_/B _13209_/B _13209_/C _13209_/D vssd1 vssd1 vccd1 vccd1 _13210_/Y
+ sky130_fd_sc_hd__o22ai_4
XANTENNA__12220__B1 _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14190_ _14190_/A _14190_/B vssd1 vssd1 vccd1 vccd1 _14198_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13559__B _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13141_ _13140_/A _13140_/B _13140_/C vssd1 vssd1 vccd1 vccd1 _13142_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_21_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13072_ _13072_/A _13072_/B _13072_/C vssd1 vssd1 vccd1 vccd1 _13072_/X sky130_fd_sc_hd__or3_1
XFILLER_0_20_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16900_ _16951_/A _16997_/A vssd1 vssd1 vccd1 vccd1 _16952_/A sky130_fd_sc_hd__and2_1
X_12023_ _12023_/A _12071_/A vssd1 vssd1 vccd1 vccd1 _12077_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__19987__B1 _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16589__C _16870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17880_ _17746_/A _17745_/B _17743_/X vssd1 vssd1 vccd1 vccd1 _17881_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_40_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16265__A2 _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16831_ _17041_/A _17141_/C _17493_/A _16899_/B vssd1 vssd1 vccd1 vccd1 _16832_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13294__B _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout580 _21727_/Q vssd1 vssd1 vccd1 vccd1 _13525_/A sky130_fd_sc_hd__buf_4
Xfanout591 _11549_/A vssd1 vssd1 vccd1 vccd1 _11224_/A sky130_fd_sc_hd__buf_4
XANTENNA__19262__A _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19550_ _19549_/B _19700_/B _19549_/A vssd1 vssd1 vccd1 vccd1 _19551_/C sky130_fd_sc_hd__a21o_1
X_16762_ _16759_/X _16762_/B vssd1 vssd1 vccd1 vccd1 _16828_/B sky130_fd_sc_hd__and2b_1
X_13974_ _14138_/A _16328_/B _16399_/B _13975_/B vssd1 vssd1 vccd1 vccd1 _13974_/Y
+ sky130_fd_sc_hd__a22oi_1
X_18501_ _18500_/B _18500_/C _18500_/A vssd1 vssd1 vccd1 vccd1 _18503_/B sky130_fd_sc_hd__a21o_1
X_15713_ _15713_/A _15713_/B vssd1 vssd1 vccd1 vccd1 _15724_/A sky130_fd_sc_hd__or2_1
XFILLER_0_88_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12925_ _12924_/B _12924_/C _12924_/A vssd1 vssd1 vccd1 vccd1 _12925_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_77_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19481_ _19469_/A _19469_/B _19468_/A vssd1 vssd1 vccd1 vccd1 _19634_/A sky130_fd_sc_hd__a21bo_1
X_16693_ _16662_/A _16662_/C _16662_/B vssd1 vssd1 vccd1 vccd1 _16694_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_88_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18432_ _20317_/D _19644_/A _19227_/C _19227_/D vssd1 vssd1 vccd1 vccd1 _18588_/A
+ sky130_fd_sc_hd__and4_1
X_15644_ _15645_/A _15645_/B vssd1 vssd1 vccd1 vccd1 _15644_/Y sky130_fd_sc_hd__nand2_1
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12039__B1 _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12856_ _12856_/A _12856_/B vssd1 vssd1 vccd1 vccd1 _12865_/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18363_ _18363_/A _18363_/B _18363_/C vssd1 vssd1 vccd1 vccd1 _18363_/Y sky130_fd_sc_hd__nand3_2
X_11807_ _12458_/A _12357_/C _12444_/B _12443_/A vssd1 vssd1 vccd1 vccd1 _11810_/A
+ sky130_fd_sc_hd__nand4_1
X_15575_ _15702_/D _21787_/Q _15575_/C _15575_/D vssd1 vssd1 vccd1 vccd1 _15700_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_51_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12787_ _12787_/A _12787_/B _12787_/C vssd1 vssd1 vccd1 vccd1 _12790_/A sky130_fd_sc_hd__nand3_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17314_ _17315_/A _17315_/B vssd1 vssd1 vccd1 vccd1 _17314_/X sky130_fd_sc_hd__and2_2
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14526_ _14526_/A _14526_/B _14526_/C vssd1 vssd1 vccd1 vccd1 _14526_/X sky130_fd_sc_hd__and3_1
XANTENNA__11262__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11262__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18294_ _19373_/B _19068_/C _19238_/C _19051_/A vssd1 vssd1 vccd1 vccd1 _18294_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_44_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11738_ _12261_/A _12357_/C _13155_/B _13157_/A vssd1 vssd1 vccd1 vccd1 _11741_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_12_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17245_ _17245_/A _17245_/B _17245_/C vssd1 vssd1 vccd1 vccd1 _17248_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_71_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14457_ _14936_/D _14774_/D _16084_/D vssd1 vssd1 vccd1 vccd1 _14457_/X sky130_fd_sc_hd__and3_1
XFILLER_0_4_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11669_ _11670_/B _11670_/A vssd1 vssd1 vccd1 vccd1 _11669_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_71_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13408_ _13858_/A _13858_/B _14354_/C _14663_/D vssd1 vssd1 vccd1 vccd1 _13409_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_107_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17176_ _16721_/A _16721_/C _16721_/B vssd1 vssd1 vccd1 vccd1 _17267_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_148_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14388_ _15373_/B _14217_/D _15093_/B _15373_/A vssd1 vssd1 vccd1 vccd1 _14391_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16127_ _16127_/A _16127_/B vssd1 vssd1 vccd1 vccd1 _16128_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_109_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13339_ _13338_/B _13338_/C _13338_/A vssd1 vssd1 vccd1 vccd1 _13339_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_122_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20590__B _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19690__A2 _19692_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16058_ _16284_/A _16177_/B _16286_/B _16173_/A vssd1 vssd1 vccd1 vccd1 _16062_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14503__A2 _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15009_ _15006_/X _15007_/Y _14881_/B _14883_/B vssd1 vssd1 vccd1 vccd1 _15012_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16499__C _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19817_ _19818_/A _19818_/B vssd1 vssd1 vccd1 vccd1 _19817_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_155_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19748_ _20103_/A _19906_/D vssd1 vssd1 vccd1 vccd1 _19749_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14019__A1 _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19679_ _19679_/A _19679_/B vssd1 vssd1 vccd1 vccd1 _19681_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_56_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21710_ _22105_/CLK _21710_/D vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_154_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17123__C _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21641_ _21722_/CLK hold287/X fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[104]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout243_A _19692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11253__A1 _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11253__B2 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21572_ mstream_o[35] _11051_/Y _21579_/S vssd1 vssd1 vccd1 vccd1 _22099_/D sky130_fd_sc_hd__mux2_1
XANTENNA_10 _11331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_21 _11339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_32 _11412_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_43 _11445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20523_ _20910_/A _21256_/B _20523_/C _20523_/D vssd1 vssd1 vccd1 vccd1 _20686_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA_54 hold275/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout410_A _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12564__A _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16036__A _16036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_65 hold274/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_76 hold277/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout508_A _21742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_87 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_98 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20454_ _20845_/D _21286_/B _21296_/B _20721_/D vssd1 vssd1 vccd1 vccd1 _20458_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12753__A1 _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20385_ _20386_/A _20386_/B vssd1 vssd1 vccd1 vccd1 _20914_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22055_ _22063_/CLK _22055_/D vssd1 vssd1 vccd1 vccd1 hold270/A sky130_fd_sc_hd__dfxtp_4
XFILLER_0_101_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold288_A hold288/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21006_ _21005_/B _21005_/C _21005_/A vssd1 vssd1 vccd1 vccd1 _21006_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__17444__A1 _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17444__B2 _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21528__A0 hold270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19197__A1 _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19197__B2 _18894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10971_ _10971_/A _10971_/B vssd1 vssd1 vccd1 vccd1 _10972_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_134_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14657__C _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12710_ _12957_/B _12710_/B vssd1 vssd1 vccd1 vccd1 _21343_/B sky130_fd_sc_hd__xnor2_4
X_21908_ _21945_/CLK hold159/X vssd1 vssd1 vccd1 vccd1 hold158/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13561__C _21734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13690_ _13690_/A _13690_/B _13690_/C vssd1 vssd1 vccd1 vccd1 _13690_/X sky130_fd_sc_hd__and3_1
XANTENNA__11492__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12458__B _12785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12641_ _12641_/A _12641_/B vssd1 vssd1 vccd1 vccd1 _12651_/A sky130_fd_sc_hd__and2_1
X_21839_ _21845_/CLK _21839_/D vssd1 vssd1 vccd1 vccd1 _21839_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_93_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_21_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_400 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15360_ _15363_/A _15222_/B _15085_/A vssd1 vssd1 vccd1 vccd1 _15365_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_109_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12572_ _12572_/A _12572_/B _12572_/C vssd1 vssd1 vccd1 vccd1 _12575_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14311_ _14311_/A _14311_/B vssd1 vssd1 vccd1 vccd1 _14316_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12992__A1 _21735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20394__C _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12992__B2 _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11523_ _11544_/A1 t2x[24] v1z[24] fanout21/X _11522_/X vssd1 vssd1 vccd1 vccd1 _11523_/X
+ sky130_fd_sc_hd__a221o_1
X_15291_ _15292_/A _15292_/B vssd1 vssd1 vccd1 vccd1 _15291_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_110_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13595__A1_N _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17030_ _17030_/A vssd1 vssd1 vccd1 vccd1 _17058_/A sky130_fd_sc_hd__inv_2
X_14242_ _14713_/A _14713_/B _15234_/C vssd1 vssd1 vccd1 vccd1 _14242_/X sky130_fd_sc_hd__and3_1
XANTENNA__13289__B _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11454_ _21718_/D t2x[1] v1z[1] fanout17/X _11453_/X vssd1 vssd1 vccd1 vccd1 _11454_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14173_ _14173_/A _14173_/B vssd1 vssd1 vccd1 vccd1 _14273_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_1_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19257__A _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11385_ hold316/X fanout29/X _11384_/X vssd1 vssd1 vccd1 vccd1 _11385_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_150_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13124_ _13124_/A _13124_/B _13124_/C vssd1 vssd1 vccd1 vccd1 _13126_/A sky130_fd_sc_hd__and3_1
XANTENNA__16486__A2 _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18981_ _18815_/X _18817_/X _18979_/Y _18980_/X vssd1 vssd1 vccd1 vccd1 _18981_/X
+ sky130_fd_sc_hd__a211o_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15694__B1 _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ _13054_/A _13054_/B _13054_/C vssd1 vssd1 vccd1 vccd1 _13056_/C sky130_fd_sc_hd__a21o_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17932_ _17932_/A _17932_/B _17932_/C vssd1 vssd1 vccd1 vccd1 _17935_/A sky130_fd_sc_hd__nand3_1
XANTENNA__17435__A1 _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12006_ _12897_/C _12214_/C _12403_/B _12897_/D vssd1 vssd1 vccd1 vccd1 _12007_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17863_ _17861_/X _17863_/B vssd1 vssd1 vccd1 vccd1 _17864_/B sky130_fd_sc_hd__and2b_1
XANTENNA__17435__B2 _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14249__A1 _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11180__A0 _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19602_ _18789_/A _20242_/C _19603_/C _19729_/A vssd1 vssd1 vccd1 vccd1 _19604_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21519__A0 hold234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16814_ _16813_/A _17063_/C _17019_/C _17029_/B vssd1 vssd1 vccd1 vccd1 _16815_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17794_ _17794_/A _17794_/B _17794_/C vssd1 vssd1 vccd1 vccd1 _17797_/A sky130_fd_sc_hd__nand3_1
XANTENNA__20722__A1_N _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16745_ _16813_/A _16743_/C _17013_/D _16743_/B vssd1 vssd1 vccd1 vccd1 _16746_/B
+ sky130_fd_sc_hd__a22o_1
X_19533_ _19535_/A _20416_/A _20416_/B _19695_/A vssd1 vssd1 vccd1 vccd1 _19538_/C
+ sky130_fd_sc_hd__a22o_1
X_13957_ _13956_/B _13956_/C _13956_/A vssd1 vssd1 vccd1 vccd1 _13958_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_89_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17224__B _17417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17738__A2 _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12908_ _14384_/C _12907_/X _12906_/X vssd1 vssd1 vccd1 vccd1 _12909_/B sky130_fd_sc_hd__a21bo_1
X_19464_ _19464_/A _19464_/B vssd1 vssd1 vccd1 vccd1 _19465_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11483__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16676_ _16676_/A _16676_/B _16676_/C vssd1 vssd1 vccd1 vccd1 _16676_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13888_ _13730_/Y _13733_/X _13886_/Y _13887_/X vssd1 vssd1 vccd1 vccd1 _13948_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__20107__A1_N _20249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15627_ _21725_/D hold185/X _10946_/Y fanout5/X vssd1 vssd1 vccd1 vccd1 _15627_/X
+ sky130_fd_sc_hd__a22o_1
X_18415_ _18260_/X _18262_/Y _18413_/A _18414_/X vssd1 vssd1 vccd1 vccd1 _18415_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_124_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12839_ _13822_/B _13983_/B _14176_/C _13402_/D vssd1 vssd1 vccd1 vccd1 _12839_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_9_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19395_ _19395_/A _19395_/B _19395_/C vssd1 vssd1 vccd1 vccd1 _19398_/A sky130_fd_sc_hd__nand3_1
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18336__A _19732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11235__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18346_ _19438_/B _19868_/B _19414_/C _19438_/A vssd1 vssd1 vccd1 vccd1 _18347_/B
+ sky130_fd_sc_hd__a22o_1
X_15558_ _15558_/A _15558_/B vssd1 vssd1 vccd1 vccd1 _15560_/C sky130_fd_sc_hd__xnor2_1
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_126_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14509_ _14353_/X _14356_/X _14506_/X _14508_/Y vssd1 vssd1 vccd1 vccd1 _14509_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16174__A1 _16284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18277_ _18277_/A _18277_/B vssd1 vssd1 vccd1 vccd1 _18378_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15489_ _15490_/A _15490_/B vssd1 vssd1 vccd1 vccd1 _15625_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_12_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17228_ _17229_/A _17229_/B vssd1 vssd1 vccd1 vccd1 _17317_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17894__B _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15695__A _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17159_ _17159_/A _17159_/B _17159_/C _17159_/D vssd1 vssd1 vccd1 vccd1 _17159_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_13_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12534__D _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19663__A2 _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20170_ _20590_/D _20462_/D _20838_/C _20838_/D vssd1 vssd1 vccd1 vccd1 _20314_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__13927__B _21759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20106__A _21831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11171__A0 _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout193_A _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12559__A _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout458_A _21755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14477__C _14477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11474__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout625_A _21822_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17788__C _17924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11226__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21624_ _21939_/CLK _21624_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[87] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_90_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11226__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14493__B _14494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21555_ mstream_o[18] hold17/X _21562_/S vssd1 vssd1 vccd1 vccd1 _22082_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_105_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17300__D _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_2__f_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_2__f_clk_i/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_16_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20506_ _20503_/Y _20504_/X _20357_/Y _20359_/Y vssd1 vssd1 vccd1 vccd1 _20506_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15912__A1 _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14715__A2 _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21486_ hold202/X sstream_i[63] _21507_/S vssd1 vssd1 vccd1 vccd1 _22013_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_99_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12444__D _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20437_ _20438_/A _20438_/B vssd1 vssd1 vccd1 vccd1 _20571_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_114_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11170_ hold198/X fanout22/X _11169_/X vssd1 vssd1 vccd1 vccd1 _11170_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13837__B _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20368_ _20220_/A _20220_/B _20221_/X vssd1 vssd1 vccd1 vccd1 _20370_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_105_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19227__D _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20299_ _20299_/A _20299_/B vssd1 vssd1 vccd1 vccd1 _20301_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_101_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13151__A1 _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22038_ _22038_/CLK _22038_/D vssd1 vssd1 vccd1 vccd1 hold271/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13151__B2 _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14860_ _14860_/A _14860_/B _14976_/B vssd1 vssd1 vccd1 vccd1 _14862_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_89_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13811_ _13818_/B _13809_/Y _13656_/B _13656_/Y vssd1 vssd1 vccd1 vccd1 _13812_/B
+ sky130_fd_sc_hd__a211o_1
X_14791_ _14791_/A _14791_/B _14946_/B vssd1 vssd1 vccd1 vccd1 _14793_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_98_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16530_ _16530_/A _16530_/B vssd1 vssd1 vccd1 vccd1 _16531_/B sky130_fd_sc_hd__nor2_1
X_13742_ _14365_/A _14367_/A _14384_/A _14212_/B vssd1 vssd1 vccd1 vccd1 _13743_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__11465__A1 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10954_ hold78/A hold276/A _10952_/X _10953_/Y vssd1 vssd1 vccd1 vccd1 _10959_/A
+ sky130_fd_sc_hd__a211o_2
XANTENNA__11465__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16883__B _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16461_ _16743_/C _16460_/X _16459_/X vssd1 vssd1 vccd1 vccd1 _16462_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13673_ _13985_/A _16404_/B vssd1 vssd1 vccd1 vccd1 _13674_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12619__D _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10885_ _10885_/A _10885_/B _10885_/C vssd1 vssd1 vccd1 vccd1 _10886_/B sky130_fd_sc_hd__and3_1
XFILLER_0_156_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18200_ _18200_/A _18200_/B vssd1 vssd1 vccd1 vccd1 _18209_/A sky130_fd_sc_hd__xnor2_2
X_15412_ _15547_/A _16040_/C _15933_/C _15412_/D vssd1 vssd1 vccd1 vccd1 _15547_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_39_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19180_ _19013_/C _19179_/X _19178_/X vssd1 vssd1 vccd1 vccd1 _19182_/A sky130_fd_sc_hd__a21bo_2
X_12624_ _12732_/B _12622_/X _12530_/C _12532_/A vssd1 vssd1 vccd1 vccd1 _12625_/B
+ sky130_fd_sc_hd__o211ai_1
X_16392_ _16392_/A _16392_/B vssd1 vssd1 vccd1 vccd1 _16393_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18131_ _18849_/A _18849_/B _19221_/C vssd1 vssd1 vccd1 vccd1 _18131_/X sky130_fd_sc_hd__and3_1
X_15343_ _15192_/A _15192_/B _15151_/A vssd1 vssd1 vccd1 vccd1 _15345_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_109_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16156__A1 _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12555_ _12556_/A _12556_/B vssd1 vssd1 vccd1 vccd1 _12653_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_124_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11312__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11506_ _11505_/X _19227_/C _11545_/S vssd1 vssd1 vccd1 vccd1 _21840_/D sky130_fd_sc_hd__mux2_1
X_18062_ _18062_/A _18062_/B vssd1 vssd1 vccd1 vccd1 _18071_/A sky130_fd_sc_hd__xnor2_2
X_15274_ _15931_/A _15931_/B _16040_/C _16396_/A vssd1 vssd1 vccd1 vccd1 _15406_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12486_ _12381_/Y _12383_/Y _12484_/X _12485_/Y vssd1 vssd1 vccd1 vccd1 _12825_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_145_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17013_ _17146_/A _17141_/B _17013_/C _17013_/D vssd1 vssd1 vccd1 vccd1 _17016_/A
+ sky130_fd_sc_hd__nand4_2
X_14225_ _14224_/B _14224_/C _14224_/A vssd1 vssd1 vccd1 vccd1 _14226_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_34_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11437_ _11436_/X _21278_/B _11470_/S vssd1 vssd1 vccd1 vccd1 _21817_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_123_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16404__A _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16459__A2 _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17656__A1 _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14156_ _14306_/A _16328_/B _14157_/C _14157_/D vssd1 vssd1 vccd1 vccd1 _14156_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17656__B2 _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11368_ _11367_/X _17086_/C _11401_/S vssd1 vssd1 vccd1 vccd1 _21794_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_42_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11548__A _11549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13107_ _13107_/A _13244_/B vssd1 vssd1 vccd1 vccd1 _13109_/A sky130_fd_sc_hd__or2_1
XFILLER_0_81_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14087_ _14087_/A _14250_/B vssd1 vssd1 vccd1 vccd1 _14090_/A sky130_fd_sc_hd__nand2_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18964_ _18964_/A _18964_/B _18964_/C vssd1 vssd1 vccd1 vccd1 _18967_/A sky130_fd_sc_hd__or3_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ fanout58/X v0z[18] fanout18/X _11298_/X vssd1 vssd1 vccd1 vccd1 _11299_/X
+ sky130_fd_sc_hd__a31o_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ _13038_/A _13169_/B _13038_/C vssd1 vssd1 vccd1 vccd1 _13040_/B sky130_fd_sc_hd__nand3_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17915_ _17915_/A _18787_/A _18787_/B _17915_/D vssd1 vssd1 vccd1 vccd1 _18047_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__11153__A0 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18895_ _18895_/A _18895_/B vssd1 vssd1 vccd1 vccd1 _18905_/A sky130_fd_sc_hd__and2_1
XANTENNA__14859__A _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17846_ _17847_/A _17847_/B _17847_/C vssd1 vssd1 vccd1 vccd1 _18127_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14989_ _14990_/A _14990_/B _14990_/C vssd1 vssd1 vccd1 vccd1 _15012_/A sky130_fd_sc_hd__a21oi_2
X_17777_ _17777_/A _17777_/B vssd1 vssd1 vccd1 vccd1 _17785_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13913__D _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18908__A1 _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18908__B2 _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11456__A1 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19516_ _19356_/B _19358_/B _19676_/A _19515_/Y vssd1 vssd1 vccd1 vccd1 _19676_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_152_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16728_ _16727_/B _16727_/C _16727_/A vssd1 vssd1 vccd1 vccd1 _16730_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__11456__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16659_ _17141_/A _17141_/B _17434_/B _17433_/A vssd1 vssd1 vccd1 vccd1 _16662_/A
+ sky130_fd_sc_hd__nand4_1
X_19447_ _19448_/B _19448_/A vssd1 vssd1 vccd1 vccd1 _19447_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_14_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_119_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19378_ _19535_/B _19379_/B _20416_/A _19691_/D vssd1 vssd1 vccd1 vccd1 _19378_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18136__A2 _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18329_ _18176_/X _18178_/X _18327_/X _18328_/Y vssd1 vssd1 vccd1 vccd1 _18368_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11730__B _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11222__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21340_ _21349_/A _21340_/B vssd1 vssd1 vccd1 vccd1 _21340_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17895__A1 _18030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17895__B2 _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21271_ _21271_/A _21271_/B vssd1 vssd1 vccd1 vccd1 _21281_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16314__A _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout206_A _21816_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20222_ _20222_/A _20222_/B _20220_/Y vssd1 vssd1 vccd1 vccd1 _20223_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17129__B _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20153_ _20153_/A _20153_/B vssd1 vssd1 vccd1 vccd1 _20156_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13133__A1 _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20084_ _19636_/A _15210_/B _21393_/B _20770_/B vssd1 vssd1 vccd1 vccd1 _20084_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11144__A0 _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13673__A _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17145__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11695__A1 _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16083__B1 _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14633__A1 _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11447__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12644__B1 _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20986_ _20986_/A _20986_/B vssd1 vssd1 vccd1 vccd1 _20994_/A sky130_fd_sc_hd__nand2_1
XANTENNA__16386__A1 _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout21_A _11224_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19324__A1 _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15702__A_N _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21607_ _21906_/CLK _21607_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[70] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11132__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12340_ _12899_/B _12637_/A _11713_/B _11711_/X vssd1 vssd1 vccd1 vccd1 _12350_/A
+ sky130_fd_sc_hd__a31o_1
X_21538_ mstream_o[1] hold9/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22065_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_63_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1016 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14951__B _15174_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12271_ _12271_/A _12271_/B vssd1 vssd1 vccd1 vccd1 _12271_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_65_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21469_ hold198/X sstream_i[46] _21481_/S vssd1 vssd1 vccd1 vccd1 _21996_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19238__C _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14010_ _14007_/Y _14008_/Y _13845_/Y _13847_/Y vssd1 vssd1 vccd1 vccd1 _14011_/D
+ sky130_fd_sc_hd__a211oi_2
X_11222_ hold313/X _11221_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21757_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17638__A1 _18008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17638__B2 _18008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19535__A _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11153_ _12637_/B _11152_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21734_/D sky130_fd_sc_hd__mux2_1
X_15961_ _14813_/A _21788_/Q hold319/A _15961_/D vssd1 vssd1 vccd1 vccd1 _15964_/A
+ sky130_fd_sc_hd__and4b_2
X_11084_ _10965_/Y hold56/X _11084_/S vssd1 vssd1 vccd1 vccd1 _21679_/D sky130_fd_sc_hd__mux2_1
XANTENNA__11135__A0 _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21198__A1 _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18796__D _19753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14872__A1 _15093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14912_ _14913_/B vssd1 vssd1 vccd1 vccd1 _14912_/Y sky130_fd_sc_hd__inv_2
X_17700_ _17700_/A _17700_/B vssd1 vssd1 vccd1 vccd1 _17703_/A sky130_fd_sc_hd__nand2_2
XANTENNA__17055__A _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15892_ _15892_/A _15892_/B _16027_/B vssd1 vssd1 vccd1 vccd1 _15894_/A sky130_fd_sc_hd__and3_1
XANTENNA__12883__B1 _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18680_ _18525_/C _18525_/Y _18678_/X _18679_/X vssd1 vssd1 vccd1 vccd1 _18682_/A
+ sky130_fd_sc_hd__o211a_1
X_14843_ _14840_/Y _14841_/X _14709_/A _14710_/Y vssd1 vssd1 vccd1 vccd1 _14844_/C
+ sky130_fd_sc_hd__a211o_1
X_17631_ _17630_/B _17630_/C _17630_/A vssd1 vssd1 vccd1 vccd1 _17631_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_98_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11438__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17562_ _17562_/A _17562_/B _17562_/C vssd1 vssd1 vccd1 vccd1 _17564_/B sky130_fd_sc_hd__nand3_1
XANTENNA__19012__B1 _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14774_ _14621_/D _15838_/B _16314_/D _14774_/D vssd1 vssd1 vccd1 vccd1 _14777_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_58_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11986_ _11986_/A _11986_/B _11986_/C vssd1 vssd1 vccd1 vccd1 _12043_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_58_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16513_ _16989_/C _17619_/A _16512_/C _16564_/A vssd1 vssd1 vccd1 vccd1 _16513_/X
+ sky130_fd_sc_hd__a22o_1
X_19301_ _19139_/A _19139_/C _19139_/B vssd1 vssd1 vccd1 vccd1 _19303_/B sky130_fd_sc_hd__a21bo_1
X_13725_ _13591_/D _13592_/B _13723_/Y _13724_/X vssd1 vssd1 vccd1 vccd1 _13883_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__21305__A _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10937_ hold79/A hold101/A vssd1 vssd1 vccd1 vccd1 _10945_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17502__B _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17493_ _17493_/A _21256_/A _17493_/C _17493_/D vssd1 vssd1 vccd1 vccd1 _17614_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__21370__A1 _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14388__B1 _15093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15303__A _15439_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16444_ _16444_/A _16697_/A vssd1 vssd1 vccd1 vccd1 _16456_/A sky130_fd_sc_hd__nor2_1
X_19232_ _19228_/X _19230_/Y _19056_/X _19059_/X vssd1 vssd1 vccd1 vccd1 _19233_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_156_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14927__A2 _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13656_ _13656_/A _13656_/B _13656_/C vssd1 vssd1 vccd1 vccd1 _13656_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_14_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10868_ mstream_o[45] _10867_/X _10992_/S vssd1 vssd1 vccd1 vccd1 _21582_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_27_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11550__B _11550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19163_ _19161_/Y _19163_/B vssd1 vssd1 vccd1 vccd1 _19788_/A sky130_fd_sc_hd__nand2b_2
X_12607_ _13682_/C _13822_/B _21776_/Q _13258_/D vssd1 vssd1 vccd1 vccd1 _12728_/A
+ sky130_fd_sc_hd__and4_1
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16375_ _16333_/A _16332_/B _16330_/Y vssd1 vssd1 vccd1 vccd1 _16376_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13587_ _13583_/X _13584_/Y _13428_/A _13428_/Y vssd1 vssd1 vccd1 vccd1 _13648_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_87_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ mstream_o[114] _10790_/Y _11027_/S vssd1 vssd1 vccd1 vccd1 _21722_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_82_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20863__B _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18114_ _18114_/A _18253_/B _18114_/C vssd1 vssd1 vccd1 vccd1 _18114_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15326_ _15326_/A _15326_/B vssd1 vssd1 vccd1 vccd1 _15328_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19094_ _19095_/A _19095_/B _19095_/C vssd1 vssd1 vccd1 vccd1 _19097_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_42_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12538_ _12750_/A _13157_/B _12429_/B _12427_/X vssd1 vssd1 vccd1 vccd1 _12540_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__15957__B _21787_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21040__A _21040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18045_ _18044_/B _18044_/C _18044_/A vssd1 vssd1 vccd1 vccd1 _18046_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15257_ _16087_/A _15913_/B _15258_/C _15451_/A vssd1 vssd1 vccd1 vccd1 _15259_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12469_ _12468_/A _12468_/B _12468_/C vssd1 vssd1 vccd1 vccd1 _12471_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_112_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14208_ _14208_/A _14208_/B vssd1 vssd1 vccd1 vccd1 _14268_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_111_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15188_ _15296_/B _15186_/X _15046_/Y _15050_/C vssd1 vssd1 vccd1 vccd1 _15188_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11913__A2 _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14139_ _16084_/D _14138_/X _14137_/X vssd1 vssd1 vccd1 vccd1 _14141_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__19445__A _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout409 _14698_/A vssd1 vssd1 vccd1 vccd1 _13155_/C sky130_fd_sc_hd__buf_4
X_19996_ _19898_/A _19898_/C _19898_/B vssd1 vssd1 vccd1 vccd1 _19997_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18947_ _18947_/A _18947_/B vssd1 vssd1 vccd1 vccd1 _18955_/A sky130_fd_sc_hd__nand2_1
XANTENNA__21189__A1 _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21189__B2 _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11677__A1 _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18878_ _18867_/Y _18878_/B _18878_/C vssd1 vssd1 vccd1 vccd1 _18878_/X sky130_fd_sc_hd__and3b_2
XANTENNA__20103__B _21815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17829_ _17830_/A _17830_/B _17837_/B vssd1 vssd1 vccd1 vccd1 _17831_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__11725__B _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19003__B1 _14126_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11429__A1 _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20840_ _20975_/D _21291_/B _20841_/C _20841_/D vssd1 vssd1 vccd1 vccd1 _20842_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_49_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20771_ _11550_/B _15888_/Y _20769_/Y _11550_/A _20770_/X vssd1 vssd1 vccd1 vccd1
+ _20771_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_18_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout156_A _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout27 _11348_/S vssd1 vssd1 vccd1 vccd1 _11352_/S sky130_fd_sc_hd__buf_6
Xfanout38 _21422_/X vssd1 vssd1 vccd1 vccd1 _21490_/S sky130_fd_sc_hd__buf_4
XANTENNA__20476__D _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout49 _11123_/X vssd1 vssd1 vccd1 vccd1 fanout49/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18109__A2 _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout323_A _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21323_ _21323_/A _21323_/B vssd1 vssd1 vccd1 vccd1 _21324_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21254_ _21247_/B _21248_/A _21253_/X _21246_/B vssd1 vssd1 vccd1 vccd1 _21324_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12291__B _12291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18897__C _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20205_ _20205_/A _20205_/B vssd1 vssd1 vccd1 vccd1 _20206_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_64_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12722__D _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21185_ _21185_/A _21185_/B vssd1 vssd1 vccd1 vccd1 _21186_/B sky130_fd_sc_hd__or2_1
XFILLER_0_111_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20136_ _21291_/A _20419_/A _20136_/C _20136_/D vssd1 vssd1 vccd1 vccd1 _20275_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__11117__A0 _10965_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14499__A _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20067_ _19929_/A _19929_/B _19927_/X vssd1 vssd1 vccd1 vccd1 _20069_/B sky130_fd_sc_hd__a21o_1
XANTENNA_hold270_A hold270/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout69_A _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19802__B _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14606__A1 _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14606__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_303 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _11840_/A _11840_/B _11834_/A vssd1 vssd1 vccd1 vccd1 _11840_/X sky130_fd_sc_hd__or3b_1
XANTENNA_314 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_325 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_336 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19545__A1 _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19545__B2 _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _11772_/A _11772_/B _11772_/C vssd1 vssd1 vccd1 vccd1 _11771_/X sky130_fd_sc_hd__and3_1
XFILLER_0_68_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20969_ _21087_/D _21291_/B _20969_/C _20969_/D vssd1 vssd1 vccd1 vccd1 _21085_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_68_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13510_ _13511_/A _13511_/B vssd1 vssd1 vccd1 vccd1 _13662_/A sky130_fd_sc_hd__or2_2
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17020__A2 _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14490_ _14491_/A _14491_/B vssd1 vssd1 vccd1 vccd1 _14490_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_95_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15031__A1 _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15031__B2 _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14384__D _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13441_ _14365_/A _15514_/B _14365_/D _15514_/A vssd1 vssd1 vccd1 vccd1 _13443_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16160_ _16380_/A _16371_/A _21753_/Q _16369_/B vssd1 vssd1 vccd1 vccd1 _16275_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__13593__A1 _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12396__A2 _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13593__B2 _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13372_ _13361_/A _13512_/A _13361_/C _13518_/C _13368_/B vssd1 vssd1 vccd1 vccd1
+ _13513_/A sky130_fd_sc_hd__o32a_2
XFILLER_0_23_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15111_ _16084_/A _15653_/C _15112_/D _16087_/A vssd1 vssd1 vccd1 vccd1 _15115_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12323_ _12403_/A _13012_/B _12320_/Y _12322_/B vssd1 vssd1 vccd1 vccd1 _12324_/B
+ sky130_fd_sc_hd__a22oi_1
X_16091_ _16091_/A _16091_/B vssd1 vssd1 vccd1 vccd1 _16095_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_121_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15042_ _15040_/A _15040_/B _15040_/C vssd1 vssd1 vccd1 vccd1 _15044_/C sky130_fd_sc_hd__a21o_1
X_12254_ _12250_/X _12254_/B vssd1 vssd1 vccd1 vccd1 _12259_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_121_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11205_ hold119/X fanout51/X fanout48/X hold272/A vssd1 vssd1 vccd1 vccd1 _11205_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18284__A1 _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19850_ _19723_/A _19723_/C _19586_/X vssd1 vssd1 vccd1 vccd1 _20091_/A sky130_fd_sc_hd__a21o_2
XFILLER_0_102_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18284__B2 _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12185_ _12185_/A _12185_/B _12185_/C vssd1 vssd1 vccd1 vccd1 _12193_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18801_ _19123_/A _19123_/B _21258_/B _20247_/C vssd1 vssd1 vccd1 vccd1 _18802_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA__11108__A0 _10903_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ hold317/X _11126_/A _11126_/B hold192/X vssd1 vssd1 vccd1 vccd1 _11136_/X
+ sky130_fd_sc_hd__a22o_1
X_19781_ _19782_/A _19782_/B vssd1 vssd1 vccd1 vccd1 _19942_/B sky130_fd_sc_hd__nand2_1
X_16993_ _16982_/A _16982_/B _16982_/C vssd1 vssd1 vccd1 vccd1 _16994_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__18036__A1 _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18732_ _19644_/A _19487_/A _18732_/C _18894_/B vssd1 vssd1 vccd1 vccd1 _18733_/B
+ sky130_fd_sc_hd__and4_1
X_15944_ _15776_/A _15777_/Y _15942_/A _15943_/Y vssd1 vssd1 vccd1 vccd1 _15944_/Y
+ sky130_fd_sc_hd__a211oi_4
X_11067_ _11066_/Y hold81/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21662_/D sky130_fd_sc_hd__mux2_1
X_15875_ _15874_/A _15874_/B _15874_/C _15874_/D vssd1 vssd1 vccd1 vccd1 _15875_/Y
+ sky130_fd_sc_hd__o22ai_2
X_18663_ _18664_/A _18664_/B _18664_/C vssd1 vssd1 vccd1 vccd1 _18663_/X sky130_fd_sc_hd__and3_1
XFILLER_0_153_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14826_ _16027_/A _16328_/A _14692_/X _14693_/X _16418_/A vssd1 vssd1 vccd1 vccd1
+ _14831_/A sky130_fd_sc_hd__a32o_1
X_17614_ _17614_/A _17614_/B vssd1 vssd1 vccd1 vccd1 _17616_/B sky130_fd_sc_hd__or2_2
XFILLER_0_116_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18594_ _18594_/A _18594_/B vssd1 vssd1 vccd1 vccd1 _18603_/A sky130_fd_sc_hd__or2_1
XTAP_3870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19536__A1 _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14757_ _14758_/A _14758_/B vssd1 vssd1 vccd1 vccd1 _14757_/Y sky130_fd_sc_hd__nand2_1
X_17545_ _19951_/A _17543_/X _17544_/X vssd1 vssd1 vccd1 vccd1 _17546_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__17232__B _18058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11969_ _11969_/A _11969_/B _11969_/C vssd1 vssd1 vccd1 vccd1 _11970_/B sky130_fd_sc_hd__or3_1
XFILLER_0_114_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13820__A2 _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13708_ _13708_/A _13708_/B vssd1 vssd1 vccd1 vccd1 _13718_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17476_ _17366_/A _17366_/B _17364_/Y vssd1 vssd1 vccd1 vccd1 _17478_/B sky130_fd_sc_hd__o21ai_2
X_14688_ _14688_/A _14688_/B vssd1 vssd1 vccd1 vccd1 _14689_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_74_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19215_ _19216_/B _19216_/A vssd1 vssd1 vccd1 vccd1 _19327_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_156_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16427_ _16286_/B _16283_/A _16286_/D _16027_/B _16286_/A vssd1 vssd1 vccd1 vccd1
+ _16429_/A sky130_fd_sc_hd__o2111a_1
XFILLER_0_128_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13639_ _13638_/B _13638_/C _13638_/A vssd1 vssd1 vccd1 vccd1 _13639_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__18344__A _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11711__D _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16358_ _16359_/A _16359_/B vssd1 vssd1 vccd1 vccd1 _16360_/A sky130_fd_sc_hd__and2_1
X_19146_ _18981_/X _18983_/X _19143_/X _19144_/Y vssd1 vssd1 vccd1 vccd1 _19148_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15309_ _21735_/Q _15838_/B _16374_/B _15159_/D vssd1 vssd1 vccd1 vccd1 _15310_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_14_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16289_ _16289_/A _16289_/B vssd1 vssd1 vccd1 vccd1 _16290_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_125_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19077_ _19076_/A _19076_/B _19076_/C vssd1 vssd1 vccd1 vccd1 _19078_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12392__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11500__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18028_ _19664_/B _18769_/B vssd1 vssd1 vccd1 vccd1 _18032_/A sky130_fd_sc_hd__and2_1
XFILLER_0_2_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11347__B1 _11346_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout206 _21816_/Q vssd1 vssd1 vccd1 vccd1 _19751_/C sky130_fd_sc_hd__buf_4
Xfanout217 _21040_/A vssd1 vssd1 vccd1 vccd1 _21305_/A sky130_fd_sc_hd__buf_4
Xfanout228 _19703_/C vssd1 vssd1 vccd1 vccd1 _19546_/D sky130_fd_sc_hd__buf_4
XFILLER_0_5_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout239 _17915_/D vssd1 vssd1 vccd1 vccd1 _19692_/B sky130_fd_sc_hd__clkbuf_4
X_19979_ _19979_/A _20098_/B _19979_/C vssd1 vssd1 vccd1 vccd1 _20126_/A sky130_fd_sc_hd__and3_1
XANTENNA__18578__A2 _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21941_ _21942_/CLK _21941_/D vssd1 vssd1 vccd1 vccd1 hold95/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout273_A _21800_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21872_ _21938_/CLK hold84/X vssd1 vssd1 vccd1 vccd1 hold83/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_82_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20823_ _20823_/A _20823_/B _20823_/C vssd1 vssd1 vccd1 vccd1 _20824_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_82_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout440_A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout538_A _15439_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20754_ _20750_/Y _20751_/X _20621_/B _20621_/Y vssd1 vssd1 vccd1 vccd1 _20755_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18750__A2 _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20685_ _20685_/A _20685_/B vssd1 vssd1 vccd1 vccd1 _20696_/A sky130_fd_sc_hd__or2_1
XFILLER_0_134_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21098__B1 _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11586__B1 _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18404__D _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16513__A1 _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11410__S _11446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12733__C _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21306_ _21163_/A _21163_/B _21162_/A vssd1 vssd1 vccd1 vccd1 _21307_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_66_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21237_ _21255_/B _21237_/B vssd1 vssd1 vccd1 vccd1 _21240_/A sky130_fd_sc_hd__nand2_1
Xhold260 hold260/A vssd1 vssd1 vccd1 vccd1 hold260/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 hold271/A vssd1 vssd1 vccd1 vccd1 hold271/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 hold282/A vssd1 vssd1 vccd1 vccd1 hold282/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold293 hold293/A vssd1 vssd1 vccd1 vccd1 hold293/X sky130_fd_sc_hd__dlygate4sd3_1
X_21168_ _21168_/A vssd1 vssd1 vccd1 vccd1 _21171_/C sky130_fd_sc_hd__inv_2
XANTENNA__14827__A1 _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14827__B2 _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_9_clk_i _21806_/CLK vssd1 vssd1 vccd1 vccd1 _22005_/CLK sky130_fd_sc_hd__clkbuf_16
X_20119_ _20119_/A _20119_/B vssd1 vssd1 vccd1 vccd1 _20121_/B sky130_fd_sc_hd__xnor2_2
X_13990_ _14149_/B _13990_/B vssd1 vssd1 vccd1 vccd1 _13992_/C sky130_fd_sc_hd__nand2_1
X_21099_ _21286_/A _21311_/A _21283_/B _21305_/B vssd1 vssd1 vccd1 vccd1 _21208_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_102_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12941_ _12938_/Y _12939_/X _12813_/B _12812_/Y vssd1 vssd1 vccd1 vccd1 _12942_/C
+ sky130_fd_sc_hd__a211o_1
XTAP_3111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21573__A1 _11053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18429__A _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15660_ _16369_/A _16326_/A _15661_/C _15661_/D vssd1 vssd1 vccd1 vccd1 _15662_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_3144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_100 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12872_ _12869_/X _12870_/Y _12765_/X _12768_/Y vssd1 vssd1 vccd1 vccd1 _12872_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_3166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_111 sstream_i[64] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14611_ _14611_/A _14611_/B vssd1 vssd1 vccd1 vccd1 _14751_/A sky130_fd_sc_hd__or2_2
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_122 v0z[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_133 v1z[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11823_ _11823_/A _11823_/B _11823_/C vssd1 vssd1 vccd1 vccd1 _11823_/Y sky130_fd_sc_hd__nand3_2
X_15591_ _16374_/A _16087_/A _15717_/C _15976_/D vssd1 vssd1 vccd1 vccd1 _15713_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17052__B _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_144 v1z[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21325__A1 _11550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_155 v2z[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_166 v2z[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17330_ _17331_/A _17331_/B vssd1 vssd1 vccd1 vccd1 _17427_/B sky130_fd_sc_hd__nand2_2
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14542_ _15375_/A _16418_/A _14543_/C _14543_/D vssd1 vssd1 vccd1 vccd1 _14542_/Y
+ sky130_fd_sc_hd__a22oi_2
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_177 v2z[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_188 hold239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11754_ _11753_/B _11753_/C _11753_/A vssd1 vssd1 vccd1 vccd1 _11754_/Y sky130_fd_sc_hd__a21oi_2
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_199 hold268/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15788__A _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17261_ _17363_/A _17260_/C _17260_/A vssd1 vssd1 vccd1 vccd1 _17261_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_37_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14473_ _14361_/A _14360_/B _14358_/X vssd1 vssd1 vccd1 vccd1 _14473_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11685_ _11685_/A _11685_/B _11685_/C vssd1 vssd1 vccd1 vccd1 _11770_/A sky130_fd_sc_hd__and3_1
XFILLER_0_71_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16212_ _16212_/A _16212_/B vssd1 vssd1 vccd1 vccd1 _16223_/A sky130_fd_sc_hd__or2_1
X_19000_ _19000_/A _19000_/B vssd1 vssd1 vccd1 vccd1 _19001_/B sky130_fd_sc_hd__nor2_2
X_13424_ _13425_/A _13425_/B vssd1 vssd1 vccd1 vccd1 _13580_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_154_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17192_ _17387_/A _20797_/A vssd1 vssd1 vccd1 vccd1 _17194_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_24_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16143_ _16143_/A _16143_/B vssd1 vssd1 vccd1 vccd1 _16144_/B sky130_fd_sc_hd__or2_1
XFILLER_0_106_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15300__B _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13355_ _13213_/B _13213_/Y _13352_/X _13354_/Y vssd1 vssd1 vccd1 vccd1 _13509_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_107_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11320__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14515__B1 _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12306_ _12306_/A _12306_/B vssd1 vssd1 vccd1 vccd1 _12307_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__12643__C _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16074_ _16071_/A _16072_/Y _15902_/A _15905_/A vssd1 vssd1 vccd1 vccd1 _16075_/B
+ sky130_fd_sc_hd__o211ai_1
X_13286_ _13373_/B _13286_/B vssd1 vssd1 vccd1 vccd1 _13348_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13458__D _14218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15025_ _14816_/X _14819_/X _15023_/X _15024_/Y vssd1 vssd1 vccd1 vccd1 _15025_/X
+ sky130_fd_sc_hd__o211a_1
X_19902_ _19902_/A _19902_/B vssd1 vssd1 vccd1 vccd1 _19917_/A sky130_fd_sc_hd__xnor2_1
X_12237_ _12203_/X _12211_/Y _12234_/A _12241_/A vssd1 vssd1 vccd1 vccd1 _12238_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15954__C _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19833_ _19669_/B _19671_/B _19830_/X _19831_/Y vssd1 vssd1 vccd1 vccd1 _19833_/X
+ sky130_fd_sc_hd__a211o_1
X_12168_ _12168_/A _12168_/B _12168_/C vssd1 vssd1 vccd1 vccd1 _12168_/X sky130_fd_sc_hd__or3_1
XANTENNA__14818__A1 _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_16_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15673__D _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18009__A1 _18008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18009__B2 _18008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11119_ _10978_/Y hold61/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21713_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12829__B1 _11055_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19723__A _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19764_ _19742_/Y _19743_/X _19763_/C _19763_/D vssd1 vssd1 vccd1 vccd1 _19765_/B
+ sky130_fd_sc_hd__a2bb2o_1
X_16976_ _17096_/A _17124_/C _16974_/Y _16983_/A vssd1 vssd1 vccd1 vccd1 _16978_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_12099_ _12093_/A _12093_/B _12093_/C vssd1 vssd1 vccd1 vccd1 _12100_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_120_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18715_ _18712_/Y _18713_/X _18581_/D _18582_/B vssd1 vssd1 vccd1 vccd1 _18716_/B
+ sky130_fd_sc_hd__o211ai_1
X_15927_ _15927_/A _15927_/B vssd1 vssd1 vccd1 vccd1 _15938_/A sky130_fd_sc_hd__or2_1
X_19695_ _19695_/A _20419_/A _19695_/C _19695_/D vssd1 vssd1 vccd1 vccd1 _19695_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11706__D _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13771__A _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18646_ _19587_/B _19866_/D _19874_/B _19587_/A vssd1 vssd1 vccd1 vccd1 _18646_/X
+ sky130_fd_sc_hd__a22o_1
X_15858_ _15859_/A _15859_/B vssd1 vssd1 vccd1 vccd1 _15860_/A sky130_fd_sc_hd__nand2_1
XANTENNA__18058__B _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14809_ _14809_/A _14809_/B vssd1 vssd1 vccd1 vccd1 _14844_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_118_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18577_ _18693_/A _18576_/C _18576_/A vssd1 vssd1 vccd1 vccd1 _18678_/B sky130_fd_sc_hd__o21a_1
X_15789_ _15789_/A _15973_/B vssd1 vssd1 vccd1 vccd1 _15800_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13921__D _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17528_ _17526_/X _17528_/B vssd1 vssd1 vccd1 vccd1 _17529_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_129_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17459_ _17458_/A _17458_/B _17458_/C vssd1 vssd1 vccd1 vccd1 _17461_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20470_ _20470_/A _20470_/B vssd1 vssd1 vccd1 vccd1 _20471_/B sky130_fd_sc_hd__and2_1
XFILLER_0_14_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15210__B _15210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19129_ _19129_/A _19291_/A _19129_/C vssd1 vssd1 vccd1 vccd1 _19130_/C sky130_fd_sc_hd__or3_1
XFILLER_0_14_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout119_A _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20770__C _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_22071_ _22080_/CLK _22071_/D fanout639/X vssd1 vssd1 vccd1 vccd1 mstream_o[7] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_61_1030 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21022_ _21135_/A _21020_/X _20851_/Y _20856_/A vssd1 vssd1 vccd1 vccd1 _21022_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11335__A3 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13665__B _21364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout390_A _21771_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout488_A _21747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11740__B1 _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17759__B1 _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11616__D _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21924_ _21926_/CLK _21924_/D vssd1 vssd1 vccd1 vccd1 hold96/A sky130_fd_sc_hd__dfxtp_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21855_ _21923_/CLK _21855_/D vssd1 vssd1 vccd1 vccd1 hold206/A sky130_fd_sc_hd__dfxtp_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17303__D _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20806_ _20806_/A _20806_/B vssd1 vssd1 vccd1 vccd1 _20807_/B sky130_fd_sc_hd__nand2_1
X_21786_ _21788_/CLK _21786_/D vssd1 vssd1 vccd1 vccd1 _21786_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20737_ _20738_/B _20738_/A vssd1 vssd1 vccd1 vccd1 _20737_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_80_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17931__B1 _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11470_ _11469_/X _19951_/A _11470_/S vssd1 vssd1 vccd1 vccd1 _21828_/D sky130_fd_sc_hd__mux2_1
X_20668_ _21151_/A _20924_/A _21301_/A _21286_/A vssd1 vssd1 vccd1 vccd1 _20671_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11559__B1 _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15120__B _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12220__A1 _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12220__B2 _12242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13559__C _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20599_ _20600_/A _20600_/B vssd1 vssd1 vccd1 vccd1 _20601_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_150_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16498__B1 _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13140_ _13140_/A _13140_/B _13140_/C vssd1 vssd1 vccd1 vccd1 _13142_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13071_ _13072_/A _13072_/B _13072_/C vssd1 vssd1 vccd1 vccd1 _13071_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_143_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16232__A _16232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12022_ _12023_/A _12071_/A vssd1 vssd1 vccd1 vccd1 _12036_/B sky130_fd_sc_hd__nand2_1
XANTENNA__19987__A1 _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19987__B2 _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16589__D _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17998__B1 _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11731__B1 _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16830_ _16833_/A vssd1 vssd1 vccd1 vccd1 _16830_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13294__C _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11807__C _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout570 _21729_/Q vssd1 vssd1 vccd1 vccd1 _12403_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__20689__A _20689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout581 _12269_/D vssd1 vssd1 vccd1 vccd1 _12312_/A sky130_fd_sc_hd__buf_4
Xfanout592 _21724_/Q vssd1 vssd1 vccd1 vccd1 _11549_/A sky130_fd_sc_hd__buf_8
X_13973_ _13973_/A _13973_/B vssd1 vssd1 vccd1 vccd1 _14015_/A sky130_fd_sc_hd__or2_1
X_16761_ _17041_/A _17123_/C _17282_/A _16899_/B vssd1 vssd1 vccd1 vccd1 _16762_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19262__B _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13591__A _13875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18500_ _18500_/A _18500_/B _18500_/C vssd1 vssd1 vccd1 vccd1 _18503_/A sky130_fd_sc_hd__nand3_1
X_15712_ _15712_/A _15712_/B vssd1 vssd1 vccd1 vccd1 _15733_/A sky130_fd_sc_hd__xor2_2
X_12924_ _12924_/A _12924_/B _12924_/C vssd1 vssd1 vccd1 vccd1 _12924_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__17063__A _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16692_ _16691_/B _16691_/C _16691_/A vssd1 vssd1 vccd1 vccd1 _16694_/B sky130_fd_sc_hd__a21bo_1
X_19480_ _19476_/A _19476_/B _19471_/X vssd1 vssd1 vccd1 vccd1 _19635_/A sky130_fd_sc_hd__o21a_1
X_18431_ _20317_/D _19227_/C _19227_/D _19644_/A vssd1 vssd1 vccd1 vccd1 _18431_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__18962__A2 _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15643_ _16031_/A _15643_/B vssd1 vssd1 vccd1 vccd1 _15645_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_87_148 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12855_ _12855_/A _12855_/B vssd1 vssd1 vccd1 vccd1 _12869_/A sky130_fd_sc_hd__xor2_2
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11806_ _11805_/B _11805_/C _11805_/A vssd1 vssd1 vccd1 vccd1 _11806_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_56_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15574_ _15702_/D _15698_/B _15575_/C _15575_/D vssd1 vssd1 vccd1 vccd1 _15576_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_96_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18362_ _18363_/A _18363_/B _18363_/C vssd1 vssd1 vccd1 vccd1 _18362_/X sky130_fd_sc_hd__and3_1
XFILLER_0_28_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ _12785_/B _14384_/D _14391_/B _14248_/A vssd1 vssd1 vccd1 vccd1 _12787_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14525_ _14524_/A _14524_/B _14524_/C vssd1 vssd1 vccd1 vccd1 _14526_/C sky130_fd_sc_hd__a21o_1
X_17313_ _17313_/A _17313_/B vssd1 vssd1 vccd1 vccd1 _17315_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _11736_/B _11736_/C _11736_/A vssd1 vssd1 vccd1 vccd1 _11750_/B sky130_fd_sc_hd__a21o_1
XANTENNA__12357__D _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18293_ _18293_/A _18293_/B vssd1 vssd1 vccd1 vccd1 _18302_/A sky130_fd_sc_hd__or2_1
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14456_ _14936_/D _16084_/C _16084_/D _14306_/A vssd1 vssd1 vccd1 vccd1 _14456_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17244_ _17243_/A _17243_/B _17243_/C vssd1 vssd1 vccd1 vccd1 _17245_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_142_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11668_ _12316_/B _11668_/B vssd1 vssd1 vccd1 vccd1 _11670_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13407_ _13858_/A _14354_/C _14663_/D _21734_/Q vssd1 vssd1 vccd1 vccd1 _13409_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17175_ _17172_/Y _17173_/Y _17174_/X fanout3/X hold194/X vssd1 vssd1 vccd1 vccd1
+ _21886_/D sky130_fd_sc_hd__o32a_1
X_14387_ _14387_/A _14387_/B vssd1 vssd1 vccd1 vccd1 _14395_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18622__A _19092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11599_ _11596_/X _11599_/B vssd1 vssd1 vccd1 vccd1 _11874_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_113_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16126_ _16123_/Y _16124_/X _15991_/B _15992_/Y vssd1 vssd1 vccd1 vccd1 _16127_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_109_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13338_ _13338_/A _13338_/B _13338_/C vssd1 vssd1 vccd1 vccd1 _13338_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_24_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20590__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16057_ _16027_/A _16286_/B _16028_/A _15894_/A vssd1 vssd1 vccd1 vccd1 _16064_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_150_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13766__A _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15161__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17238__A _17557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13269_ _13864_/B _13867_/A _13269_/C _13269_/D vssd1 vssd1 vccd1 vccd1 _13416_/A
+ sky130_fd_sc_hd__and4_1
X_15008_ _14881_/B _14883_/B _15006_/X _15007_/Y vssd1 vssd1 vccd1 vccd1 _15012_/C
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__16499__D _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19816_ _19816_/A _19816_/B vssd1 vssd1 vccd1 vccd1 _19818_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16661__B1 _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19747_ _19866_/C _19746_/X _19745_/X vssd1 vssd1 vccd1 vccd1 _19749_/A sky130_fd_sc_hd__a21bo_1
X_16959_ _16956_/A _16956_/Y _16958_/X vssd1 vssd1 vccd1 vccd1 _16961_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_155_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19678_ _19678_/A _19678_/B vssd1 vssd1 vccd1 vccd1 _19679_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__15216__A1 _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14019__A2 _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18629_ _18630_/A _18630_/B vssd1 vssd1 vccd1 vccd1 _18629_/X sky130_fd_sc_hd__or2_1
XFILLER_0_149_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17123__D _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21640_ _21722_/CLK hold310/X fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[103]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21571_ mstream_o[34] _11048_/Y _21579_/S vssd1 vssd1 vccd1 vccd1 _22098_/D sky130_fd_sc_hd__mux2_1
XANTENNA_11 _11331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12845__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_22 _11339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout236_A _20991_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_33 _11412_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20522_ _20910_/A _21256_/B _20523_/C _20523_/D vssd1 vssd1 vccd1 vccd1 _20528_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA_44 hold247/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_55 hold275/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_66 hold274/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12564__B _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_77 hold277/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_88 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20453_ _20450_/X _20451_/Y _20302_/B _20302_/Y vssd1 vssd1 vccd1 vccd1 _20499_/B
+ sky130_fd_sc_hd__a211oi_4
XANTENNA_99 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout403_A _21769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13379__C _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22069__RESET_B fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20384_ _20245_/A _20428_/B _20254_/B _20252_/Y vssd1 vssd1 vccd1 vccd1 _20403_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15152__B1 _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22054_ _22063_/CLK _22054_/D vssd1 vssd1 vccd1 vccd1 hold286/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__16987__A _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21005_ _21005_/A _21005_/B _21005_/C vssd1 vssd1 vccd1 vccd1 _21005_/X sky130_fd_sc_hd__or3_2
XANTENNA__11627__C _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21633__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19197__A2 _19053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10970_ hold76/A hold100/A vssd1 vssd1 vccd1 vccd1 _10971_/B sky130_fd_sc_hd__nand2_1
XANTENNA_fanout51_A _11122_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21907_ _21939_/CLK _21907_/D vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__15115__B _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_12_clk_i _21806_/CLK vssd1 vssd1 vccd1 vccd1 _22049_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__19810__B _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13561__D _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11135__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12458__C _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17611__A _17854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12640_ _12528_/B _15768_/A _12639_/C _12639_/D vssd1 vssd1 vccd1 vccd1 _12641_/B
+ sky130_fd_sc_hd__a22o_1
X_21838_ _21845_/CLK _21838_/D vssd1 vssd1 vccd1 vccd1 _21838_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12441__A1 _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12571_ _12570_/A _12570_/B _12570_/C vssd1 vssd1 vccd1 vccd1 _12572_/C sky130_fd_sc_hd__a21o_1
X_21769_ _21789_/CLK _21769_/D vssd1 vssd1 vccd1 vccd1 _21769_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14310_ _16084_/D _14138_/X _14141_/A _14141_/B vssd1 vssd1 vccd1 vccd1 _14311_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_68_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11522_ _21723_/D t1y[24] t0x[24] _11223_/A vssd1 vssd1 vccd1 vccd1 _11522_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_136_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15290_ _15290_/A _15290_/B vssd1 vssd1 vccd1 vccd1 _15292_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12992__A2 _13269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_27_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21923_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14241_ _14713_/B _14557_/D _15234_/C _14713_/A vssd1 vssd1 vccd1 vccd1 _14241_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14194__A1 _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11453_ _21718_/Q t1y[1] t0x[1] _21724_/D vssd1 vssd1 vccd1 vccd1 _11453_/X sky130_fd_sc_hd__a22o_1
XANTENNA__19538__A _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13289__C _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20691__B _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14172_ _14173_/A _14173_/B vssd1 vssd1 vccd1 vccd1 _14172_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_1_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19257__B _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11384_ _11124_/A hold278/X fanout45/X hold210/X vssd1 vssd1 vccd1 vccd1 _11384_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13123_ _13975_/B _14018_/C _12982_/B _12980_/X vssd1 vssd1 vccd1 vccd1 _13124_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_132_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18980_ _18979_/B _18979_/C _18979_/A vssd1 vssd1 vccd1 vccd1 _18980_/X sky130_fd_sc_hd__o21a_1
XANTENNA__15694__A1 _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ _13054_/A _13054_/B _13054_/C vssd1 vssd1 vccd1 vccd1 _13056_/B sky130_fd_sc_hd__nand3_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17931_ _19123_/B _19262_/C _19414_/C _19123_/A vssd1 vssd1 vccd1 vccd1 _17932_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12005_ _12899_/B _12246_/D vssd1 vssd1 vccd1 vccd1 _12055_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17435__A2 _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17862_ _18873_/A _19227_/C _19227_/D _18849_/A vssd1 vssd1 vccd1 vccd1 _17863_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14249__A2 _21759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19601_ _19732_/A _19732_/B _19972_/C _21258_/B vssd1 vssd1 vccd1 vccd1 _19729_/A
+ sky130_fd_sc_hd__nand4_2
X_16813_ _16813_/A _17029_/B _17063_/C _17086_/C vssd1 vssd1 vccd1 vccd1 _16815_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13457__B1 _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17793_ _19123_/B _18789_/B _19262_/C _19123_/A vssd1 vssd1 vccd1 vccd1 _17794_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19532_ _19532_/A _19532_/B vssd1 vssd1 vccd1 vccd1 _19542_/A sky130_fd_sc_hd__xor2_1
X_16744_ _21830_/Q _17019_/C vssd1 vssd1 vccd1 vccd1 _16818_/A sky130_fd_sc_hd__nand2_1
X_13956_ _13956_/A _13956_/B _13956_/C vssd1 vssd1 vccd1 vccd1 _13958_/A sky130_fd_sc_hd__nor3_2
XFILLER_0_89_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17224__C _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12907_ _14712_/A _14712_/B _14386_/B vssd1 vssd1 vccd1 vccd1 _12907_/X sky130_fd_sc_hd__and3_1
X_19463_ _19464_/B _19464_/A vssd1 vssd1 vccd1 vccd1 _19463_/Y sky130_fd_sc_hd__nand2b_1
X_13887_ _13884_/Y _13885_/X _13757_/X _13795_/A vssd1 vssd1 vccd1 vccd1 _13887_/X
+ sky130_fd_sc_hd__a211o_1
X_16675_ _16676_/A _16676_/B _16676_/C vssd1 vssd1 vccd1 vccd1 _16675_/X sky130_fd_sc_hd__and3_1
XFILLER_0_33_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18414_ _18414_/A _18414_/B _18414_/C vssd1 vssd1 vccd1 vccd1 _18414_/X sky130_fd_sc_hd__and3_1
XFILLER_0_69_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15626_ _15626_/A _15626_/B vssd1 vssd1 vccd1 vccd1 _15626_/Y sky130_fd_sc_hd__xnor2_2
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12838_ _13083_/A _12838_/B vssd1 vssd1 vccd1 vccd1 _12938_/A sky130_fd_sc_hd__and2_1
XFILLER_0_115_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19394_ _19393_/B _19543_/B _19393_/A vssd1 vssd1 vccd1 vccd1 _19395_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_57_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21043__A _21267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18336__B _19732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18345_ _19438_/A _19438_/B _19262_/C _19414_/C vssd1 vssd1 vccd1 vccd1 _18345_/X
+ sky130_fd_sc_hd__and4_1
X_15557_ _15558_/A _15558_/B vssd1 vssd1 vccd1 vccd1 _15682_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_139_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_663 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12769_ _12765_/X _12766_/Y _12648_/X _12650_/X vssd1 vssd1 vccd1 vccd1 _12803_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14508_ _14508_/A _15022_/B _14508_/C _14508_/D vssd1 vssd1 vccd1 vccd1 _14508_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_12_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15488_ _15351_/A _15351_/B _15349_/X vssd1 vssd1 vccd1 vccd1 _15490_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18276_ _18277_/A _18277_/B vssd1 vssd1 vccd1 vccd1 _18398_/B sky130_fd_sc_hd__and2_1
XFILLER_0_72_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17227_ _17227_/A _17227_/B vssd1 vssd1 vccd1 vccd1 _17229_/B sky130_fd_sc_hd__xnor2_2
X_14439_ _14439_/A _14439_/B vssd1 vssd1 vccd1 vccd1 _14442_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17894__C _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12196__B1 _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17158_ _17158_/A _17158_/B vssd1 vssd1 vccd1 vccd1 _17159_/D sky130_fd_sc_hd__nand2_1
X_16109_ _16110_/B _16110_/A vssd1 vssd1 vccd1 vccd1 _16109_/Y sky130_fd_sc_hd__nand2b_1
X_17089_ _17089_/A _17089_/B _17089_/C vssd1 vssd1 vccd1 vccd1 _17089_/X sky130_fd_sc_hd__or3_1
XANTENNA__13927__C _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20106__B _21832_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18623__A1 _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16600__A _18058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout186_A _21824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12559__B _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14477__D _14635_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout353_A _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13381__D _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14948__B1 _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14774__B _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21623_ _21939_/CLK _21623_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[86] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_75_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout520_A _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout618_A _21717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_814 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21554_ mstream_o[17] hold32/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22081_/D sky130_fd_sc_hd__mux2_1
XANTENNA__20792__A _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10985__A1 _10984_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20505_ _20357_/Y _20359_/Y _20503_/Y _20504_/X vssd1 vssd1 vccd1 vccd1 _20639_/A
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__15912__A2 _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14790__A _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21485_ hold201/X sstream_i[62] _21507_/S vssd1 vssd1 vccd1 vccd1 _22012_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_31_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12187__B1 _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12726__A2 _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20436_ _20436_/A _20436_/B vssd1 vssd1 vccd1 vccd1 _20438_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21806__CLK _21806_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17665__A2 _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11919__A _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20367_ _20367_/A _20367_/B vssd1 vssd1 vccd1 vccd1 _20370_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13837__C _14477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout99_A _19060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22106_ _22106_/CLK _22106_/D _11089_/A vssd1 vssd1 vccd1 vccd1 mstream_o[42] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20298_ _20449_/B _20296_/X _20115_/X _20118_/Y vssd1 vssd1 vccd1 vccd1 _20299_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_101_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22037_ _22049_/CLK _22037_/D vssd1 vssd1 vccd1 vccd1 hold233/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13151__A2 _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17606__A _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19093__A _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14949__B _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13810_ _13656_/B _13656_/Y _13818_/B _13809_/Y vssd1 vssd1 vccd1 vccd1 _13962_/A
+ sky130_fd_sc_hd__o211ai_4
X_14790_ _15153_/B _15978_/B _14790_/C _14946_/A vssd1 vssd1 vccd1 vccd1 _14946_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__15161__A1_N _21734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13741_ _14365_/A _14384_/A _14212_/B _14367_/A vssd1 vssd1 vccd1 vccd1 _13744_/A
+ sky130_fd_sc_hd__a22o_1
X_10953_ _10945_/A _10945_/B _10945_/C _10950_/A vssd1 vssd1 vccd1 vccd1 _10953_/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__12662__A1 _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13672_ _16399_/B _13671_/X _13670_/X vssd1 vssd1 vccd1 vccd1 _13674_/A sky130_fd_sc_hd__a21bo_1
X_16460_ _17041_/A _16899_/B _17013_/D vssd1 vssd1 vccd1 vccd1 _16460_/X sky130_fd_sc_hd__and3_1
X_10884_ _10885_/A _10885_/B _10885_/C vssd1 vssd1 vccd1 vccd1 _10886_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20690__A2_N _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15411_ _15808_/C _16040_/C _15409_/Y _15547_/A vssd1 vssd1 vccd1 vccd1 _15413_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_66_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12623_ _12530_/C _12532_/A _12732_/B _12622_/X vssd1 vssd1 vccd1 vccd1 _12743_/A
+ sky130_fd_sc_hd__a211o_1
X_16391_ _16391_/A _16391_/B vssd1 vssd1 vccd1 vccd1 _16392_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_155_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15342_ _15342_/A _15342_/B vssd1 vssd1 vccd1 vccd1 _15345_/A sky130_fd_sc_hd__xnor2_4
X_18130_ _18849_/A _18732_/C _19221_/C _18849_/B vssd1 vssd1 vccd1 vccd1 _18130_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12554_ _12554_/A _12554_/B vssd1 vssd1 vccd1 vccd1 _12556_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__16156__A2 _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11505_ _11224_/A t2x[18] v1z[18] fanout21/X _11504_/X vssd1 vssd1 vccd1 vccd1 _11505_/X
+ sky130_fd_sc_hd__a221o_1
X_15273_ _15931_/B _16040_/C _16396_/A _15931_/A vssd1 vssd1 vccd1 vccd1 _15273_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_123_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18061_ _18061_/A _18061_/B vssd1 vssd1 vccd1 vccd1 _18062_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_145_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12485_ _12484_/B _12484_/C _12484_/A vssd1 vssd1 vccd1 vccd1 _12485_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14224_ _14224_/A _14224_/B _14224_/C vssd1 vssd1 vccd1 vccd1 _14226_/B sky130_fd_sc_hd__nand3_2
XANTENNA__13914__A1 _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17012_ _16971_/A _16971_/C _16971_/B vssd1 vssd1 vccd1 vccd1 _17018_/B sky130_fd_sc_hd__a21o_1
X_11436_ hold238/A fanout28/X _11435_/X vssd1 vssd1 vccd1 vccd1 _11436_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_145_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16404__B _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14155_ _15159_/D _14936_/D _14155_/C _14155_/D vssd1 vssd1 vccd1 vccd1 _14157_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_145_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17656__A2 _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ hold165/X fanout29/X _11366_/X vssd1 vssd1 vccd1 vccd1 _11367_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_104_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18900__A _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13106_ _13104_/A _13104_/B _13104_/C vssd1 vssd1 vccd1 vccd1 _13244_/B sky130_fd_sc_hd__a21oi_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14086_ _14086_/A _14086_/B vssd1 vssd1 vccd1 vccd1 _14095_/A sky130_fd_sc_hd__xor2_2
X_18963_ _19123_/A _20247_/D _20721_/C vssd1 vssd1 vccd1 vccd1 _18964_/C sky130_fd_sc_hd__and3_1
XFILLER_0_81_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11298_ _11224_/A t1x[18] v2z[18] _11507_/B2 _11297_/X vssd1 vssd1 vccd1 vccd1 _11298_/X
+ sky130_fd_sc_hd__a221o_2
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ _14367_/A _15217_/A _13169_/A _13036_/D vssd1 vssd1 vccd1 vccd1 _13038_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17914_ _19439_/A _17915_/D _17787_/X _17788_/X _17670_/B vssd1 vssd1 vccd1 vccd1
+ _17919_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18894_ _20178_/D _18894_/B _18894_/C _18894_/D vssd1 vssd1 vccd1 vccd1 _18895_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__20412__A1 _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17845_ _18121_/A _17845_/B vssd1 vssd1 vccd1 vccd1 _17847_/C sky130_fd_sc_hd__or2_1
XANTENNA__11564__A _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17776_ _17776_/A _17776_/B vssd1 vssd1 vccd1 vccd1 _17810_/A sky130_fd_sc_hd__nand2_1
X_14988_ _14865_/B _14865_/C _14865_/D _14851_/X vssd1 vssd1 vccd1 vccd1 _14990_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_152_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18908__A2 _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19515_ _19514_/B _19514_/C _19503_/Y vssd1 vssd1 vccd1 vccd1 _19515_/Y sky130_fd_sc_hd__a21boi_1
X_16727_ _16727_/A _16727_/B _16727_/C vssd1 vssd1 vccd1 vccd1 _16800_/A sky130_fd_sc_hd__nand3_1
X_13939_ _13939_/A _13939_/B _13939_/C vssd1 vssd1 vccd1 vccd1 _13939_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_89_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19446_ _19292_/A _19292_/B _19847_/A vssd1 vssd1 vccd1 vccd1 _19448_/B sky130_fd_sc_hd__a21oi_2
X_16658_ _17178_/B _16657_/B _16657_/C _16657_/D vssd1 vssd1 vccd1 vccd1 _16658_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15609_ _15693_/B _15606_/Y _15422_/X _15426_/C vssd1 vssd1 vccd1 vccd1 _15609_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19377_ _19535_/B _20416_/A _20416_/B _19686_/A vssd1 vssd1 vccd1 vccd1 _19382_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16589_ _16590_/A _16588_/Y _16870_/A _17526_/B vssd1 vssd1 vccd1 vccd1 _16628_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11503__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18328_ _18328_/A _18328_/B _18328_/C vssd1 vssd1 vccd1 vccd1 _18328_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_45_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17895__A2 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18259_ _18259_/A _18402_/B vssd1 vssd1 vccd1 vccd1 _18261_/B sky130_fd_sc_hd__or2_1
XFILLER_0_4_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_71_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21270_ _21174_/A _21174_/B _21270_/S vssd1 vssd1 vccd1 vccd1 _21271_/B sky130_fd_sc_hd__mux2_1
XFILLER_0_13_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11739__A _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20221_ _20222_/A _20222_/B _20220_/Y vssd1 vssd1 vccd1 vccd1 _20221_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_130_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19906__A _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20100__B1 _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout101_A _21842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17129__C _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11392__A1 _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_1128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20152_ _20153_/A _20153_/B vssd1 vssd1 vccd1 vccd1 _20294_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_110_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13133__A2 _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20083_ _20372_/A _20083_/B vssd1 vssd1 vccd1 vccd1 _21393_/B sky130_fd_sc_hd__xnor2_2
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16607__B1 _17557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13673__B _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17145__B _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11695__A2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15591__D _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout470_A _15091_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout568_A _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1068 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14633__A2 _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21382__S _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20985_ _20985_/A _20985_/B vssd1 vssd1 vccd1 vccd1 _20996_/A sky130_fd_sc_hd__or2_1
XFILLER_0_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16386__A2 _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19324__A2 _19322_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11413__S _11446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21606_ _21934_/CLK _21606_/D _11041_/A vssd1 vssd1 vccd1 vccd1 mstream_o[69] sky130_fd_sc_hd__dfrtp_4
XANTENNA_hold313_A hold313/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout14_A wire16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11080__A0 _10941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21537_ mstream_o[0] hold13/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22064_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_51_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1028 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12270_ _12217_/B _12268_/X _12269_/X vssd1 vssd1 vccd1 vccd1 _12271_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_105_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21468_ hold170/X sstream_i[45] _21481_/S vssd1 vssd1 vccd1 vccd1 _21995_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_121_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15766__D _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11221_ hold202/X fanout22/X _11220_/X vssd1 vssd1 vccd1 vccd1 _11221_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_142_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17638__A2 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20419_ _20419_/A _21286_/A _20419_/C _20419_/D vssd1 vssd1 vccd1 vccd1 _20552_/B
+ sky130_fd_sc_hd__and4_1
X_21399_ _21420_/S _21399_/B vssd1 vssd1 vccd1 vccd1 _21399_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11383__A1 _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15649__A1 _15907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11152_ hold183/X fanout23/X _11151_/X vssd1 vssd1 vccd1 vccd1 _11152_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_102_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13864__A _21738_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15960_ _15960_/A _15960_/B vssd1 vssd1 vccd1 vccd1 _15965_/A sky130_fd_sc_hd__xnor2_2
X_11083_ _10959_/Y hold3/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21678_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_41_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21198__A2 _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14911_ _14911_/A _14911_/B vssd1 vssd1 vccd1 vccd1 _14913_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17055__B _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15891_ hold208/X _15890_/X fanout2/X vssd1 vssd1 vccd1 vccd1 _21880_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12883__A1 _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12883__B2 _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17630_ _17630_/A _17630_/B _17630_/C vssd1 vssd1 vccd1 vccd1 _17630_/Y sky130_fd_sc_hd__nor3_4
X_14842_ _14709_/A _14710_/Y _14840_/Y _14841_/X vssd1 vssd1 vccd1 vccd1 _14844_/B
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__19012__A1 _19493_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17561_ _17450_/A _17450_/C _17450_/B vssd1 vssd1 vccd1 vccd1 _17562_/C sky130_fd_sc_hd__a21bo_1
X_14773_ _14773_/A _14773_/B vssd1 vssd1 vccd1 vccd1 _14778_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__19012__B2 _19337_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11985_ _12458_/A _12751_/B _12637_/B _12269_/B vssd1 vssd1 vccd1 vccd1 _11986_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14695__A _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18167__A _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19300_ _19300_/A _19300_/B vssd1 vssd1 vccd1 vccd1 _19303_/A sky130_fd_sc_hd__xnor2_2
X_16512_ _16989_/C _17619_/A _16512_/C _16564_/A vssd1 vssd1 vccd1 vccd1 _16564_/B
+ sky130_fd_sc_hd__nand4_1
X_13724_ _14027_/A _16286_/A _13724_/C _13724_/D vssd1 vssd1 vccd1 vccd1 _13724_/X
+ sky130_fd_sc_hd__and4_1
X_10936_ hold79/A hold101/A vssd1 vssd1 vccd1 vccd1 _10938_/A sky130_fd_sc_hd__or2_1
XFILLER_0_85_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21305__B _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17492_ _17490_/A _20797_/A _21258_/A _21792_/Q vssd1 vssd1 vccd1 vccd1 _17493_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17502__C _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21370__A2 _13967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18771__B1 _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14388__A1 _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19231_ _19056_/X _19059_/X _19228_/X _19230_/Y vssd1 vssd1 vccd1 vccd1 _19231_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15303__B _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16443_ _16444_/A _16442_/Y _16870_/A _16917_/C vssd1 vssd1 vccd1 vccd1 _16697_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_39_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14388__B2 _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10867_ _10873_/B _10867_/B vssd1 vssd1 vccd1 vccd1 _10867_/X sky130_fd_sc_hd__and2_2
X_13655_ _13652_/Y _13653_/X _13500_/C _13501_/X vssd1 vssd1 vccd1 vccd1 _13656_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_156_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19162_ _19162_/A _19162_/B vssd1 vssd1 vccd1 vccd1 _19163_/B sky130_fd_sc_hd__nand2_1
X_12606_ _12606_/A _12606_/B vssd1 vssd1 vccd1 vccd1 _12701_/A sky130_fd_sc_hd__xnor2_1
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16374_ _16374_/A _16374_/B vssd1 vssd1 vccd1 vccd1 _16376_/A sky130_fd_sc_hd__or2_1
X_13586_ _13428_/A _13428_/Y _13583_/X _13584_/Y vssd1 vssd1 vccd1 vccd1 _13586_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_155_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10798_ _20721_/C vssd1 vssd1 vccd1 vccd1 _10798_/Y sky130_fd_sc_hd__inv_2
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11071__A0 _10874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20863__C _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18113_ _18703_/A _19201_/B _18253_/A _18111_/Y vssd1 vssd1 vccd1 vccd1 _18114_/C
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__15337__B1 _15336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15325_ _15326_/A _15326_/B vssd1 vssd1 vccd1 vccd1 _15325_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_82_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12537_ _12537_/A _12537_/B vssd1 vssd1 vccd1 vccd1 _12540_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_81_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19093_ _20650_/A _19906_/C vssd1 vssd1 vccd1 vccd1 _19095_/C sky130_fd_sc_hd__and2_1
XFILLER_0_53_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21040__B _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18044_ _18044_/A _18044_/B _18044_/C vssd1 vssd1 vccd1 vccd1 _18046_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_2_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15256_ _16084_/A _16196_/A _15653_/C _15911_/C vssd1 vssd1 vccd1 vccd1 _15451_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_48_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12468_ _12468_/A _12468_/B _12468_/C vssd1 vssd1 vccd1 vccd1 _12471_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_151_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14207_ _14207_/A _14207_/B vssd1 vssd1 vccd1 vccd1 _14208_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_112_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11419_ _11418_/X _20270_/C _11470_/S vssd1 vssd1 vccd1 vccd1 _21811_/D sky130_fd_sc_hd__mux2_1
X_15187_ _15046_/Y _15050_/C _15296_/B _15186_/X vssd1 vssd1 vccd1 vccd1 _15346_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_105_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12399_ _12399_/A _12605_/A vssd1 vssd1 vccd1 vccd1 _12414_/A sky130_fd_sc_hd__and2_1
XFILLER_0_111_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11374__A1 _16743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14138_ _14138_/A _14463_/D _16084_/C vssd1 vssd1 vccd1 vccd1 _14138_/X sky130_fd_sc_hd__and3_1
XFILLER_0_1_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19995_ _20863_/C _20419_/A _19995_/C _20138_/A vssd1 vssd1 vccd1 vccd1 _20138_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_10_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14069_ _14209_/B _14068_/C _14068_/A vssd1 vssd1 vccd1 vccd1 _14070_/C sky130_fd_sc_hd__a21o_1
X_18946_ _18946_/A _18946_/B vssd1 vssd1 vccd1 vccd1 _18979_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18877_ _18876_/B _18876_/C _18876_/A vssd1 vssd1 vccd1 vccd1 _18878_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11677__A2 _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17828_ _17828_/A _17828_/B vssd1 vssd1 vccd1 vccd1 _17837_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19003__B2 _11550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17759_ _19664_/B _18767_/B _18616_/D _18008_/A vssd1 vssd1 vccd1 vccd1 _17759_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20770_ hold124/X _20770_/B _21142_/A vssd1 vssd1 vccd1 vccd1 _20770_/X sky130_fd_sc_hd__and3_1
XFILLER_0_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout17 fanout19/X vssd1 vssd1 vccd1 vccd1 fanout17/X sky130_fd_sc_hd__buf_4
XFILLER_0_58_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19429_ _17324_/D _20242_/C _20242_/D _19430_/A vssd1 vssd1 vccd1 vccd1 _19432_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout28 fanout29/X vssd1 vssd1 vccd1 vccd1 fanout28/X sky130_fd_sc_hd__buf_4
XFILLER_0_119_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout39 fanout40/X vssd1 vssd1 vccd1 vccd1 _21381_/B sky130_fd_sc_hd__buf_4
XFILLER_0_45_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout149_A _21832_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_249 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11062__A0 _11061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout316_A _17854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21322_ _21322_/A _21322_/B vssd1 vssd1 vccd1 vccd1 _21323_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13976__A2_N _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19636__A _19636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21253_ _21246_/A _21253_/B vssd1 vssd1 vccd1 vccd1 _21253_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_102_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11365__A1 _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20204_ _20205_/A _20205_/B vssd1 vssd1 vccd1 vccd1 _20204_/X sky130_fd_sc_hd__or2_1
X_21184_ _21185_/A _21185_/B vssd1 vssd1 vccd1 vccd1 _21186_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_111_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20135_ _21291_/A _20419_/A _20136_/C _20136_/D vssd1 vssd1 vccd1 vccd1 _20139_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__14499__B _14659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20066_ _20066_/A _20066_/B vssd1 vssd1 vccd1 vccd1 _20069_/A sky130_fd_sc_hd__xnor2_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19802__C _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_304 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_315 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_326 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_337 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19545__A2 _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11770_ _11770_/A _11770_/B vssd1 vssd1 vccd1 vccd1 _11772_/C sky130_fd_sc_hd__nor2_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20968_ _20838_/B _21291_/B _20969_/C _20969_/D vssd1 vssd1 vccd1 vccd1 _20970_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20560__B1 _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20899_ _20906_/A vssd1 vssd1 vccd1 vccd1 _20899_/Y sky130_fd_sc_hd__inv_2
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15031__A2 _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13440_ _14367_/A _15763_/A vssd1 vssd1 vccd1 vccd1 _13444_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17308__A1 _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17308__B2 _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13593__A2 _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13371_ hold315/X _13370_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _21863_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_36_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15110_ _15012_/B _15011_/Y _15107_/Y _15250_/B vssd1 vssd1 vccd1 vccd1 _15147_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_23_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12322_ _12401_/A _12322_/B _12403_/A _15768_/A vssd1 vssd1 vccd1 vccd1 _12401_/B
+ sky130_fd_sc_hd__and4b_1
X_16090_ _16091_/A _16091_/B vssd1 vssd1 vccd1 vccd1 _16207_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15041_ _15044_/B vssd1 vssd1 vccd1 vccd1 _15041_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_32_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14542__A1 _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12253_ _12217_/X _12244_/Y _12245_/X _12248_/X vssd1 vssd1 vccd1 vccd1 _12254_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_121_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19546__A _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__A1 _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11204_ _14234_/C _11203_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21751_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_31_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18284__A2 _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12184_ _12183_/B _12183_/C _12183_/A vssd1 vssd1 vccd1 vccd1 _12185_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_102_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18800_ _19123_/B _20249_/B _20247_/C _19123_/A vssd1 vssd1 vccd1 vccd1 _18802_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13594__A _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17492__B1 _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11135_ _12246_/D _11134_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21728_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19780_ _19942_/A _19780_/B vssd1 vssd1 vccd1 vccd1 _19782_/B sky130_fd_sc_hd__and2_1
X_16992_ _16992_/A _16992_/B vssd1 vssd1 vccd1 vccd1 _16994_/B sky130_fd_sc_hd__xor2_1
X_18731_ _19644_/A _18732_/C _18894_/B _19487_/A vssd1 vssd1 vccd1 vccd1 _18733_/A
+ sky130_fd_sc_hd__a22oi_1
X_15943_ _16078_/A _15941_/C _15941_/A vssd1 vssd1 vccd1 vccd1 _15943_/Y sky130_fd_sc_hd__a21oi_2
X_11066_ _11066_/A _11066_/B vssd1 vssd1 vccd1 vccd1 _11066_/Y sky130_fd_sc_hd__nor2_4
XANTENNA__18036__A2 _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16047__A1 _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19281__A _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18662_ _18661_/A _18661_/B _18661_/C vssd1 vssd1 vccd1 vccd1 _18664_/C sky130_fd_sc_hd__a21o_1
X_15874_ _15874_/A _15874_/B _15874_/C _15874_/D vssd1 vssd1 vccd1 vccd1 _15874_/X
+ sky130_fd_sc_hd__or4_2
X_17613_ _17732_/B _17613_/B vssd1 vssd1 vccd1 vccd1 _17616_/A sky130_fd_sc_hd__or2_2
X_14825_ _14825_/A _14825_/B vssd1 vssd1 vccd1 vccd1 _14833_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_153_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18593_ _18720_/B _18593_/B vssd1 vssd1 vccd1 vccd1 _18608_/A sky130_fd_sc_hd__and2_1
XTAP_3860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_116_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19536__A2 _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17544_ _20583_/A _19951_/A _19951_/B _19892_/A vssd1 vssd1 vccd1 vccd1 _17544_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14756_ _14758_/A _14758_/B vssd1 vssd1 vccd1 vccd1 _14756_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11968_ _11969_/B _11969_/C _11969_/A vssd1 vssd1 vccd1 vccd1 _11979_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11292__A0 _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13707_ _14306_/A _13997_/C _13707_/C _13707_/D vssd1 vssd1 vccd1 vccd1 _13708_/B
+ sky130_fd_sc_hd__nand4_1
X_10919_ _10919_/A _10919_/B vssd1 vssd1 vccd1 vccd1 _10919_/X sky130_fd_sc_hd__xor2_4
X_17475_ _17475_/A _17475_/B vssd1 vssd1 vccd1 vccd1 _17478_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_58_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14687_ _14809_/B _14685_/X _14549_/Y _14553_/A vssd1 vssd1 vccd1 vccd1 _14688_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_6_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11899_ _11899_/A _11899_/B _11899_/C vssd1 vssd1 vccd1 vccd1 _11900_/B sky130_fd_sc_hd__and3_1
XFILLER_0_15_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_12_clk_i_A _21806_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19214_ _19214_/A _19214_/B vssd1 vssd1 vccd1 vccd1 _19216_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16426_ _16291_/A _16291_/B _16294_/A vssd1 vssd1 vccd1 vccd1 _16430_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13638_ _13638_/A _13638_/B _13638_/C vssd1 vssd1 vccd1 vccd1 _13638_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__13033__A1 _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13033__B2 _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11044__A0 _11043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19145_ _18981_/X _18983_/X _19143_/X _19144_/Y vssd1 vssd1 vccd1 vccd1 _19145_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16357_ _16250_/A _16250_/B _16248_/A vssd1 vssd1 vccd1 vccd1 _16359_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_27_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16145__A fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13569_ _13569_/A _13569_/B vssd1 vssd1 vccd1 vccd1 _13578_/A sky130_fd_sc_hd__or2_1
XANTENNA__12673__A _12784_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15308_ _21734_/Q _15838_/B _16314_/D _21735_/Q vssd1 vssd1 vccd1 vccd1 _15449_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_81_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19076_ _19076_/A _19076_/B _19076_/C vssd1 vssd1 vccd1 vccd1 _19078_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_70_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16288_ _16287_/B _16287_/C _16287_/A vssd1 vssd1 vccd1 vccd1 _16289_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_2_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12392__B _12392_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18027_ _17921_/A _17921_/C _17921_/B vssd1 vssd1 vccd1 vccd1 _18042_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_48_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15239_ _15240_/A _15240_/B vssd1 vssd1 vccd1 vccd1 _15384_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11347__A1 _21407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout207 _21816_/Q vssd1 vssd1 vccd1 vccd1 _21046_/B sky130_fd_sc_hd__buf_4
XFILLER_0_10_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout218 hold323/X vssd1 vssd1 vccd1 vccd1 _21040_/A sky130_fd_sc_hd__buf_4
Xfanout229 _20273_/A vssd1 vssd1 vccd1 vccd1 _19703_/C sky130_fd_sc_hd__clkbuf_4
X_19978_ _20098_/A _19977_/C _19977_/A vssd1 vssd1 vccd1 vccd1 _19979_/C sky130_fd_sc_hd__a21o_1
XANTENNA__14297__B1 _10881_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18929_ _21833_/Q _18929_/B _19546_/D vssd1 vssd1 vccd1 vccd1 _18929_/X sky130_fd_sc_hd__and3_1
XFILLER_0_66_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11228__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21940_ _21942_/CLK _21940_/D vssd1 vssd1 vccd1 vccd1 hold167/A sky130_fd_sc_hd__dfxtp_1
X_21871_ _21934_/CLK _21871_/D vssd1 vssd1 vccd1 vccd1 hold216/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20130__A _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout266_A _18030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20822_ _20824_/B vssd1 vssd1 vccd1 vccd1 _20822_/Y sky130_fd_sc_hd__inv_2
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11283__B1 _11282_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15549__B1 _14698_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20753_ _20753_/A vssd1 vssd1 vccd1 vccd1 _20755_/C sky130_fd_sc_hd__inv_2
XFILLER_0_119_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout433_A _14712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_465 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20684_ _20872_/B _20684_/B vssd1 vssd1 vccd1 vccd1 _20699_/A sky130_fd_sc_hd__and2_1
XFILLER_0_134_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16761__A2 _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21098__A1 _21311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21098__B2 _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11586__A1 _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11586__B2 _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16513__A2 _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21305_ _21305_/A _21305_/B vssd1 vssd1 vccd1 vccd1 _21307_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12535__B1 _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21236_ _21236_/A _21236_/B _21236_/C vssd1 vssd1 vccd1 vccd1 _21237_/B sky130_fd_sc_hd__or3_1
XFILLER_0_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold250 hold250/A vssd1 vssd1 vccd1 vccd1 hold250/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold261 hold261/A vssd1 vssd1 vccd1 vccd1 hold261/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold272 hold272/A vssd1 vssd1 vccd1 vccd1 hold272/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 hold283/A vssd1 vssd1 vccd1 vccd1 hold283/X sky130_fd_sc_hd__buf_4
Xhold294 hold294/A vssd1 vssd1 vccd1 vccd1 hold294/X sky130_fd_sc_hd__dlygate4sd3_1
X_21167_ _21056_/A _21169_/A _21056_/B vssd1 vssd1 vccd1 vccd1 _21168_/A sky130_fd_sc_hd__o21ai_1
XANTENNA_fanout81_A _19030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14827__A2 _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20118_ _20118_/A vssd1 vssd1 vccd1 vccd1 _20118_/Y sky130_fd_sc_hd__inv_2
X_21098_ _21311_/A _21283_/B _21305_/B _21286_/A vssd1 vssd1 vccd1 vccd1 _21102_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11138__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20049_ _20049_/A _20049_/B _20188_/B vssd1 vssd1 vccd1 vccd1 _20186_/A sky130_fd_sc_hd__or3_1
X_12940_ _12813_/B _12812_/Y _12938_/Y _12939_/X vssd1 vssd1 vccd1 vccd1 _12961_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_3112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11510__A1 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18429__B _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ _12765_/X _12768_/Y _12869_/X _12870_/Y vssd1 vssd1 vccd1 vccd1 _12971_/A
+ sky130_fd_sc_hd__a211o_2
XANTENNA_101 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_112 sstream_i[65] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14610_ _14469_/A _14469_/B _14472_/A vssd1 vssd1 vccd1 vccd1 _14755_/A sky130_fd_sc_hd__a21o_2
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_123 v0z[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18148__C _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_134 v1z[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11822_ _11823_/A _11823_/B _11823_/C vssd1 vssd1 vccd1 vccd1 _11822_/X sky130_fd_sc_hd__and3_1
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15590_ _15593_/D vssd1 vssd1 vccd1 vccd1 _15590_/Y sky130_fd_sc_hd__inv_2
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17052__C _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_145 v1z[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_156 v2z[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_167 v2z[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14541_ _14543_/D vssd1 vssd1 vccd1 vccd1 _14541_/Y sky130_fd_sc_hd__inv_2
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_178 v2z[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11753_ _11753_/A _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11753_/Y sky130_fd_sc_hd__nand3_2
XANTENNA_189 hold247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13015__A1 _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17260_ _17260_/A _17363_/A _17260_/C vssd1 vssd1 vccd1 vccd1 _17363_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_154_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15788__B _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14472_ _14472_/A _14472_/B vssd1 vssd1 vccd1 vccd1 _14492_/A sky130_fd_sc_hd__or2_2
XFILLER_0_3_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11684_ _11705_/B _11682_/C _11682_/A vssd1 vssd1 vccd1 vccd1 _11685_/C sky130_fd_sc_hd__a21o_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16211_ _16211_/A _16211_/B vssd1 vssd1 vccd1 vccd1 _16232_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_153_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13589__A _21742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13423_ _13580_/A _13423_/B vssd1 vssd1 vccd1 vccd1 _13425_/B sky130_fd_sc_hd__and2_1
XFILLER_0_64_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17191_ _17191_/A _17191_/B vssd1 vssd1 vccd1 vccd1 _17194_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_52_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12493__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16142_ _16142_/A _16142_/B vssd1 vssd1 vccd1 vccd1 _16144_/A sky130_fd_sc_hd__nor2_1
X_13354_ _13353_/B _13353_/C _13353_/A vssd1 vssd1 vccd1 vccd1 _13354_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15300__C _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12305_ _12306_/A _12305_/B _12304_/B vssd1 vssd1 vccd1 vccd1 _12305_/X sky130_fd_sc_hd__or3b_1
XANTENNA__14515__A1 _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12643__D _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16073_ _15902_/A _15905_/A _16071_/A _16072_/Y vssd1 vssd1 vccd1 vccd1 _16075_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__14515__B2 _16173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13285_ _13373_/A _13283_/Y _13139_/X _13142_/X vssd1 vssd1 vccd1 vccd1 _13286_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11329__B2 _11089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15024_ _15024_/A _15024_/B _15024_/C vssd1 vssd1 vccd1 vccd1 _15024_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_121_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12236_ _12234_/A _12241_/A _12203_/X _12211_/Y vssd1 vssd1 vccd1 vccd1 _12238_/B
+ sky130_fd_sc_hd__o211ai_1
X_19901_ _19899_/X _19901_/B vssd1 vssd1 vccd1 vccd1 _19902_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__15954__D _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19832_ _19669_/B _19671_/B _19830_/X _19831_/Y vssd1 vssd1 vccd1 vccd1 _19832_/Y
+ sky130_fd_sc_hd__a211oi_1
X_12167_ _12168_/A _12168_/B _12168_/C vssd1 vssd1 vccd1 vccd1 _12167_/Y sky130_fd_sc_hd__nor3_1
X_11118_ _10972_/Y hold5/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21712_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18009__A2 _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11556__B _12242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19763_ _19742_/Y _19743_/X _19763_/C _19763_/D vssd1 vssd1 vccd1 vccd1 _19763_/X
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__12829__A1 _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16975_ _17144_/A _17129_/B _17013_/D _17019_/C vssd1 vssd1 vccd1 vccd1 _16983_/A
+ sky130_fd_sc_hd__and4_1
X_12098_ _12098_/A _12098_/B vssd1 vssd1 vccd1 vccd1 _12100_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__12829__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18714_ _18581_/D _18582_/B _18712_/Y _18713_/X vssd1 vssd1 vccd1 vccd1 _18716_/A
+ sky130_fd_sc_hd__a211o_1
X_15926_ _16114_/B _15926_/B vssd1 vssd1 vccd1 vccd1 _15941_/A sky130_fd_sc_hd__and2_1
X_11049_ _11048_/Y hold143/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21654_/D sky130_fd_sc_hd__mux2_1
X_19694_ _19695_/A _20419_/A _19695_/C _19695_/D vssd1 vssd1 vccd1 vccd1 _19694_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__11501__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13771__B _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21046__A _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18645_ _19439_/A _19414_/C vssd1 vssd1 vccd1 vccd1 _18649_/A sky130_fd_sc_hd__nand2_1
X_15857_ _15857_/A _15857_/B vssd1 vssd1 vccd1 vccd1 _15859_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14808_ _14808_/A _14808_/B vssd1 vssd1 vccd1 vccd1 _14897_/A sky130_fd_sc_hd__xnor2_1
X_18576_ _18576_/A _18693_/A _18576_/C vssd1 vssd1 vccd1 vccd1 _18693_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_52_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15788_ _16409_/A _15788_/B _15788_/C _15973_/A vssd1 vssd1 vccd1 vccd1 _15973_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_148_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17527_ _21802_/Q _17417_/C _17417_/D _17526_/B vssd1 vssd1 vccd1 vccd1 _17528_/B
+ sky130_fd_sc_hd__a22o_1
X_14739_ _14739_/A _14739_/B vssd1 vssd1 vccd1 vccd1 _14742_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15698__B _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17458_ _17458_/A _17458_/B _17458_/C vssd1 vssd1 vccd1 vccd1 _17461_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_7_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16409_ _16409_/A _16409_/B vssd1 vssd1 vccd1 vccd1 _16410_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17389_ _17488_/A _17488_/B vssd1 vssd1 vccd1 vccd1 _17489_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19128_ _19291_/A _19129_/C _19129_/A vssd1 vssd1 vccd1 vccd1 _19130_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19693__A1 _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14506__A1 _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19059_ _19373_/B _19060_/B _19060_/C _19060_/D vssd1 vssd1 vccd1 vccd1 _19059_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_125_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22070_ _22080_/CLK _22070_/D fanout639/X vssd1 vssd1 vccd1 vccd1 mstream_o[6] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_125_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_516 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21021_ _20851_/Y _20856_/A _21135_/A _21020_/X vssd1 vssd1 vccd1 vccd1 _21135_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout383_A _16173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17434__A _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17759__A1 _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17759__B2 _18008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21923_ _21923_/CLK _21923_/D vssd1 vssd1 vccd1 vccd1 hold163/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout550_A _21733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21854_ _22106_/CLK _21854_/D vssd1 vssd1 vccd1 vccd1 hold212/A sky130_fd_sc_hd__dfxtp_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11256__A0 _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20805_ _20806_/A _20806_/B vssd1 vssd1 vccd1 vccd1 _20999_/B sky130_fd_sc_hd__or2_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20515__B1 _15626_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21785_ _21788_/CLK _21785_/D vssd1 vssd1 vccd1 vccd1 _21785_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_38_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20736_ _20736_/A _20857_/B vssd1 vssd1 vccd1 vccd1 _20738_/B sky130_fd_sc_hd__or2_1
XFILLER_0_37_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16195__B1 _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17931__A1 _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20667_ _20667_/A _20667_/B vssd1 vssd1 vccd1 vccd1 _20708_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12220__A2 _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20598_ _20598_/A vssd1 vssd1 vccd1 vccd1 _20600_/B sky130_fd_sc_hd__inv_2
XANTENNA__13559__D _14663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16498__B2 _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13070_ _13067_/X _13068_/Y _12929_/B _12928_/Y vssd1 vssd1 vccd1 vccd1 _13072_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_130_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12021_ _12070_/A _12118_/A vssd1 vssd1 vccd1 vccd1 _12071_/A sky130_fd_sc_hd__and2_1
X_21219_ _21220_/B _21220_/A vssd1 vssd1 vccd1 vccd1 _21275_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__19987__A2 fanout96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17998__A1 _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17998__B2 _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14968__A _14968_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13294__D _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout560 _21731_/Q vssd1 vssd1 vccd1 vccd1 _14621_/D sky130_fd_sc_hd__buf_4
XANTENNA__20689__B _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout571 _12268_/B vssd1 vssd1 vccd1 vccd1 _12246_/D sky130_fd_sc_hd__buf_4
X_16760_ _17206_/B _17277_/A vssd1 vssd1 vccd1 vccd1 _16828_/A sky130_fd_sc_hd__nand2_1
Xfanout582 _13985_/A vssd1 vssd1 vccd1 vccd1 _12269_/D sky130_fd_sc_hd__clkbuf_8
X_13972_ _13972_/A _13972_/B vssd1 vssd1 vccd1 vccd1 _14117_/A sky130_fd_sc_hd__nor2_1
Xfanout593 _11122_/A vssd1 vssd1 vccd1 vccd1 _11325_/A1 sky130_fd_sc_hd__buf_4
X_15711_ _15712_/A _15711_/B vssd1 vssd1 vccd1 vccd1 _15711_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13591__B _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ _12924_/A _12924_/B _12924_/C vssd1 vssd1 vccd1 vccd1 _12923_/X sky130_fd_sc_hd__and3_1
XANTENNA__17063__B _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16691_ _16691_/A _16691_/B _16691_/C vssd1 vssd1 vccd1 vccd1 _16730_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_115_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18430_ _18430_/A _18430_/B vssd1 vssd1 vccd1 vccd1 _18440_/A sky130_fd_sc_hd__nand2_1
X_15642_ _16031_/A _15643_/B vssd1 vssd1 vccd1 vccd1 _15642_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_154_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ _12855_/A _12855_/B vssd1 vssd1 vccd1 vccd1 _12966_/B sky130_fd_sc_hd__or2_1
XANTENNA__12039__A2 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20909__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11247__B1 _11246_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18361_ _18360_/A _18360_/B _18360_/C vssd1 vssd1 vccd1 vccd1 _18363_/C sky130_fd_sc_hd__a21o_1
X_11805_ _11805_/A _11805_/B _11805_/C vssd1 vssd1 vccd1 vccd1 _11805_/X sky130_fd_sc_hd__and3_2
XFILLER_0_150_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15573_ _15700_/A vssd1 vssd1 vccd1 vccd1 _15575_/D sky130_fd_sc_hd__inv_2
XFILLER_0_96_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ _14248_/A _12785_/B _14384_/D _14391_/B vssd1 vssd1 vccd1 vccd1 _12787_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19372__B1 _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17312_ _17313_/A _17313_/B vssd1 vssd1 vccd1 vccd1 _17312_/X sky130_fd_sc_hd__and2_2
XFILLER_0_28_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14524_ _14524_/A _14524_/B _14524_/C vssd1 vssd1 vccd1 vccd1 _14526_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_12_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18292_ _18292_/A _18292_/B vssd1 vssd1 vccd1 vccd1 _18292_/Y sky130_fd_sc_hd__xnor2_2
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11736_ _11736_/A _11736_/B _11736_/C vssd1 vssd1 vccd1 vccd1 _11750_/A sky130_fd_sc_hd__nand3_2
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17243_ _17243_/A _17243_/B _17243_/C vssd1 vssd1 vccd1 vccd1 _17245_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_154_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14455_ _14379_/A _14379_/C _14379_/B vssd1 vssd1 vccd1 vccd1 _14494_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ _11667_/A _11667_/B vssd1 vssd1 vccd1 vccd1 _11668_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20809__A1 _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13406_ _13860_/A _14018_/C vssd1 vssd1 vccd1 vccd1 _13410_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17174_ hold156/X fanout7/X _11553_/Y vssd1 vssd1 vccd1 vccd1 _17174_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_141_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14386_ _14537_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _14387_/B sky130_fd_sc_hd__and2_1
XFILLER_0_107_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11598_ _12020_/A _12403_/A _12511_/A _12326_/D vssd1 vssd1 vccd1 vccd1 _11599_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18622__B _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16125_ _15991_/B _15992_/Y _16123_/Y _16124_/X vssd1 vssd1 vccd1 vccd1 _16127_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13337_ _13338_/A _13338_/B _13338_/C vssd1 vssd1 vccd1 vccd1 _13337_/X sky130_fd_sc_hd__and3_1
XFILLER_0_106_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20590__D _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16056_ _16056_/A _16056_/B vssd1 vssd1 vccd1 vccd1 _16067_/A sky130_fd_sc_hd__or2_1
XFILLER_0_122_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13766__B _14218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15161__B2 _21733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13268_ _13154_/A _13153_/A _13153_/B vssd1 vssd1 vccd1 vccd1 _13273_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__17238__B _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15007_ _15006_/B _15006_/C _15006_/A vssd1 vssd1 vccd1 vccd1 _15007_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_20_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12219_ _12219_/A _12219_/B _12219_/C vssd1 vssd1 vccd1 vccd1 _12226_/A sky130_fd_sc_hd__nand3_1
XANTENNA__19734__A _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13199_ _13199_/A _13199_/B _13199_/C vssd1 vssd1 vccd1 vccd1 _13199_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__20319__A2_N _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19815_ _19654_/A _19653_/A _19653_/B _19649_/B _19649_/A vssd1 vssd1 vccd1 vccd1
+ _19816_/B sky130_fd_sc_hd__o32ai_4
XANTENNA__14878__A _21769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16958_ _16958_/A _16958_/B vssd1 vssd1 vccd1 vccd1 _16958_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_1070 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19746_ _20101_/A _20101_/B _19868_/B vssd1 vssd1 vccd1 vccd1 _19746_/X sky130_fd_sc_hd__and3_1
XFILLER_0_56_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15909_ _15909_/A _15909_/B vssd1 vssd1 vccd1 vccd1 _15948_/A sky130_fd_sc_hd__or2_1
XFILLER_0_79_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19677_ _19678_/A _19678_/B vssd1 vssd1 vccd1 vccd1 _19677_/Y sky130_fd_sc_hd__nor2_1
X_16889_ _16876_/A _16876_/C _16876_/B vssd1 vssd1 vccd1 vccd1 _16890_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11506__S _11545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17610__B1 _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18628_ _18628_/A _18628_/B vssd1 vssd1 vccd1 vccd1 _18630_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18559_ _18559_/A _18559_/B vssd1 vssd1 vccd1 vccd1 _18561_/B sky130_fd_sc_hd__and2_1
XFILLER_0_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21570_ mstream_o[33] _11045_/X _21579_/S vssd1 vssd1 vccd1 vccd1 _22097_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_90_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_12 _11331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_23 _11339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20521_ _20686_/A vssd1 vssd1 vccd1 vccd1 _20523_/D sky130_fd_sc_hd__inv_2
XFILLER_0_144_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_34 _11412_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout131_A _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_45 hold247/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_56 hold270/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_67 hold274/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_78 hold277/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20452_ _20302_/B _20302_/Y _20450_/X _20451_/Y vssd1 vssd1 vccd1 vccd1 _20499_/A
+ sky130_fd_sc_hd__o211a_2
XANTENNA_89 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11410__A0 _11409_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20383_ _20788_/A _21146_/B vssd1 vssd1 vccd1 vccd1 _20918_/A sky130_fd_sc_hd__or2_2
XFILLER_0_28_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15152__B2 _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22053_ _22063_/CLK _22053_/D vssd1 vssd1 vccd1 vccd1 hold309/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__19644__A _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21004_ _21000_/Y _21001_/X _20871_/X _20873_/X vssd1 vssd1 vccd1 vccd1 _21005_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16987__B _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14788__A _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11627__D _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11416__S _11446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21906_ _21906_/CLK _21906_/D vssd1 vssd1 vccd1 vccd1 hold89/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13823__A1_N _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19810__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_672 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12458__D _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17611__B _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21837_ _21837_/CLK _21837_/D vssd1 vssd1 vccd1 vccd1 _21837_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_65_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12570_ _12570_/A _12570_/B _12570_/C vssd1 vssd1 vccd1 vccd1 _12572_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21768_ _21789_/CLK _21768_/D vssd1 vssd1 vccd1 vccd1 _21768_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__12441__A2 _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12755__B _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20719_ _20719_/A _20719_/B vssd1 vssd1 vccd1 vccd1 _20720_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_81_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11521_ _11520_/X _19223_/B _11521_/S vssd1 vssd1 vccd1 vccd1 _21845_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_25_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15915__B1 _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21699_ _22096_/CLK _21699_/D vssd1 vssd1 vccd1 vccd1 hold106/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14240_ _14240_/A _14240_/B vssd1 vssd1 vccd1 vccd1 _14260_/A sky130_fd_sc_hd__xor2_2
X_11452_ _11451_/X _17557_/A _11470_/S vssd1 vssd1 vccd1 vccd1 _21822_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14194__A2 _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19538__B _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13289__D _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20691__C _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13867__A _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14171_ _14171_/A _14171_/B vssd1 vssd1 vccd1 vccd1 _14173_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_104_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11383_ _11382_/X _16860_/C _11401_/S vssd1 vssd1 vccd1 vccd1 _21799_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12771__A _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19257__C _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13122_ _13121_/B _13121_/C _13121_/A vssd1 vssd1 vccd1 vccd1 _13124_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_104_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15694__A2 _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13053_ _12913_/A _12913_/C _12913_/B vssd1 vssd1 vccd1 vccd1 _13054_/C sky130_fd_sc_hd__a21bo_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17930_ _19123_/A _19123_/B _19262_/C _19414_/C vssd1 vssd1 vccd1 vccd1 _17932_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_30_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12004_ _12897_/C _12155_/B _12214_/C _12403_/B vssd1 vssd1 vccd1 vccd1 _12004_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_79_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17861_ _18873_/A _18849_/A _19227_/C _19227_/D vssd1 vssd1 vccd1 vccd1 _17861_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_139_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14698__A _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16812_ _17029_/A _17029_/B _17063_/C _17086_/C vssd1 vssd1 vccd1 vccd1 _16816_/A
+ sky130_fd_sc_hd__and4_1
X_19600_ _19732_/B _19972_/C _20249_/B _19732_/A vssd1 vssd1 vccd1 vccd1 _19603_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13457__A1 _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17792_ _19123_/A _19123_/B _18789_/B _21040_/A vssd1 vssd1 vccd1 vccd1 _17794_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13457__B2 _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout390 _21771_/Q vssd1 vssd1 vccd1 vccd1 _12420_/D sky130_fd_sc_hd__buf_4
X_19531_ _19531_/A _20671_/B vssd1 vssd1 vccd1 vccd1 _19532_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16743_ _16813_/A _16743_/B _16743_/C _17013_/D vssd1 vssd1 vccd1 vccd1 _16743_/X
+ sky130_fd_sc_hd__and4_1
X_13955_ _13952_/Y _13953_/X _13802_/Y _13804_/X vssd1 vssd1 vccd1 vccd1 _13956_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_17_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17224__D _17324_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12906_ _14712_/B _14386_/B _14384_/C _14712_/A vssd1 vssd1 vccd1 vccd1 _12906_/X
+ sky130_fd_sc_hd__a22o_1
X_19462_ _19308_/A _19308_/B _19306_/X vssd1 vssd1 vccd1 vccd1 _19464_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16674_ _16674_/A _16674_/B vssd1 vssd1 vccd1 vccd1 _16676_/C sky130_fd_sc_hd__xnor2_1
X_13886_ _13757_/X _13795_/A _13884_/Y _13885_/X vssd1 vssd1 vccd1 vccd1 _13886_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_124_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18413_ _18413_/A vssd1 vssd1 vccd1 vccd1 _18413_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_154_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15625_ _15625_/A _15625_/B vssd1 vssd1 vccd1 vccd1 _15626_/B sky130_fd_sc_hd__or2_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19393_ _19393_/A _19393_/B _19543_/B vssd1 vssd1 vccd1 vccd1 _19395_/B sky130_fd_sc_hd__nand3_1
X_12837_ _12837_/A _12837_/B _12837_/C vssd1 vssd1 vccd1 vccd1 _12838_/B sky130_fd_sc_hd__or3_1
XFILLER_0_124_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16418__A _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11850__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18344_ _19723_/A _19092_/C vssd1 vssd1 vccd1 vccd1 _18348_/A sky130_fd_sc_hd__nand2_1
X_15556_ _15556_/A _15556_/B vssd1 vssd1 vccd1 vccd1 _15558_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__16159__B1 _21754_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21043__B _21841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11235__A3 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ _12648_/X _12650_/X _12765_/X _12766_/Y vssd1 vssd1 vccd1 vccd1 _12768_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_83_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_675 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14507_ _14508_/A _15022_/B _14508_/C _14508_/D vssd1 vssd1 vccd1 vccd1 _14507_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18275_ _18275_/A _18275_/B vssd1 vssd1 vccd1 vccd1 _18277_/B sky130_fd_sc_hd__xnor2_1
X_11719_ _12781_/D _12444_/B vssd1 vssd1 vccd1 vccd1 _11723_/A sky130_fd_sc_hd__nand2_1
X_15487_ _15487_/A _15487_/B vssd1 vssd1 vccd1 vccd1 _15490_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_154_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12699_ _12585_/Y _12587_/X _12696_/X _12698_/Y vssd1 vssd1 vccd1 vccd1 _12701_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17226_ _17224_/X _17226_/B vssd1 vssd1 vccd1 vccd1 _17227_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_114_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14438_ _14438_/A _14438_/B vssd1 vssd1 vccd1 vccd1 _14439_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12196__A1 _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12196__B2 _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17157_ _17156_/A _17156_/B _17156_/C vssd1 vssd1 vccd1 vccd1 _17158_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_4_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14369_ _14368_/B _14513_/B _14368_/A vssd1 vssd1 vccd1 vccd1 _14370_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_80_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15695__C _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16108_ _16108_/A _16212_/B vssd1 vssd1 vccd1 vccd1 _16110_/B sky130_fd_sc_hd__or2_1
X_17088_ _17146_/A _17086_/C _17123_/C _17146_/B vssd1 vssd1 vccd1 vccd1 _17089_/C
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_40_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20106__C _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16039_ _16414_/A _16040_/C _16268_/B _16391_/A vssd1 vssd1 vccd1 vccd1 _16042_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18623__A2 _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16600__B _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19729_ _19729_/A _19729_/B vssd1 vssd1 vccd1 vccd1 _19737_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11236__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout179_A _17443_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13017__A _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21391__A0 _15070_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14948__B2 _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16328__A _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout346_A _16396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_379 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21622_ _21939_/CLK _21622_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[85] sky130_fd_sc_hd__dfrtp_4
XANTENNA__14774__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21553_ mstream_o[16] hold73/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22080_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_63_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout513_A _21741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20792__B _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20504_ _20501_/Y _20502_/X _20351_/Y _20353_/X vssd1 vssd1 vccd1 vccd1 _20504_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21484_ hold180/X sstream_i[61] _21507_/S vssd1 vssd1 vccd1 vccd1 _22011_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_7_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16570__B1 _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14790__B _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12187__A1 _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12187__B2 _12242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20435_ _20436_/B _20436_/A vssd1 vssd1 vccd1 vccd1 _20571_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_16_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11934__A1 _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11919__B _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20366_ _20366_/A _20366_/B vssd1 vssd1 vccd1 vccd1 _20367_/B sky130_fd_sc_hd__or2_1
XFILLER_0_3_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22105_ _22105_/CLK _22105_/D _11089_/A vssd1 vssd1 vccd1 vccd1 mstream_o[41] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20297_ _20115_/X _20118_/Y _20449_/B _20296_/X vssd1 vssd1 vccd1 vccd1 _20299_/A
+ sky130_fd_sc_hd__o211a_1
X_22036_ _22038_/CLK _22036_/D vssd1 vssd1 vccd1 vccd1 hold305/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__21409__A _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19093__B _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17606__B _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20032__B _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13740_ _13736_/Y _13737_/X _13581_/A _13581_/Y vssd1 vssd1 vccd1 vccd1 _13800_/B
+ sky130_fd_sc_hd__a211oi_2
X_10952_ hold78/A hold276/A hold263/A hold273/A vssd1 vssd1 vccd1 vccd1 _10952_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__21382__A0 _14605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13671_ _14133_/D _13983_/B _16409_/B vssd1 vssd1 vccd1 vccd1 _13671_/X sky130_fd_sc_hd__and3_1
X_10883_ hold243/A hold252/A vssd1 vssd1 vccd1 vccd1 _10885_/C sky130_fd_sc_hd__xnor2_1
X_15410_ _15931_/A _15931_/B _16396_/A _16266_/C vssd1 vssd1 vccd1 vccd1 _15547_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_38_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12622_ _12621_/C _13573_/D _12732_/A _12620_/Y vssd1 vssd1 vccd1 vccd1 _12622_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_16390_ _16390_/A _16390_/B vssd1 vssd1 vccd1 vccd1 _16392_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15341_ _15342_/A _15342_/B vssd1 vssd1 vccd1 vccd1 _15341_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_93_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12553_ _12551_/X _12553_/B vssd1 vssd1 vccd1 vccd1 _12554_/B sky130_fd_sc_hd__and2b_1
XANTENNA__14981__A _21766_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1192 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11504_ _11507_/A1 t1y[18] t0x[18] _11507_/B2 vssd1 vssd1 vccd1 vccd1 _11504_/X sky130_fd_sc_hd__a22o_1
X_18060_ _19438_/B _18640_/B _19092_/C _19438_/A vssd1 vssd1 vccd1 vccd1 _18061_/B
+ sky130_fd_sc_hd__a22oi_2
X_15272_ _15001_/B _15091_/X _15094_/A _15094_/B vssd1 vssd1 vccd1 vccd1 _15279_/A
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_136_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12484_ _12484_/A _12484_/B _12484_/C vssd1 vssd1 vccd1 vccd1 _12484_/X sky130_fd_sc_hd__and3_1
XFILLER_0_81_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17011_ _16980_/A _16980_/C _16980_/B vssd1 vssd1 vccd1 vccd1 _17028_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14223_ _14222_/A _14222_/B _14222_/C vssd1 vssd1 vccd1 vccd1 _14224_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_124_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13914__A2 _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11435_ _11447_/A1 hold220/A fanout48/X hold161/A vssd1 vssd1 vccd1 vccd1 _11435_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16313__B1 _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14154_ _15159_/D _14155_/C _14155_/D _14936_/D vssd1 vssd1 vccd1 vccd1 _14157_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11366_ _11124_/A hold249/A fanout45/X hold177/X vssd1 vssd1 vccd1 vccd1 _11366_/X
+ sky130_fd_sc_hd__a22o_1
X_13105_ _13250_/C vssd1 vssd1 vccd1 vccd1 _13107_/A sky130_fd_sc_hd__inv_2
XFILLER_0_46_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14085_ _14557_/D _14084_/X _14083_/X vssd1 vssd1 vccd1 vccd1 _14086_/B sky130_fd_sc_hd__a21bo_1
X_11297_ _11325_/A1 t2y[18] t0y[18] _11507_/A1 vssd1 vssd1 vccd1 vccd1 _11297_/X sky130_fd_sc_hd__a22o_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18962_ _19123_/A _20247_/D _20721_/C vssd1 vssd1 vccd1 vccd1 _18964_/B sky130_fd_sc_hd__a21oi_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14875__B1 _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ _14367_/A _15217_/A _13169_/A _13036_/D vssd1 vssd1 vccd1 vccd1 _13169_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17913_ _17913_/A _17913_/B vssd1 vssd1 vccd1 vccd1 _17921_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11689__B1 _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18893_ _20178_/D _18894_/B _18894_/C _18894_/D vssd1 vssd1 vccd1 vccd1 _18895_/A
+ sky130_fd_sc_hd__a22o_1
X_17844_ _18703_/A _19030_/C _17720_/X _17725_/A vssd1 vssd1 vccd1 vccd1 _17845_/B
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__20412__A2 _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11564__B _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17775_ _17772_/Y _17773_/X _17647_/X _17649_/X vssd1 vssd1 vccd1 vccd1 _17776_/B
+ sky130_fd_sc_hd__a211o_1
X_14987_ _15085_/A _15502_/A _14984_/Y _14985_/X vssd1 vssd1 vccd1 vccd1 _14990_/B
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_135_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11056__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16726_ _17146_/A _17526_/B _17223_/A _17146_/B vssd1 vssd1 vccd1 vccd1 _16727_/C
+ sky130_fd_sc_hd__a22o_1
X_19514_ _19503_/Y _19514_/B _19514_/C vssd1 vssd1 vccd1 vccd1 _19676_/A sky130_fd_sc_hd__and3b_1
XFILLER_0_152_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13938_ _13939_/A _13939_/B _13939_/C vssd1 vssd1 vccd1 vccd1 _13938_/X sky130_fd_sc_hd__and3_1
XANTENNA__16919__A2 _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19445_ _19445_/A _19445_/B vssd1 vssd1 vccd1 vccd1 _19847_/A sky130_fd_sc_hd__and2_2
X_16657_ _17178_/B _16657_/B _16657_/C _16657_/D vssd1 vssd1 vccd1 vccd1 _16657_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__11861__B1 _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13869_ _13865_/X _13867_/Y _13710_/X _13713_/B vssd1 vssd1 vccd1 vccd1 _13870_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_1081 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11580__A _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15608_ _15422_/X _15426_/C _15693_/B _15606_/Y vssd1 vssd1 vccd1 vccd1 _15608_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19376_ _19376_/A _19376_/B vssd1 vssd1 vccd1 vccd1 _19386_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_29_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16588_ _21825_/Q _17434_/B _17433_/A _16734_/B vssd1 vssd1 vccd1 vccd1 _16588_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_146_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18327_ _18328_/A _18328_/B _18328_/C vssd1 vssd1 vccd1 vccd1 _18327_/X sky130_fd_sc_hd__a21o_2
X_15539_ _16369_/A _16399_/A _15539_/C _15539_/D vssd1 vssd1 vccd1 vccd1 _15663_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_60_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18258_ _18255_/Y _18402_/A _18857_/B _19201_/B vssd1 vssd1 vccd1 vccd1 _18402_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_127_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17209_ _17207_/X _17209_/B vssd1 vssd1 vccd1 vccd1 _17210_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18189_ _18187_/Y _18332_/A _18789_/A _19089_/B vssd1 vssd1 vccd1 vccd1 _18332_/B
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__16314__C _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12842__C _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20220_ _20220_/A _20220_/B vssd1 vssd1 vccd1 vccd1 _20220_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16304__B1 _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11739__B _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20100__A1 _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19906__B _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20100__B2 _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_11_clk_i _21806_/CLK vssd1 vssd1 vccd1 vccd1 _22038_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_12_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17129__D _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20151_ _20151_/A _20151_/B vssd1 vssd1 vccd1 vccd1 _20153_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_100_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16611__A _21824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16968__D _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20082_ _19792_/B _20081_/Y _20080_/X vssd1 vssd1 vccd1 vccd1 _20083_/B sky130_fd_sc_hd__o21a_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20133__A _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16607__A1 _17557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout296_A _21796_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16607__B2 _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21888_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16083__A2 _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17280__A1 _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout463_A _21753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18538__A _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17442__A _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20984_ _20984_/A _20984_/B vssd1 vssd1 vccd1 vccd1 _21005_/A sky130_fd_sc_hd__or2_1
XFILLER_0_79_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12644__A2 _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11921__C _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_984 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21605_ _21934_/CLK _21605_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[68] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15112__D _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21536_ hold283/X sstream_i[113] _21536_/S vssd1 vssd1 vccd1 vccd1 _22063_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_91_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_hold306_A hold306/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21467_ hold123/X sstream_i[44] _21494_/S vssd1 vssd1 vccd1 vccd1 _21994_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14306__A _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ hold148/X fanout51/X fanout48/X hold251/A vssd1 vssd1 vccd1 vccd1 _11220_/X
+ sky130_fd_sc_hd__a22o_1
X_20418_ _21842_/Q _20270_/C _20419_/C _20419_/D vssd1 vssd1 vccd1 vccd1 _20420_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_102_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21398_ hold167/X _21397_/X _21403_/S vssd1 vssd1 vccd1 vccd1 _21940_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_120_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11151_ hold248/X _11126_/A fanout45/X hold298/A vssd1 vssd1 vccd1 vccd1 _11151_/X
+ sky130_fd_sc_hd__a22o_1
X_20349_ _20498_/A _20348_/C _20348_/A vssd1 vssd1 vccd1 vccd1 _20350_/B sky130_fd_sc_hd__o21a_1
XANTENNA__16521__A _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19535__C _19692_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13864__B _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11082_ _10950_/Y hold62/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21677_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_41_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14910_ _14910_/A _14910_/B vssd1 vssd1 vccd1 vccd1 _15206_/A sky130_fd_sc_hd__nor2_2
X_22019_ _22020_/CLK _22019_/D vssd1 vssd1 vccd1 vccd1 hold186/A sky130_fd_sc_hd__dfxtp_1
X_15890_ _12291_/B _15888_/Y _15889_/X vssd1 vssd1 vccd1 vccd1 _15890_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12883__A2 _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14841_ _14840_/B _14840_/C _14840_/A vssd1 vssd1 vccd1 vccd1 _14841_/X sky130_fd_sc_hd__a21o_1
XANTENNA__14085__A1 _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17560_ _17559_/B _17559_/C _17559_/A vssd1 vssd1 vccd1 vccd1 _17562_/B sky130_fd_sc_hd__a21o_1
X_14772_ _15829_/C _14615_/X _14618_/A _14618_/B vssd1 vssd1 vccd1 vccd1 _14773_/B
+ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__19012__A2 _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11984_ _12268_/A _12639_/A vssd1 vssd1 vccd1 vccd1 _11986_/B sky130_fd_sc_hd__and2_1
XFILLER_0_59_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14695__B _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18167__B _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16511_ _17029_/A _17029_/B _16860_/C _16917_/C vssd1 vssd1 vccd1 vccd1 _16564_/A
+ sky130_fd_sc_hd__nand4_2
X_13723_ _14027_/A _16286_/A _13724_/C _13724_/D vssd1 vssd1 vccd1 vccd1 _13723_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_105_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17491_ _17614_/A vssd1 vssd1 vccd1 vccd1 _17493_/C sky130_fd_sc_hd__inv_2
X_10935_ mstream_o[54] _10934_/Y _10992_/S vssd1 vssd1 vccd1 vccd1 _21591_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17502__D _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18771__A1 _19092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19230_ _19230_/A _19382_/B _19230_/C _19230_/D vssd1 vssd1 vccd1 vccd1 _19230_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_129_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16442_ _16868_/A _17223_/A _16860_/C _16734_/B vssd1 vssd1 vccd1 vccd1 _16442_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__18771__B2 _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14388__A2 _14217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13654_ _13500_/C _13501_/X _13652_/Y _13653_/X vssd1 vssd1 vccd1 vccd1 _13656_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_155_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10866_ _10866_/A _10866_/B _10864_/Y vssd1 vssd1 vccd1 vccd1 _10867_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_14_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19161_ _19162_/A _19162_/B vssd1 vssd1 vccd1 vccd1 _19161_/Y sky130_fd_sc_hd__nor2_1
X_12605_ _12605_/A _12605_/B _12606_/B vssd1 vssd1 vccd1 vccd1 _12818_/A sky130_fd_sc_hd__or3_2
X_16373_ _16373_/A _16373_/B vssd1 vssd1 vccd1 vccd1 _16379_/A sky130_fd_sc_hd__xnor2_2
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19279__A _19430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13585_ _13428_/A _13428_/Y _13583_/X _13584_/Y vssd1 vssd1 vccd1 vccd1 _13648_/A
+ sky130_fd_sc_hd__o211a_1
X_10797_ _16314_/D vssd1 vssd1 vccd1 vccd1 _10797_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18112_ _18253_/A _18111_/Y _18703_/A _19201_/B vssd1 vssd1 vccd1 vccd1 _18253_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_53_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15324_ _15324_/A _15324_/B vssd1 vssd1 vccd1 vccd1 _15326_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_147_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19092_ _19092_/A _19092_/B _19092_/C _19262_/C vssd1 vssd1 vccd1 vccd1 _19095_/B
+ sky130_fd_sc_hd__nand4_1
X_12536_ _12534_/X _12536_/B vssd1 vssd1 vccd1 vccd1 _12537_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_81_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18043_ _18164_/B _18042_/C _18042_/A vssd1 vssd1 vccd1 vccd1 _18044_/C sky130_fd_sc_hd__a21o_1
X_15255_ _16196_/A _15653_/C _15911_/C _16374_/A vssd1 vssd1 vccd1 vccd1 _15258_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12467_ _12364_/A _12364_/C _12364_/B vssd1 vssd1 vccd1 vccd1 _12468_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_22_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18911__A _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14206_ _14203_/X _14204_/Y _14070_/B _14072_/A vssd1 vssd1 vccd1 vccd1 _14207_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_111_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11418_ hold280/A fanout28/X _11417_/X vssd1 vssd1 vccd1 vccd1 _11418_/X sky130_fd_sc_hd__a21o_1
X_15186_ _15296_/A _15185_/C _15185_/A vssd1 vssd1 vccd1 vccd1 _15186_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_1_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12398_ _12398_/A vssd1 vssd1 vccd1 vccd1 _12605_/A sky130_fd_sc_hd__inv_2
X_14137_ _14138_/A _16084_/C _16084_/D _14463_/D vssd1 vssd1 vccd1 vccd1 _14137_/X
+ sky130_fd_sc_hd__a22o_1
X_11349_ _11349_/A1 t2y[31] t0y[31] _11089_/B vssd1 vssd1 vccd1 vccd1 _11349_/X sky130_fd_sc_hd__a22o_1
X_19994_ _20863_/C _20419_/A _19995_/C _20138_/A vssd1 vssd1 vccd1 vccd1 _19997_/A
+ sky130_fd_sc_hd__a22o_1
X_14068_ _14068_/A _14209_/B _14068_/C vssd1 vssd1 vccd1 vccd1 _14070_/B sky130_fd_sc_hd__nand3_2
X_18945_ _18944_/B _18944_/C _18944_/A vssd1 vssd1 vccd1 vccd1 _18946_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_20_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12323__A1 _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__A _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13019_ _13155_/B _13155_/C _21768_/Q _13018_/B vssd1 vssd1 vccd1 vccd1 _13020_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18876_ _18876_/A _18876_/B _18876_/C vssd1 vssd1 vccd1 vccd1 _18878_/B sky130_fd_sc_hd__nand3_2
X_17827_ _17828_/A _17828_/B vssd1 vssd1 vccd1 vccd1 _17967_/A sky130_fd_sc_hd__nor2_2
XANTENNA__14076__A1 _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11725__D _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19003__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17758_ _19664_/B _18008_/A _18616_/D vssd1 vssd1 vccd1 vccd1 _17758_/X sky130_fd_sc_hd__and3_1
XFILLER_0_7_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16709_ _16675_/X _16706_/Y _16705_/Y _16705_/A vssd1 vssd1 vccd1 vccd1 _16712_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_49_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17689_ _17689_/A _17689_/B _17689_/C _17689_/D vssd1 vssd1 vccd1 vccd1 _17689_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_76_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout18 fanout19/X vssd1 vssd1 vccd1 vccd1 fanout18/X sky130_fd_sc_hd__clkbuf_4
X_19428_ _19439_/A _20242_/D _19286_/X _19117_/X _20247_/C vssd1 vssd1 vccd1 vccd1
+ _19433_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_18_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout29 _11124_/Y vssd1 vssd1 vccd1 vccd1 fanout29/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_58_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19359_ _19358_/B _19358_/C _19347_/Y vssd1 vssd1 vccd1 vccd1 _19359_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_73_932 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16606__A _17557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15510__A _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20128__A _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21321_ _21321_/A _21321_/B vssd1 vssd1 vccd1 vccd1 _21322_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout211_A _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout309_A _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21252_ hold171/X _11553_/Y _21250_/X _21251_/X vssd1 vssd1 vccd1 vccd1 hold172/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18278__B1 _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19636__B _19636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20203_ _20053_/X _20203_/B vssd1 vssd1 vccd1 vccd1 _20205_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_25_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21183_ _21183_/A _21183_/B vssd1 vssd1 vccd1 vccd1 _21185_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20134_ _20275_/A vssd1 vssd1 vccd1 vccd1 _20136_/D sky130_fd_sc_hd__inv_2
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout580_A _21727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14499__C _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20065_ _20216_/B _20065_/B vssd1 vssd1 vccd1 vccd1 _20066_/B sky130_fd_sc_hd__or2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19802__D _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17172__A _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_305 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold256_A hold256/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_316 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_327 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_338 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20967_ _21085_/A vssd1 vssd1 vccd1 vccd1 _20969_/D sky130_fd_sc_hd__inv_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20560__A1 _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20898_ _20898_/A _20898_/B vssd1 vssd1 vccd1 vccd1 _20906_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__20560__B2 _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21422__A _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19702__B1 _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18434__C _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13370_ _16363_/A hold190/X _11063_/X fanout6/X _13369_/Y vssd1 vssd1 vccd1 vccd1
+ _13370_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_118_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12321_ _12530_/A _12319_/C _12420_/D _14621_/D vssd1 vssd1 vccd1 vccd1 _12322_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__10800__B2 _10792_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21519_ hold234/X sstream_i[96] _21528_/S vssd1 vssd1 vccd1 vccd1 _22046_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_106_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15040_ _15040_/A _15040_/B _15040_/C vssd1 vssd1 vccd1 vccd1 _15044_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_142_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14542__A2 _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12252_ _12258_/A _12252_/B vssd1 vssd1 vccd1 vccd1 _12259_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19546__B _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13875__A _21741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11203_ hold207/X fanout22/X _11202_/X vssd1 vssd1 vccd1 vccd1 _11203_/X sky130_fd_sc_hd__a21o_1
XANTENNA__20027__A2_N _20841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12183_ _12183_/A _12183_/B _12183_/C vssd1 vssd1 vccd1 vccd1 _12219_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_43_1135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17492__A1 _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13594__B _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ hold209/X fanout23/X _11133_/X vssd1 vssd1 vccd1 vccd1 _11134_/X sky130_fd_sc_hd__a21o_1
X_16991_ _16992_/B _16992_/A vssd1 vssd1 vccd1 vccd1 _16999_/B sky130_fd_sc_hd__and2b_1
XANTENNA__17492__B2 _21792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15942_ _15942_/A vssd1 vssd1 vccd1 vccd1 _16078_/B sky130_fd_sc_hd__inv_2
X_11065_ _11065_/A _11065_/B _11065_/C vssd1 vssd1 vccd1 vccd1 _11066_/B sky130_fd_sc_hd__and3_1
X_18730_ _18846_/A _18728_/X _18569_/Y _18572_/X vssd1 vssd1 vccd1 vccd1 _18826_/B
+ sky130_fd_sc_hd__o211a_1
X_18661_ _18661_/A _18661_/B _18661_/C vssd1 vssd1 vccd1 vccd1 _18664_/B sky130_fd_sc_hd__nand3_2
X_15873_ _15870_/A _15871_/X _15733_/B _15732_/Y vssd1 vssd1 vccd1 vccd1 _15874_/D
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__19281__B _19753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14824_ _14824_/A _14824_/B vssd1 vssd1 vccd1 vccd1 _14840_/A sky130_fd_sc_hd__xnor2_2
X_17612_ _17854_/B _21256_/A _17611_/C _17611_/D vssd1 vssd1 vccd1 vccd1 _17613_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_116_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18592_ _18592_/A _18592_/B vssd1 vssd1 vccd1 vccd1 _18593_/B sky130_fd_sc_hd__nand2_1
XTAP_3850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17543_ _20583_/A _19892_/A _19951_/B vssd1 vssd1 vccd1 vccd1 _17543_/X sky130_fd_sc_hd__and3_1
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14755_ _14755_/A _14755_/B vssd1 vssd1 vccd1 vccd1 _14758_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11967_ _11892_/X _11965_/Y _11964_/X _11944_/Y vssd1 vssd1 vccd1 vccd1 _11971_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_114_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13706_ _14306_/A _13997_/C _13707_/C _13707_/D vssd1 vssd1 vccd1 vccd1 _13708_/A
+ sky130_fd_sc_hd__a22o_1
X_10918_ _10917_/A _10917_/B _10919_/A vssd1 vssd1 vccd1 vccd1 _10924_/B sky130_fd_sc_hd__o21ba_1
X_17474_ _17474_/A _17474_/B vssd1 vssd1 vccd1 vccd1 _17475_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_128_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14686_ _14549_/Y _14553_/A _14809_/B _14685_/X vssd1 vssd1 vccd1 vccd1 _14688_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11898_ _11899_/A _11899_/B _11899_/C vssd1 vssd1 vccd1 vccd1 _11900_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16425_ _16344_/A _16344_/B _16342_/X vssd1 vssd1 vccd1 vccd1 _16431_/A sky130_fd_sc_hd__a21o_1
X_19213_ _19213_/A _19213_/B vssd1 vssd1 vccd1 vccd1 _19214_/B sky130_fd_sc_hd__xnor2_1
X_13637_ _13638_/A _13638_/B _13638_/C vssd1 vssd1 vccd1 vccd1 _13637_/X sky130_fd_sc_hd__and3_1
XFILLER_0_6_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13033__A2 _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10849_ _11065_/B _11065_/C _11065_/A vssd1 vssd1 vccd1 vccd1 _11066_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_26_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19144_ _19143_/B _19143_/C _19143_/A vssd1 vssd1 vccd1 vccd1 _19144_/Y sky130_fd_sc_hd__a21oi_2
X_16356_ _16356_/A _16356_/B vssd1 vssd1 vccd1 vccd1 _16359_/A sky130_fd_sc_hd__xnor2_2
X_13568_ _13690_/B _13568_/B vssd1 vssd1 vccd1 vccd1 _13568_/X sky130_fd_sc_hd__and2_1
XFILLER_0_41_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12673__B _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15307_ _15307_/A _15307_/B vssd1 vssd1 vccd1 vccd1 _15311_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_42_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19075_ _18914_/A _18914_/C _18914_/B vssd1 vssd1 vccd1 vccd1 _19076_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_42_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12519_ _12519_/A _12519_/B vssd1 vssd1 vccd1 vccd1 _12521_/C sky130_fd_sc_hd__xnor2_2
X_16287_ _16287_/A _16287_/B _16287_/C vssd1 vssd1 vccd1 vccd1 _16289_/A sky130_fd_sc_hd__and3_1
XFILLER_0_140_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13499_ _13496_/X _13497_/Y _13348_/B _13347_/Y vssd1 vssd1 vccd1 vccd1 _13500_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18026_ _18026_/A _18026_/B vssd1 vssd1 vccd1 vccd1 _18044_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15238_ _15238_/A _15238_/B vssd1 vssd1 vccd1 vccd1 _15240_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13741__B1 _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15169_ _15169_/A _15169_/B vssd1 vssd1 vccd1 vccd1 _15177_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout208 _19753_/B vssd1 vssd1 vccd1 vccd1 _19866_/D sky130_fd_sc_hd__clkbuf_8
Xfanout219 _18789_/B vssd1 vssd1 vccd1 vccd1 _19092_/C sky130_fd_sc_hd__buf_4
XANTENNA__14297__A1 _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19977_ _19977_/A _20098_/A _19977_/C vssd1 vssd1 vccd1 vccd1 _20098_/B sky130_fd_sc_hd__nand3_1
XANTENNA__14297__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11509__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18928_ _18767_/B _18773_/B _19546_/D _21833_/Q vssd1 vssd1 vccd1 vccd1 _18928_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18859_ _18859_/A _21261_/B _18859_/C _18859_/D vssd1 vssd1 vccd1 vccd1 _18860_/B
+ sky130_fd_sc_hd__nor4_1
XANTENNA__20411__A _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21870_ _21934_/CLK _21870_/D vssd1 vssd1 vccd1 vccd1 hold243/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__20130__B _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20821_ _20823_/A _20823_/B _20823_/C vssd1 vssd1 vccd1 vccd1 _20824_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout161_A _17324_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11244__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout259_A _19230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15549__A1 _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17720__A _17854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15549__B2 _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20752_ _20621_/B _20621_/Y _20750_/Y _20751_/X vssd1 vssd1 vccd1 vccd1 _20753_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_15_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20683_ _20683_/A _20683_/B vssd1 vssd1 vccd1 vccd1 _20684_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_135_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout426_A _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11035__A1 hold262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21098__A2 _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11586__A2 _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21304_ _21286_/A _21311_/B _21214_/A _21212_/B vssd1 vssd1 vccd1 vccd1 _21308_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21627__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21235_ _21236_/A _21236_/B _21236_/C vssd1 vssd1 vccd1 vccd1 _21255_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__12535__B2 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold240 hold240/A vssd1 vssd1 vccd1 vccd1 hold240/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 hold251/A vssd1 vssd1 vccd1 vccd1 hold251/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 hold262/A vssd1 vssd1 vccd1 vccd1 hold262/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold273 hold273/A vssd1 vssd1 vccd1 vccd1 hold273/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold284 hold284/A vssd1 vssd1 vccd1 vccd1 hold284/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21166_ _21059_/A _21061_/B _21059_/B vssd1 vssd1 vccd1 vccd1 _21270_/S sky130_fd_sc_hd__o21ba_1
Xhold295 hold295/A vssd1 vssd1 vccd1 vccd1 hold295/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20117_ _20119_/B _20119_/A vssd1 vssd1 vccd1 vccd1 _20118_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__11419__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21097_ _21097_/A _21097_/B vssd1 vssd1 vccd1 vccd1 _21105_/A sky130_fd_sc_hd__nand2_1
XANTENNA__15118__C _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout74_A _21849_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20048_ _20045_/Y _20188_/A _20590_/D _20193_/D vssd1 vssd1 vccd1 vccd1 _20188_/B
+ sky130_fd_sc_hd__and4bb_1
XTAP_3102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20230__B1 _15356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15415__A _15415_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12870_ _12869_/B _12869_/C _12869_/A vssd1 vssd1 vccd1 vccd1 _12870_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_38_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_102 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_113 sstream_i[66] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11821_ _11821_/A _11821_/B vssd1 vssd1 vccd1 vccd1 _11823_/C sky130_fd_sc_hd__xor2_2
XFILLER_0_96_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18148__D _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_124 v0z[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_135 v1z[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_146 v1z[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17052__D _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21999_ _22005_/CLK _21999_/D vssd1 vssd1 vccd1 vccd1 hold184/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_138_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20975__B _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_157 v2z[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14540_ _15373_/A _15373_/B _16268_/B _16266_/C vssd1 vssd1 vccd1 vccd1 _14543_/D
+ sky130_fd_sc_hd__nand4_2
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11274__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_168 v2z[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11752_ _11753_/A _11753_/B _11753_/C vssd1 vssd1 vccd1 vccd1 _11752_/X sky130_fd_sc_hd__and3_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_179 v2z[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14471_ _14471_/A _14471_/B vssd1 vssd1 vccd1 vccd1 _14472_/B sky130_fd_sc_hd__and2_1
XFILLER_0_95_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ _11683_/A _11683_/B vssd1 vssd1 vccd1 vccd1 _11685_/B sky130_fd_sc_hd__nand2_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16210_ _16211_/B vssd1 vssd1 vccd1 vccd1 _16210_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_3_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11026__A1 hold290/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13422_ _13419_/X _13569_/B _13290_/D _13292_/A vssd1 vssd1 vccd1 vccd1 _13423_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__13589__B _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17190_ _17191_/A _17191_/B vssd1 vssd1 vccd1 vccd1 _17190_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_52_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12493__B _12493_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12774__A1 _13018_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16141_ _16142_/B vssd1 vssd1 vccd1 vccd1 _16141_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_36_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13353_ _13353_/A _13353_/B _13353_/C vssd1 vssd1 vccd1 vccd1 _13353_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_3_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15300__D _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12304_ _12305_/B _12304_/B vssd1 vssd1 vccd1 vccd1 _12306_/B sky130_fd_sc_hd__and2b_1
X_16072_ _16070_/B _16070_/C _16070_/A vssd1 vssd1 vccd1 vccd1 _16072_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13284_ _13139_/X _13142_/X _13373_/A _13283_/Y vssd1 vssd1 vccd1 vccd1 _13373_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15023_ _15024_/A _15024_/B _15024_/C vssd1 vssd1 vccd1 vccd1 _15023_/X sky130_fd_sc_hd__a21o_1
X_19900_ _19897_/X _19898_/Y _19691_/X _19694_/X vssd1 vssd1 vccd1 vccd1 _19901_/B
+ sky130_fd_sc_hd__a211o_1
X_12235_ _12234_/A _12241_/A _12203_/X _12211_/Y vssd1 vssd1 vccd1 vccd1 _12235_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19831_ _19830_/B _19830_/C _19830_/A vssd1 vssd1 vccd1 vccd1 _19831_/Y sky130_fd_sc_hd__a21oi_2
X_12166_ _12115_/X _12133_/Y _12160_/A _12159_/Y vssd1 vssd1 vccd1 vccd1 _12168_/C
+ sky130_fd_sc_hd__a211oi_1
X_11117_ _10965_/Y hold45/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21711_/D sky130_fd_sc_hd__mux2_1
X_19762_ _19759_/A _19760_/Y _19578_/B _19581_/B vssd1 vssd1 vccd1 vccd1 _19763_/D
+ sky130_fd_sc_hd__o211ai_1
X_16974_ _17144_/A _17013_/D _17019_/C _17129_/B vssd1 vssd1 vccd1 vccd1 _16974_/Y
+ sky130_fd_sc_hd__a22oi_1
X_12097_ _12223_/A _12246_/C vssd1 vssd1 vccd1 vccd1 _12098_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11556__C _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18713_ _19337_/D _19201_/B _18713_/C _18713_/D vssd1 vssd1 vccd1 vccd1 _18713_/X
+ sky130_fd_sc_hd__and4_1
X_15925_ _15925_/A _15925_/B vssd1 vssd1 vccd1 vccd1 _15926_/B sky130_fd_sc_hd__nand2_1
X_11048_ _11048_/A _11048_/B vssd1 vssd1 vccd1 vccd1 _11048_/Y sky130_fd_sc_hd__xnor2_4
X_19693_ _19695_/A _20419_/A _19695_/C _19695_/D vssd1 vssd1 vccd1 vccd1 _19693_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15228__B1 _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15856_ _15857_/B _15857_/A vssd1 vssd1 vccd1 vccd1 _15856_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__21046__B _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18644_ _18644_/A _18644_/B vssd1 vssd1 vccd1 vccd1 _18664_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14807_ _14808_/A _14808_/B vssd1 vssd1 vccd1 vccd1 _14924_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_99_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15787_ _16409_/A _15788_/B _15788_/C _15973_/A vssd1 vssd1 vccd1 vccd1 _15789_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18575_ _18571_/Y _18573_/X _18456_/X _18459_/Y vssd1 vssd1 vccd1 vccd1 _18576_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_3680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12999_ _12865_/A _12864_/B _12862_/X vssd1 vssd1 vccd1 vccd1 _13000_/C sky130_fd_sc_hd__a21o_1
XTAP_3691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11064__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11265__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14738_ _14738_/A _14738_/B vssd1 vssd1 vccd1 vccd1 _14739_/B sky130_fd_sc_hd__xor2_4
X_17526_ _21802_/Q _17526_/B _18319_/B _18622_/B vssd1 vssd1 vccd1 vccd1 _17526_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_54_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17457_ _17345_/A _17345_/C _17345_/B vssd1 vssd1 vccd1 vccd1 _17458_/C sky130_fd_sc_hd__a21bo_1
X_14669_ _14667_/X _14669_/B vssd1 vssd1 vccd1 vccd1 _14670_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_28_943 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16408_ _16408_/A _16408_/B vssd1 vssd1 vccd1 vccd1 _16410_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17388_ _17388_/A _17388_/B vssd1 vssd1 vccd1 vccd1 _17488_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16339_ _16388_/B _16337_/Y _16225_/Y _16227_/Y vssd1 vssd1 vccd1 vccd1 _16340_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_6_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19127_ _19126_/A _19126_/B _19126_/C vssd1 vssd1 vccd1 vccd1 _19129_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19693__A2 _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19058_ _19373_/B _19060_/B _19060_/C _19060_/D vssd1 vssd1 vccd1 vccd1 _19058_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18009_ _18008_/A _19906_/A _20146_/B _18008_/B vssd1 vssd1 vccd1 vccd1 _18010_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21020_ _21129_/B _21018_/X _20886_/X _20888_/Y vssd1 vssd1 vccd1 vccd1 _21020_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21252__A2 _11553_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11740__A2 _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17208__A1 _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17208__B2 _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17434__B _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout376_A _14828_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17759__A2 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21922_ _21926_/CLK _21922_/D vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21853_ _21853_/CLK _21853_/D vssd1 vssd1 vccd1 vccd1 _21853_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_136_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout543_A _21735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20804_ _20999_/A _20804_/B vssd1 vssd1 vccd1 vccd1 _20806_/B sky130_fd_sc_hd__nand2_1
XANTENNA__12453__B1 _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20515__B2 _11550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21784_ _21821_/CLK _21784_/D vssd1 vssd1 vccd1 vccd1 _21784_/Q sky130_fd_sc_hd__dfxtp_2
X_20735_ _20857_/A _21311_/B _21261_/A _20735_/D vssd1 vssd1 vccd1 vccd1 _20857_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_136_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20666_ _20788_/A _20665_/B _20665_/C vssd1 vssd1 vccd1 vccd1 _20667_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__11559__A2 _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20597_ _20597_/A _20597_/B vssd1 vssd1 vccd1 vccd1 _20598_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18281__A _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16498__A2 _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17724__A1_N _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12020_ _12020_/A _12326_/D _12302_/A _12312_/A vssd1 vssd1 vccd1 vccd1 _12118_/A
+ sky130_fd_sc_hd__and4_1
X_21218_ _21218_/A _21218_/B vssd1 vssd1 vccd1 vccd1 _21220_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11192__A0 _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17998__A2 _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11731__A2 _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21149_ _21033_/A _21033_/B _20913_/Y vssd1 vssd1 vccd1 vccd1 _21259_/A sky130_fd_sc_hd__a21boi_4
Xfanout550 _21733_/Q vssd1 vssd1 vccd1 vccd1 _13860_/A sky130_fd_sc_hd__clkbuf_8
Xfanout561 _12621_/C vssd1 vssd1 vccd1 vccd1 _12214_/C sky130_fd_sc_hd__clkbuf_8
Xfanout572 _12268_/B vssd1 vssd1 vccd1 vccd1 _12402_/A sky130_fd_sc_hd__buf_4
XANTENNA__20689__C _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13971_ _14291_/A _13967_/B _14290_/B vssd1 vssd1 vccd1 vccd1 _14126_/A sky130_fd_sc_hd__o21ba_2
Xfanout583 _13985_/A vssd1 vssd1 vccd1 vccd1 _13394_/A sky130_fd_sc_hd__buf_4
Xfanout594 _11122_/A vssd1 vssd1 vccd1 vccd1 _11349_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__19262__D _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15710_ _15712_/B vssd1 vssd1 vccd1 vccd1 _15711_/B sky130_fd_sc_hd__inv_2
X_12922_ _12921_/A _12921_/B _12921_/C vssd1 vssd1 vccd1 vccd1 _12924_/C sky130_fd_sc_hd__a21o_1
X_16690_ _17141_/A _17433_/A _17526_/B _17141_/B vssd1 vssd1 vccd1 vccd1 _16691_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11495__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17063__C _17063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15641_ _15641_/A _15641_/B vssd1 vssd1 vccd1 vccd1 _15643_/B sky130_fd_sc_hd__xnor2_4
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12853_ _12853_/A _12853_/B vssd1 vssd1 vccd1 vccd1 _12855_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_115_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11247__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18360_ _18360_/A _18360_/B _18360_/C vssd1 vssd1 vccd1 vccd1 _18363_/B sky130_fd_sc_hd__nand3_4
X_11804_ _11776_/X _11777_/Y _11801_/A _11800_/Y vssd1 vssd1 vccd1 vccd1 _11805_/C
+ sky130_fd_sc_hd__a211o_1
X_15572_ _21740_/Q _15838_/D _16084_/C _16084_/D vssd1 vssd1 vccd1 vccd1 _15700_/A
+ sky130_fd_sc_hd__and4_1
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ _12784_/A _14384_/C vssd1 vssd1 vccd1 vccd1 _12787_/A sky130_fd_sc_hd__and2_1
XFILLER_0_95_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17311_ _17619_/A _17206_/B _17209_/B _17207_/X vssd1 vssd1 vccd1 vccd1 _17313_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__19372__A1 _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14523_ _14370_/A _14370_/C _14370_/B vssd1 vssd1 vccd1 vccd1 _14524_/C sky130_fd_sc_hd__a21bo_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19372__B2 _19531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18291_ _18292_/A _18292_/B vssd1 vssd1 vccd1 vccd1 _18414_/B sky130_fd_sc_hd__nand2b_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11735_ _11734_/A _11734_/B _11734_/C vssd1 vssd1 vccd1 vccd1 _11736_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_154_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17242_ _16608_/A _16608_/C _16608_/B vssd1 vssd1 vccd1 vccd1 _17243_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14454_ _14341_/A _14341_/B _14339_/Y vssd1 vssd1 vccd1 vccd1 _14496_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_3_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11666_ _11666_/A _11666_/B vssd1 vssd1 vccd1 vccd1 _12316_/B sky130_fd_sc_hd__nand2_1
X_13405_ _13405_/A _13405_/B vssd1 vssd1 vccd1 vccd1 _13415_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_272 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17173_ _21142_/A _17173_/B vssd1 vssd1 vccd1 vccd1 _17173_/Y sky130_fd_sc_hd__nor2_1
X_14385_ _14385_/A _14385_/B vssd1 vssd1 vccd1 vccd1 _14387_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_84_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11597_ _12426_/B _12402_/A vssd1 vssd1 vccd1 vccd1 _11874_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_109_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16124_ _16120_/A _16121_/Y _15944_/Y _15948_/B vssd1 vssd1 vccd1 vccd1 _16124_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_40_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13336_ _13335_/A _13335_/B _13335_/C vssd1 vssd1 vccd1 vccd1 _13338_/C sky130_fd_sc_hd__a21o_1
XANTENNA__18622__C _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_938 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16055_ _16226_/B _16055_/B vssd1 vssd1 vccd1 vccd1 _16070_/A sky130_fd_sc_hd__and2_1
X_13267_ _13267_/A _13267_/B vssd1 vssd1 vccd1 vccd1 _13275_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_122_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17238__C _17557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15006_ _15006_/A _15006_/B _15006_/C vssd1 vssd1 vccd1 vccd1 _15006_/X sky130_fd_sc_hd__and3_2
XANTENNA__12670__C _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12218_ _12217_/B _12217_/C _12217_/A vssd1 vssd1 vccd1 vccd1 _12219_/C sky130_fd_sc_hd__o21bai_1
XANTENNA__11183__A0 _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13198_ _13199_/A _13199_/B _13199_/C vssd1 vssd1 vccd1 vccd1 _13198_/X sky130_fd_sc_hd__and3_1
X_19814_ _19814_/A _19814_/B vssd1 vssd1 vccd1 vccd1 _19816_/A sky130_fd_sc_hd__xnor2_2
X_12149_ _12148_/B _12148_/C _12148_/A vssd1 vssd1 vccd1 vccd1 _12150_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__14878__B _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16661__A2 _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19745_ _20101_/B _19868_/B _19866_/C _20101_/A vssd1 vssd1 vccd1 vccd1 _19745_/X
+ sky130_fd_sc_hd__a22o_1
X_16957_ _16903_/A _16903_/C _16903_/B vssd1 vssd1 vccd1 vccd1 _16958_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14672__A1 _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14672__B2 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15908_ _15907_/A _15907_/B _15907_/C vssd1 vssd1 vccd1 vccd1 _15909_/B sky130_fd_sc_hd__o21a_1
XANTENNA__11486__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19676_ _19676_/A _19676_/B vssd1 vssd1 vccd1 vccd1 _19678_/B sky130_fd_sc_hd__nor2_1
X_16888_ _16888_/A _16888_/B vssd1 vssd1 vccd1 vccd1 _16890_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17610__A1 _19337_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17610__B2 _18851_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18627_ _18628_/A _18628_/B vssd1 vssd1 vccd1 vccd1 _18627_/Y sky130_fd_sc_hd__nand2b_1
X_15839_ _15838_/D _15838_/B _10797_/Y _14659_/A vssd1 vssd1 vccd1 vccd1 _15841_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11238__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11238__B2 _11459_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18558_ _18555_/X _18709_/B _18429_/D _18430_/B vssd1 vssd1 vccd1 vccd1 _18559_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17509_ _17510_/A _17510_/B vssd1 vssd1 vccd1 vccd1 _17629_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21170__A1 _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18489_ _18489_/A _18489_/B vssd1 vssd1 vccd1 vccd1 _18491_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_145_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_13 _11331_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12845__C _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20520_ _20774_/A _20774_/B _21258_/B _21171_/B vssd1 vssd1 vccd1 vccd1 _20686_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_145_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_24 _11339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_35 _11430_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_46 hold247/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_57 hold270/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20451_ _20450_/B _20450_/C _20450_/A vssd1 vssd1 vccd1 vccd1 _20451_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA_68 hold268/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_79 hold277/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout124_A _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11410__A1 _21293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20382_ _20788_/A _21146_/B vssd1 vssd1 vccd1 vccd1 _21034_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20136__A _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15152__A2 _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22052_ _22063_/CLK _22052_/D vssd1 vssd1 vccd1 vccd1 hold275/A sky130_fd_sc_hd__dfxtp_4
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11174__A0 _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout493_A _21746_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21003_ _21005_/B vssd1 vssd1 vccd1 vccd1 _21003_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16987__C _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11477__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21905_ _21938_/CLK hold127/X vssd1 vssd1 vccd1 vccd1 hold126/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11229__A1 _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11229__B2 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21836_ _21837_/CLK _21836_/D vssd1 vssd1 vccd1 vccd1 _21836_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout37_A _21490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21767_ _21767_/CLK _21767_/D vssd1 vssd1 vccd1 vccd1 _21767_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11520_ _11224_/A t2x[23] v1z[23] fanout21/X _11519_/X vssd1 vssd1 vccd1 vccd1 _11520_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15915__A1 _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20718_ _20718_/A _20843_/B vssd1 vssd1 vccd1 vccd1 _20720_/A sky130_fd_sc_hd__or2_2
XFILLER_0_0_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15915__B2 _16380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21698_ _22080_/CLK _21698_/D vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout3_A fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11451_ _11549_/A t2x[0] v1z[0] fanout17/X _11450_/X vssd1 vssd1 vccd1 vccd1 _11451_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20649_ _20650_/A _20650_/B vssd1 vssd1 vccd1 vccd1 _20916_/A sky130_fd_sc_hd__and2_1
XFILLER_0_135_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14170_ _14303_/B _14170_/B vssd1 vssd1 vccd1 vccd1 _14171_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11401__A1 _17334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13867__B _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11382_ hold308/X fanout29/X _11381_/X vssd1 vssd1 vccd1 vccd1 _11382_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12771__B _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20046__A _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19257__D _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13121_ _13121_/A _13121_/B _13121_/C vssd1 vssd1 vccd1 vccd1 _13124_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_108_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13052_ _13051_/B _13051_/C _13051_/A vssd1 vssd1 vccd1 vccd1 _13054_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11165__A0 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14979__A _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12003_ _12003_/A _12003_/B vssd1 vssd1 vccd1 vccd1 _12009_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17860_ _19337_/D _19060_/B vssd1 vssd1 vccd1 vccd1 _17864_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_100_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14698__B _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16811_ _16810_/A _16810_/C _16810_/B vssd1 vssd1 vccd1 vccd1 _16823_/B sky130_fd_sc_hd__a21o_1
X_17791_ _21824_/Q _20270_/C vssd1 vssd1 vccd1 vccd1 _17794_/A sky130_fd_sc_hd__and2_1
XANTENNA__13457__A2 _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout380 _21774_/Q vssd1 vssd1 vccd1 vccd1 _14828_/B sky130_fd_sc_hd__buf_4
XFILLER_0_75_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout391 _21771_/Q vssd1 vssd1 vccd1 vccd1 _13152_/D sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11468__A1 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19530_ _21278_/A _19529_/X _19528_/X vssd1 vssd1 vccd1 vccd1 _19532_/A sky130_fd_sc_hd__a21bo_1
X_13954_ _13802_/Y _13804_/X _13952_/Y _13953_/X vssd1 vssd1 vccd1 vccd1 _13956_/B
+ sky130_fd_sc_hd__a211oi_4
X_16742_ _16741_/A _16741_/C _16741_/B vssd1 vssd1 vccd1 vccd1 _16754_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11468__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12905_ _14716_/A _13034_/D vssd1 vssd1 vccd1 vccd1 _12909_/A sky130_fd_sc_hd__nand2_1
X_16673_ _16672_/A _16672_/C _16672_/B vssd1 vssd1 vccd1 vccd1 _16676_/B sky130_fd_sc_hd__a21o_1
X_19461_ _19461_/A _19461_/B vssd1 vssd1 vccd1 vccd1 _19464_/A sky130_fd_sc_hd__xor2_1
X_13885_ _13884_/B _13884_/C _13884_/A vssd1 vssd1 vccd1 vccd1 _13885_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_115_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18412_ _18414_/A _18414_/B _18414_/C vssd1 vssd1 vccd1 vccd1 _18413_/A sky130_fd_sc_hd__a21oi_2
X_15624_ _15622_/Y _15624_/B vssd1 vssd1 vccd1 vccd1 _15626_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_69_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12836_ _12837_/A _12837_/B _12837_/C vssd1 vssd1 vccd1 vccd1 _13083_/A sky130_fd_sc_hd__o21ai_2
X_19392_ _19692_/A _20148_/C _19392_/C _19543_/A vssd1 vssd1 vccd1 vccd1 _19543_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16418__B _16418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15555_ _15556_/B _15556_/A vssd1 vssd1 vccd1 vccd1 _15682_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__16159__A1 _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18343_ _18343_/A _18343_/B vssd1 vssd1 vccd1 vccd1 _18363_/A sky130_fd_sc_hd__xor2_2
XANTENNA__11850__B _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21152__A1 _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21043__C _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18336__D _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12767_ _12648_/X _12650_/X _12765_/X _12766_/Y vssd1 vssd1 vccd1 vccd1 _12803_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16159__B2 _16380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14506_ _14508_/A _15022_/B _14508_/C _14508_/D vssd1 vssd1 vccd1 vccd1 _14506_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18274_ _18275_/B _18275_/A vssd1 vssd1 vccd1 vccd1 _18398_/A sky130_fd_sc_hd__and2b_1
X_11718_ _11718_/A _11718_/B vssd1 vssd1 vccd1 vccd1 _11753_/A sky130_fd_sc_hd__xor2_2
X_15486_ _15487_/A _15487_/B vssd1 vssd1 vccd1 vccd1 _15486_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_84_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12698_ _12716_/B _12697_/B _12697_/C _12697_/D vssd1 vssd1 vccd1 vccd1 _12698_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_126_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21340__A _21349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14437_ _14438_/B _14438_/A vssd1 vssd1 vccd1 vccd1 _14437_/X sky130_fd_sc_hd__and2b_1
X_17225_ _17433_/A _19430_/A _17324_/D _17417_/A vssd1 vssd1 vccd1 vccd1 _17226_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11649_ _11649_/A _11649_/B vssd1 vssd1 vccd1 vccd1 _11650_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__15976__C _16396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12196__A2 _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17156_ _17156_/A _17156_/B _17156_/C vssd1 vssd1 vccd1 vccd1 _17159_/C sky130_fd_sc_hd__and3_1
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14368_ _14368_/A _14368_/B _14513_/B vssd1 vssd1 vccd1 vccd1 _14370_/B sky130_fd_sc_hd__nand3_1
XANTENNA__18856__B1 _19185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_136 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15695__D _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16107_ _16212_/A _21784_/Q _16196_/B _16107_/D vssd1 vssd1 vccd1 vccd1 _16212_/B
+ sky130_fd_sc_hd__and4b_1
X_13319_ _14716_/A _14384_/D vssd1 vssd1 vccd1 vccd1 _13323_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17087_ _17145_/A _17145_/B vssd1 vssd1 vccd1 vccd1 _17089_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_150_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14299_ hold157/X _14298_/X fanout4/X vssd1 vssd1 vccd1 vccd1 _21869_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_40_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16038_ _16038_/A _16038_/B vssd1 vssd1 vccd1 vccd1 _16079_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11156__A0 _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20106__D _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20415__B1 _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_110_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17989_ _17989_/A _17989_/B vssd1 vssd1 vccd1 vccd1 _17990_/B sky130_fd_sc_hd__xor2_2
XANTENNA__11459__A1 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19728_ _19847_/B _19844_/C _19847_/A _19592_/X vssd1 vssd1 vccd1 vccd1 _19740_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11459__B2 _11459_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13017__B _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19659_ _19659_/A _19659_/B vssd1 vssd1 vccd1 vccd1 _19679_/A sky130_fd_sc_hd__or2_1
XFILLER_0_79_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15513__A _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16328__B _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21621_ _21939_/CLK _21621_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[84] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14774__D _14774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout241_A _21293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21143__B2 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11252__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout339_A _21784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21552_ mstream_o[15] hold106/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22079_/D sky130_fd_sc_hd__mux2_1
XANTENNA__11631__A1 _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20792__C _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20503_ _20351_/Y _20353_/X _20501_/Y _20502_/X vssd1 vssd1 vccd1 vccd1 _20503_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_8_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21483_ hold181/X sstream_i[60] _21507_/S vssd1 vssd1 vccd1 vccd1 _22010_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_16_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16570__A1 _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout506_A _21743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16570__B2 _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12187__A2 _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20434_ _20434_/A _20558_/B vssd1 vssd1 vccd1 vccd1 _20436_/B sky130_fd_sc_hd__or2_1
XFILLER_0_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11934__A2 _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20365_ _20366_/A _20366_/B vssd1 vssd1 vccd1 vccd1 _20367_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_144_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22104_ _22105_/CLK _22104_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[40] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_101_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11147__A0 _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20296_ _20449_/A _20295_/C _20295_/A vssd1 vssd1 vccd1 vccd1 _20296_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_2_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22035_ _22038_/CLK _22035_/D vssd1 vssd1 vccd1 vccd1 hold280/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_hold286_A hold286/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17606__C _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14949__D _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14636__A1 _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20032__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19390__A _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10951_ mstream_o[57] _10950_/Y _10992_/S vssd1 vssd1 vccd1 vccd1 _21594_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_74_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21382__A1 _19476_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16519__A _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13670_ _14133_/D _16399_/B _16409_/B _13983_/B vssd1 vssd1 vccd1 vccd1 _13670_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10882_ mstream_o[47] _10881_/X _10992_/S vssd1 vssd1 vccd1 vccd1 _21584_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_112_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12621_ _12732_/A _12620_/Y _12621_/C _13573_/D vssd1 vssd1 vccd1 vccd1 _12732_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_109_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21819_ _21821_/CLK _21819_/D vssd1 vssd1 vccd1 vccd1 hold264/A sky130_fd_sc_hd__dfxtp_2
XFILLER_0_38_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18734__A _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11162__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15340_ _15340_/A _15340_/B vssd1 vssd1 vccd1 vccd1 _15342_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_65_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12552_ _13157_/A _12897_/C _12897_/D _13017_/A vssd1 vssd1 vccd1 vccd1 _12553_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_136_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14981__B _21755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11503_ _11502_/X _19240_/B _11521_/S vssd1 vssd1 vccd1 vccd1 _21839_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15271_ _15271_/A _15271_/B vssd1 vssd1 vccd1 vccd1 _15281_/A sky130_fd_sc_hd__or2_2
XFILLER_0_136_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12483_ _12479_/Y _12480_/X _12379_/B _12379_/Y vssd1 vssd1 vccd1 vccd1 _12484_/C
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17010_ _16994_/A _16994_/C _16994_/B vssd1 vssd1 vccd1 vccd1 _17010_/X sky130_fd_sc_hd__o21a_1
X_14222_ _14222_/A _14222_/B _14222_/C vssd1 vssd1 vccd1 vccd1 _14224_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18172__C _19379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11434_ _11433_/X _21046_/B _11470_/S vssd1 vssd1 vccd1 vccd1 _21816_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_105_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14153_ _14153_/A _14153_/B vssd1 vssd1 vccd1 vccd1 _14160_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16313__A1 _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11365_ _11364_/X _17123_/C _11401_/S vssd1 vssd1 vccd1 vccd1 _21793_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_46_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13104_ _13104_/A _13104_/B _13104_/C vssd1 vssd1 vccd1 vccd1 _13250_/C sky130_fd_sc_hd__nand3_2
X_14084_ _14572_/A _14713_/A _15234_/C vssd1 vssd1 vccd1 vccd1 _14084_/X sky130_fd_sc_hd__and3_1
XANTENNA__11138__A0 _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18961_ _19123_/B _21171_/B vssd1 vssd1 vccd1 vccd1 _18964_/A sky130_fd_sc_hd__nand2_1
X_11296_ _12402_/B _11295_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21775_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14875__A1 _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14875__B2 _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ _13173_/C _15076_/B _13034_/D _15076_/A vssd1 vssd1 vccd1 vccd1 _13036_/D
+ sky130_fd_sc_hd__a22o_1
X_17912_ _17912_/A _17912_/B vssd1 vssd1 vccd1 vccd1 _17948_/A sky130_fd_sc_hd__nand2_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11689__A1 _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18892_ _19051_/A _20026_/B _19060_/B _19051_/C vssd1 vssd1 vccd1 vccd1 _18894_/D
+ sky130_fd_sc_hd__nand4_4
XANTENNA__11689__B2 _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17843_ _17720_/X _17725_/A _18703_/A _19030_/C vssd1 vssd1 vccd1 vccd1 _18121_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18909__A _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_7_clk_i _21806_/CLK vssd1 vssd1 vccd1 vccd1 _21816_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_156_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13118__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17774_ _17647_/X _17649_/X _17772_/Y _17773_/X vssd1 vssd1 vccd1 vccd1 _17776_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11564__C _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14986_ _15085_/A _15502_/A _14984_/Y _14985_/X vssd1 vssd1 vccd1 vccd1 _14990_/A
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_135_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19513_ _19512_/B _19512_/C _19512_/A vssd1 vssd1 vccd1 vccd1 _19514_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_92_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16725_ _17145_/A _16860_/C vssd1 vssd1 vccd1 vccd1 _16727_/B sky130_fd_sc_hd__and2_1
X_13937_ _13936_/A _13936_/B _13936_/C vssd1 vssd1 vccd1 vccd1 _13939_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_152_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19444_ _19444_/A _19444_/B vssd1 vssd1 vccd1 vccd1 _19448_/A sky130_fd_sc_hd__nor2_2
X_13868_ _13710_/X _13713_/B _13865_/X _13867_/Y vssd1 vssd1 vccd1 vccd1 _13868_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_278 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16656_ _17178_/B _16657_/B _16657_/C _16657_/D vssd1 vssd1 vccd1 vccd1 _16656_/Y
+ sky130_fd_sc_hd__nor4_2
XANTENNA__11861__A1 _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11861__B2 _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15607_ _15422_/X _15426_/C _15693_/B _15606_/Y vssd1 vssd1 vccd1 vccd1 _15607_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11580__B _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ _12818_/B _12818_/C _12818_/A vssd1 vssd1 vccd1 vccd1 _12947_/C sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19375_ _19664_/B _20671_/B vssd1 vssd1 vccd1 vccd1 _19376_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_146_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13799_ _13800_/A _13800_/B _13800_/C _13800_/D vssd1 vssd1 vccd1 vccd1 _13799_/Y
+ sky130_fd_sc_hd__nor4_1
X_16587_ _21825_/Q _16734_/B _17434_/B _17433_/A vssd1 vssd1 vccd1 vccd1 _16590_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_60_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18326_ _18326_/A _18326_/B vssd1 vssd1 vccd1 vccd1 _18328_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15538_ _16369_/A _16399_/A _15539_/C _15539_/D vssd1 vssd1 vccd1 vccd1 _15540_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_84_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15469_ _15469_/A _15469_/B _15469_/C vssd1 vssd1 vccd1 vccd1 _15469_/Y sky130_fd_sc_hd__nor3_2
X_18257_ _18857_/B _19201_/B _18255_/Y _18402_/A vssd1 vssd1 vccd1 vccd1 _18259_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_71_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17208_ _17520_/A _17417_/C _17417_/D _17520_/B vssd1 vssd1 vccd1 vccd1 _17209_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18188_ _18787_/A _18787_/B _18773_/B _19546_/D vssd1 vssd1 vccd1 vccd1 _18332_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_130_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12842__D _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16314__D _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17139_ _17145_/A _17146_/C _17126_/C _17126_/D vssd1 vssd1 vccd1 vccd1 _17140_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__16304__B2 _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20100__A2 _21816_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19906__C _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20150_ _20151_/A _20151_/B vssd1 vssd1 vccd1 vccd1 _20294_/A sky130_fd_sc_hd__or2_1
XFILLER_0_69_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11129__A0 _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_976 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16611__B _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15508__A _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20081_ _20081_/A _20081_/B vssd1 vssd1 vccd1 vccd1 _20081_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20939__A1 _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20133__B _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16607__A2 _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout191_A _17557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout289_A _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17280__A2 _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18538__B _21364_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17442__B _18058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20983_ _20983_/A _20983_/B vssd1 vssd1 vccd1 vccd1 _20984_/B sky130_fd_sc_hd__and2_1
XFILLER_0_95_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11852__A1 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_259 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout623_A _17557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18554__A _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11921__D _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21604_ _21934_/CLK _21604_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[67] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21535_ hold277/X sstream_i[112] _21536_/S vssd1 vssd1 vccd1 vccd1 _22062_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_129_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17740__B1 _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21466_ hold211/X sstream_i[43] _21494_/S vssd1 vssd1 vccd1 vccd1 _21993_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_121_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14306__B _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20417_ _20552_/A vssd1 vssd1 vccd1 vccd1 _20419_/D sky130_fd_sc_hd__inv_2
X_21397_ _21720_/D _15356_/X _21396_/Y vssd1 vssd1 vccd1 vccd1 _21397_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16802__A _16870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12107__A _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _12639_/A _11149_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21733_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_113_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20348_ _20348_/A _20498_/A _20348_/C vssd1 vssd1 vccd1 vccd1 _20498_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_144_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19535__D _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11081_ _10946_/Y hold71/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21676_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13864__C _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20279_ _20279_/A _20279_/B vssd1 vssd1 vccd1 vccd1 _20280_/B sky130_fd_sc_hd__nand2_1
X_22018_ _22020_/CLK _22018_/D vssd1 vssd1 vccd1 vccd1 hold165/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14840_ _14840_/A _14840_/B _14840_/C vssd1 vssd1 vccd1 vccd1 _14840_/Y sky130_fd_sc_hd__nand3_1
X_14771_ _14771_/A _14771_/B vssd1 vssd1 vccd1 vccd1 _14773_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__13293__B1 _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11983_ _12261_/A _12269_/B _12751_/B _12637_/B vssd1 vssd1 vccd1 vccd1 _11986_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__15153__A _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13722_ _13875_/B _13877_/A _14516_/A _14365_/C vssd1 vssd1 vccd1 vccd1 _13724_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_98_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16510_ _17029_/A _16860_/C _16917_/C _16743_/B vssd1 vssd1 vccd1 vccd1 _16512_/C
+ sky130_fd_sc_hd__a22o_1
X_10934_ _10940_/B _10934_/B vssd1 vssd1 vccd1 vccd1 _10934_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17490_ _17490_/A _21792_/Q _20797_/A _21258_/A vssd1 vssd1 vccd1 vccd1 _17614_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_98_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13653_ _13652_/A _13652_/B _13652_/C _13652_/D vssd1 vssd1 vccd1 vccd1 _13653_/X
+ sky130_fd_sc_hd__o22a_1
X_16441_ _16868_/A _16734_/B _17223_/A _16860_/C vssd1 vssd1 vccd1 vccd1 _16444_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__13045__B1 _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10865_ _10866_/A _10866_/B _10864_/Y vssd1 vssd1 vccd1 vccd1 _10873_/B sky130_fd_sc_hd__o21bai_2
XANTENNA__18464__A _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12604_ _12604_/A _12604_/B vssd1 vssd1 vccd1 vccd1 _12606_/B sky130_fd_sc_hd__nor2_1
X_16372_ _16372_/A _16372_/B vssd1 vssd1 vccd1 vccd1 _16373_/B sky130_fd_sc_hd__xnor2_2
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19160_ _18995_/A _19160_/B vssd1 vssd1 vccd1 vccd1 _19162_/B sky130_fd_sc_hd__and2b_1
X_13584_ _13581_/Y _13582_/X _13450_/X _13453_/Y vssd1 vssd1 vccd1 vccd1 _13584_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_82_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10796_ _21171_/A vssd1 vssd1 vccd1 vccd1 _10796_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_82_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19279__B _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15323_ _15324_/A _15324_/B vssd1 vssd1 vccd1 vccd1 _15323_/X sky130_fd_sc_hd__or2_1
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18111_ _19008_/D _19199_/C _19199_/D _21791_/Q vssd1 vssd1 vccd1 vccd1 _18111_/Y
+ sky130_fd_sc_hd__a22oi_1
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12535_ _12877_/A _13155_/C _13155_/D _12642_/A vssd1 vssd1 vccd1 vccd1 _12536_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19091_ _19092_/B _19092_/C _19262_/C _19092_/A vssd1 vssd1 vccd1 vccd1 _19095_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15254_ _15254_/A _15254_/B vssd1 vssd1 vccd1 vccd1 _15288_/A sky130_fd_sc_hd__nor2_1
X_18042_ _18042_/A _18164_/B _18042_/C vssd1 vssd1 vccd1 vccd1 _18044_/B sky130_fd_sc_hd__nand3_2
X_12466_ _12465_/B _12465_/C _12465_/A vssd1 vssd1 vccd1 vccd1 _12468_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_124_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14205_ _14070_/B _14072_/A _14203_/X _14204_/Y vssd1 vssd1 vccd1 vccd1 _14207_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__18911__B _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11417_ _11447_/A1 hold302/A fanout47/X hold131/A vssd1 vssd1 vccd1 vccd1 _11417_/X
+ sky130_fd_sc_hd__a22o_1
X_15185_ _15185_/A _15296_/A _15185_/C vssd1 vssd1 vccd1 vccd1 _15296_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_50_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12397_ _13983_/B _13394_/A _13258_/C _13258_/D vssd1 vssd1 vccd1 vccd1 _12398_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_151_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14136_ _14136_/A vssd1 vssd1 vccd1 vccd1 _14146_/A sky130_fd_sc_hd__inv_2
X_11348_ _15838_/B _11347_/X _11348_/S vssd1 vssd1 vccd1 vccd1 _21788_/D sky130_fd_sc_hd__mux2_1
X_19993_ _20416_/A _21291_/A _20416_/B _20273_/A vssd1 vssd1 vccd1 vccd1 _20138_/A
+ sky130_fd_sc_hd__nand4_2
X_14067_ _14209_/A _14066_/C _14066_/A vssd1 vssd1 vccd1 vccd1 _14068_/C sky130_fd_sc_hd__a21o_1
X_18944_ _18944_/A _18944_/B _18944_/C vssd1 vssd1 vccd1 vccd1 _18946_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_123_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11279_ fanout58/X v0z[13] fanout17/X _11278_/X vssd1 vssd1 vccd1 vccd1 _11279_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13018_ _13155_/B _13018_/B _13155_/C _21768_/Q vssd1 vssd1 vccd1 vccd1 _13020_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_20_1114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12323__A2 _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11575__B _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18875_ _18874_/B _19028_/B _18874_/A vssd1 vssd1 vccd1 vccd1 _18876_/C sky130_fd_sc_hd__a21o_1
XANTENNA__11067__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17826_ _17704_/A _17704_/B _17702_/X vssd1 vssd1 vccd1 vccd1 _17828_/B sky130_fd_sc_hd__o21a_1
XANTENNA__17543__A _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15273__A1 _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14076__A2 _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15273__B2 _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17757_ _18008_/B _18769_/B vssd1 vssd1 vccd1 vccd1 _17761_/A sky130_fd_sc_hd__nand2_1
X_14969_ _14970_/A _14970_/B vssd1 vssd1 vccd1 vccd1 _14969_/X sky130_fd_sc_hd__and2b_1
X_16708_ _16712_/B vssd1 vssd1 vccd1 vccd1 _16708_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_18_1043 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17688_ _17689_/A _17689_/B _17689_/C _17689_/D vssd1 vssd1 vccd1 vccd1 _17688_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_147_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19427_ _19427_/A _19427_/B vssd1 vssd1 vccd1 vccd1 _19436_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_58_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16639_ _16639_/A _16639_/B _16639_/C vssd1 vssd1 vccd1 vccd1 _16665_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout19 _11224_/Y vssd1 vssd1 vccd1 vccd1 fanout19/X sky130_fd_sc_hd__buf_4
XFILLER_0_29_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19358_ _19347_/Y _19358_/B _19358_/C vssd1 vssd1 vccd1 vccd1 _19519_/A sky130_fd_sc_hd__and3b_1
XANTENNA__11598__B1 _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16606__B _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18309_ _18157_/A _18157_/Y _18307_/X _18308_/Y vssd1 vssd1 vccd1 vccd1 _18373_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19289_ _19289_/A _19289_/B vssd1 vssd1 vccd1 vccd1 _19292_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_72_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11530__S _11545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20128__B _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13311__A _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21320_ _21320_/A _21320_/B vssd1 vssd1 vccd1 vccd1 _21321_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18278__A1 _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21251_ hold195/A _11551_/Y fanout1/X vssd1 vssd1 vccd1 vccd1 _21251_/X sky130_fd_sc_hd__o21a_1
XANTENNA__18278__B2 _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout204_A _21817_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20202_ _20202_/A _20202_/B vssd1 vssd1 vccd1 vccd1 _20205_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21182_ _21182_/A _21182_/B vssd1 vssd1 vccd1 vccd1 _21183_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20133_ _20416_/A _20416_/B _20273_/A _20270_/C vssd1 vssd1 vccd1 vccd1 _20275_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_99_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20064_ _20216_/A _20062_/X _19837_/A _19838_/X vssd1 vssd1 vccd1 vccd1 _20065_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout573_A _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17172__B _21331_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_306 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_317 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_328 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_339 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20966_ _21199_/A _21293_/A _21286_/B _21296_/B vssd1 vssd1 vccd1 vccd1 _21085_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_36_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20897_ _20898_/A _20898_/B vssd1 vssd1 vccd1 vccd1 _21138_/A sky130_fd_sc_hd__and2b_1
XANTENNA__20560__A2 _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19702__A1 _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19702__B2 _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18434__D _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11440__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ _12401_/A vssd1 vssd1 vccd1 vccd1 _12320_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_133_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21518_ hold251/X sstream_i[95] _21528_/S vssd1 vssd1 vccd1 vccd1 _22045_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_90_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12251_ _12267_/A _12269_/C _12269_/D _12242_/B vssd1 vssd1 vccd1 vccd1 _12252_/B
+ sky130_fd_sc_hd__a22oi_1
X_21449_ hold119/X sstream_i[26] _21481_/S vssd1 vssd1 vccd1 vccd1 _21976_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_142_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11202_ hold293/X fanout51/X fanout48/X hold228/X vssd1 vssd1 vccd1 vccd1 _11202_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13875__B _13875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12182_ _12269_/A _12512_/A _12214_/C _12245_/B vssd1 vssd1 vccd1 vccd1 _12183_/C
+ sky130_fd_sc_hd__a22o_1
X_11133_ hold222/X _11126_/A _11126_/B hold176/X vssd1 vssd1 vccd1 vccd1 _11133_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17492__A2 _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13594__C _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16990_ _16990_/A _17033_/A vssd1 vssd1 vccd1 vccd1 _16992_/B sky130_fd_sc_hd__nor2_1
XANTENNA__20989__A _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15941_ _15941_/A _16078_/A _15941_/C vssd1 vssd1 vccd1 vccd1 _15942_/A sky130_fd_sc_hd__and3_2
X_11064_ _11063_/X hold25/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21661_/D sky130_fd_sc_hd__mux2_1
XANTENNA__21576__A1 _11059_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18660_ _18505_/A _18505_/C _18505_/B vssd1 vssd1 vccd1 vccd1 _18661_/C sky130_fd_sc_hd__a21bo_1
X_15872_ _15733_/B _15732_/Y _15870_/A _15871_/X vssd1 vssd1 vccd1 vccd1 _15874_/C
+ sky130_fd_sc_hd__o211a_2
XANTENNA__15255__B2 _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17611_ _17854_/B _21256_/A _17611_/C _17611_/D vssd1 vssd1 vccd1 vccd1 _17732_/B
+ sky130_fd_sc_hd__and4_1
X_14823_ _14821_/X _14823_/B vssd1 vssd1 vccd1 vccd1 _14824_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_153_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18591_ _18592_/A _18592_/B vssd1 vssd1 vccd1 vccd1 _18720_/B sky130_fd_sc_hd__or2_2
XTAP_3840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17542_ _21803_/Q _19432_/A vssd1 vssd1 vccd1 vccd1 _17546_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14754_ _14754_/A _14754_/B vssd1 vssd1 vccd1 vccd1 _14755_/B sky130_fd_sc_hd__xor2_4
X_11966_ _11944_/Y _11964_/X _11965_/Y _11892_/X vssd1 vssd1 vccd1 vccd1 _11971_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_54_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12300__A _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16204__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13705_ _13858_/B _13860_/A _13858_/C _16414_/A vssd1 vssd1 vccd1 vccd1 _13707_/D
+ sky130_fd_sc_hd__nand4_2
X_10917_ _10917_/A _10917_/B vssd1 vssd1 vccd1 vccd1 _10919_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14685_ _14809_/A _14684_/C _14684_/A vssd1 vssd1 vccd1 vccd1 _14685_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_10_clk_i _21806_/CLK vssd1 vssd1 vccd1 vccd1 _22013_/CLK sky130_fd_sc_hd__clkbuf_16
X_17473_ _17470_/X _17471_/X _17360_/C _17362_/A vssd1 vssd1 vccd1 vccd1 _17474_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_54_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11897_ _11897_/A _11897_/B vssd1 vssd1 vccd1 vccd1 _11899_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19212_ _19213_/A _19213_/B vssd1 vssd1 vccd1 vccd1 _19212_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_156_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16424_ _16424_/A _21784_/Q vssd1 vssd1 vccd1 vccd1 _16432_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_129_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13636_ _13635_/A _13635_/B _13635_/C vssd1 vssd1 vccd1 vccd1 _13638_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_39_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10848_ _10843_/A _10843_/B _10843_/C _11063_/B _11061_/A vssd1 vssd1 vccd1 vccd1
+ _11065_/C sky130_fd_sc_hd__a311o_1
XFILLER_0_39_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13560__A2_N _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20229__A _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19143_ _19143_/A _19143_/B _19143_/C vssd1 vssd1 vccd1 vccd1 _19143_/X sky130_fd_sc_hd__and3_1
XFILLER_0_66_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16355_ _16211_/A _16210_/Y _16209_/B vssd1 vssd1 vccd1 vccd1 _16356_/B sky130_fd_sc_hd__a21oi_2
X_13567_ _13567_/A _13567_/B vssd1 vssd1 vccd1 vccd1 _13568_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15235__A1_N _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15306_ _15306_/A _15437_/B _15307_/B vssd1 vssd1 vccd1 vccd1 _15306_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_87_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_25_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21934_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12518_ _12519_/A _12519_/B vssd1 vssd1 vccd1 vccd1 _12629_/B sky130_fd_sc_hd__nand2_1
X_16286_ _16286_/A _16286_/B _16286_/C _16286_/D vssd1 vssd1 vccd1 vccd1 _16287_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_125_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19074_ _19073_/B _19073_/C _19073_/A vssd1 vssd1 vccd1 vccd1 _19076_/B sky130_fd_sc_hd__a21o_1
X_13498_ _13348_/B _13347_/Y _13496_/X _13497_/Y vssd1 vssd1 vccd1 vccd1 _13500_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_14_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17180__A1 _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20845__A_N _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18025_ _18107_/A _18023_/X _17883_/B _17884_/Y vssd1 vssd1 vccd1 vccd1 _18087_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_23_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15237_ _15237_/A _15377_/B vssd1 vssd1 vccd1 vccd1 _15240_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12449_ _12449_/A _12449_/B vssd1 vssd1 vccd1 vccd1 _12451_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_152_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13741__A1 _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11347__A3 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15168_ _15028_/A _15027_/B _15025_/X vssd1 vssd1 vccd1 vccd1 _15179_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13741__B2 _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14119_ _13956_/B _13958_/A _14280_/B _14118_/Y vssd1 vssd1 vccd1 vccd1 _14121_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19753__A _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15099_ _14998_/X _15001_/X _15097_/X _15238_/B vssd1 vssd1 vccd1 vccd1 _15226_/A
+ sky130_fd_sc_hd__o211ai_4
Xfanout209 _21815_/Q vssd1 vssd1 vccd1 vccd1 _19753_/B sky130_fd_sc_hd__buf_4
X_19976_ _19973_/X _20110_/B _19871_/X _19874_/X vssd1 vssd1 vccd1 vccd1 _19977_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18927_ _20101_/B _19089_/B vssd1 vssd1 vccd1 vccd1 _18931_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_1012 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18858_ _18859_/A _21261_/B _18859_/C _18859_/D vssd1 vssd1 vccd1 vccd1 _18860_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_94_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20411__B _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17809_ _17810_/A _17810_/B _17810_/C vssd1 vssd1 vccd1 vccd1 _17809_/Y sky130_fd_sc_hd__nor3_1
X_18789_ _18789_/A _18789_/B _18789_/C _18947_/A vssd1 vssd1 vccd1 vccd1 _18947_/B
+ sky130_fd_sc_hd__nand4_1
X_20820_ _20951_/B _20820_/B vssd1 vssd1 vccd1 vccd1 _20823_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12848__C _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17720__B _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20751_ _20835_/B _20748_/Y _20574_/X _20578_/B vssd1 vssd1 vccd1 vccd1 _20751_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15549__A2 _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout154_A _21831_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15521__A _16031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20682_ _20683_/A _20683_/B vssd1 vssd1 vccd1 vccd1 _20872_/B sky130_fd_sc_hd__or2_1
XFILLER_0_58_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18499__A1 _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout321_A _21791_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11260__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout419_A _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21303_ _21303_/A _21303_/B vssd1 vssd1 vccd1 vccd1 _21309_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17448__A _17557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12535__A2 _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21234_ _21234_/A _21234_/B vssd1 vssd1 vccd1 vccd1 _21236_/C sky130_fd_sc_hd__xnor2_1
Xhold230 hold317/A vssd1 vssd1 vccd1 vccd1 hold230/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold241 hold241/A vssd1 vssd1 vccd1 vccd1 hold241/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 hold252/A vssd1 vssd1 vccd1 vccd1 hold252/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 hold263/A vssd1 vssd1 vccd1 vccd1 hold263/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold274 hold274/A vssd1 vssd1 vccd1 vccd1 hold274/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold285 hold285/A vssd1 vssd1 vccd1 vccd1 hold285/X sky130_fd_sc_hd__dlygate4sd3_1
X_21165_ _21172_/A _21062_/B _21065_/A vssd1 vssd1 vccd1 vccd1 _21176_/A sky130_fd_sc_hd__o21ai_1
Xhold296 hold296/A vssd1 vssd1 vccd1 vccd1 hold296/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20116_ _20116_/A _20116_/B vssd1 vssd1 vccd1 vccd1 _20119_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__19382__B _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12299__A1 _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21096_ _21096_/A _21096_/B vssd1 vssd1 vccd1 vccd1 _21107_/A sky130_fd_sc_hd__or2_1
XANTENNA__18279__A _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20047_ _20590_/D _20193_/D _20045_/Y _20188_/A vssd1 vssd1 vccd1 vccd1 _20049_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout67_A _19181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20230__B2 _11550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_103 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ _11819_/A _11819_/C _11819_/B vssd1 vssd1 vccd1 vccd1 _11823_/B sky130_fd_sc_hd__a21o_1
XTAP_3169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_114 sstream_i[67] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_125 v0z[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21998_ _22021_/CLK _21998_/D vssd1 vssd1 vccd1 vccd1 hold154/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_95_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_136 v1z[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20975__C _21853_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_147 v1z[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_158 v2z[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11751_ _11750_/A _11750_/B _11750_/C vssd1 vssd1 vccd1 vccd1 _11753_/C sky130_fd_sc_hd__a21o_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20949_ _20949_/A _20949_/B vssd1 vssd1 vccd1 vccd1 _20951_/C sky130_fd_sc_hd__xnor2_1
XANTENNA_169 v2z[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16527__A _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14470_ _14471_/A _14471_/B vssd1 vssd1 vccd1 vccd1 _14472_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_95_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11682_ _11682_/A _11705_/B _11682_/C vssd1 vssd1 vccd1 vccd1 _11685_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_48_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13421_ _13290_/D _13292_/A _13419_/X _13569_/B vssd1 vssd1 vccd1 vccd1 _13580_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_107_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13589__C _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_692 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20991__B _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16140_ _16251_/B _16138_/X _16007_/A _16009_/X vssd1 vssd1 vccd1 vccd1 _16142_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13352_ _13353_/A _13353_/B _13353_/C vssd1 vssd1 vccd1 vccd1 _13352_/X sky130_fd_sc_hd__and3_1
XANTENNA__12774__A2 _21766_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12303_ _13525_/A _12402_/B _12302_/C _12302_/D vssd1 vssd1 vccd1 vccd1 _12304_/B
+ sky130_fd_sc_hd__a22o_1
X_16071_ _16071_/A vssd1 vssd1 vccd1 vccd1 _16071_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_106_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13283_ _13280_/Y _13281_/X _13166_/B _13168_/A vssd1 vssd1 vccd1 vccd1 _13283_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_84_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15022_ _16084_/A _15022_/B vssd1 vssd1 vccd1 vccd1 _15024_/C sky130_fd_sc_hd__and2_1
XFILLER_0_121_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13723__A1 _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12234_ _12234_/A _12234_/B _12234_/C vssd1 vssd1 vccd1 vccd1 _12241_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_121_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18111__B1 _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19830_ _19830_/A _19830_/B _19830_/C vssd1 vssd1 vccd1 vccd1 _19830_/X sky130_fd_sc_hd__and3_1
X_12165_ _12165_/A _12165_/B vssd1 vssd1 vccd1 vccd1 _12168_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_124_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11116_ _10959_/Y hold12/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21710_/D sky130_fd_sc_hd__mux2_1
X_19761_ _19578_/B _19581_/B _19759_/A _19760_/Y vssd1 vssd1 vccd1 vccd1 _19763_/C
+ sky130_fd_sc_hd__a211o_2
X_16973_ _16973_/A _16973_/B _16973_/C vssd1 vssd1 vccd1 vccd1 _16980_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_21_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12096_ _12094_/X _12096_/B vssd1 vssd1 vccd1 vccd1 _12098_/A sky130_fd_sc_hd__and2b_1
XANTENNA__17093__A _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18712_ _19337_/D _19201_/B _18713_/C _18713_/D vssd1 vssd1 vccd1 vccd1 _18712_/Y
+ sky130_fd_sc_hd__a22oi_2
X_15924_ _15925_/A _15925_/B vssd1 vssd1 vccd1 vccd1 _16114_/B sky130_fd_sc_hd__or2_1
X_11047_ _11047_/A _11047_/B vssd1 vssd1 vccd1 vccd1 _11048_/B sky130_fd_sc_hd__nor2_2
X_19692_ _19692_/A _19692_/B _19692_/C _20416_/B vssd1 vssd1 vccd1 vccd1 _19695_/D
+ sky130_fd_sc_hd__nand4_1
XANTENNA__15228__A1 _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15228__B2 _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18643_ _18641_/X _18643_/B vssd1 vssd1 vccd1 vccd1 _18644_/B sky130_fd_sc_hd__and2b_1
X_15855_ _15855_/A _15972_/B vssd1 vssd1 vccd1 vccd1 _15857_/B sky130_fd_sc_hd__or2_1
XFILLER_0_87_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14806_ _14806_/A _14806_/B vssd1 vssd1 vccd1 vccd1 _14808_/B sky130_fd_sc_hd__xnor2_1
X_18574_ _18456_/X _18459_/Y _18571_/Y _18573_/X vssd1 vssd1 vccd1 vccd1 _18693_/A
+ sky130_fd_sc_hd__a211oi_2
XTAP_3670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15786_ _16328_/A _15911_/A _16424_/A _15911_/C vssd1 vssd1 vccd1 vccd1 _15973_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_87_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12998_ _12997_/B _12997_/C _12997_/A vssd1 vssd1 vccd1 vccd1 _13000_/B sky130_fd_sc_hd__a21o_1
XTAP_3692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17525_ _17525_/A _20249_/A vssd1 vssd1 vccd1 vccd1 _17529_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_54_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21343__A _21349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14737_ _14738_/A _14738_/B vssd1 vssd1 vccd1 vccd1 _14737_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_15_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11949_ _12020_/A _12326_/D _12402_/A _12302_/A vssd1 vssd1 vccd1 vccd1 _11953_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_143_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17456_ _17455_/B _17455_/C _17455_/A vssd1 vssd1 vccd1 vccd1 _17458_/B sky130_fd_sc_hd__a21o_1
X_14668_ _14664_/X _14666_/Y _14504_/X _14507_/X vssd1 vssd1 vccd1 vccd1 _14669_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16407_ _16407_/A _16407_/B vssd1 vssd1 vccd1 vccd1 _16408_/B sky130_fd_sc_hd__xnor2_1
X_13619_ _14848_/A _13913_/C vssd1 vssd1 vccd1 vccd1 _13623_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19748__A _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17387_ _17387_/A _21256_/A vssd1 vssd1 vccd1 vccd1 _17388_/B sky130_fd_sc_hd__nand2_1
X_14599_ _14599_/A _14599_/B vssd1 vssd1 vccd1 vccd1 _14911_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_82_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19126_ _19126_/A _19126_/B _19126_/C vssd1 vssd1 vccd1 vccd1 _19291_/A sky130_fd_sc_hd__and3_4
XFILLER_0_55_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16338_ _16225_/Y _16227_/Y _16388_/B _16337_/Y vssd1 vssd1 vccd1 vccd1 _16340_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19057_ _19686_/B _19529_/B _19057_/C _19057_/D vssd1 vssd1 vccd1 vccd1 _19060_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_140_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16269_ _16269_/A _16269_/B vssd1 vssd1 vccd1 vccd1 _16278_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_125_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18008_ _18008_/A _18008_/B _19906_/A _20146_/B vssd1 vssd1 vccd1 vccd1 _18144_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_51_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19959_ _19958_/B _19958_/C _19958_/A vssd1 vssd1 vccd1 vccd1 _19961_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__17434__C _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21921_ _21923_/CLK _21921_/D vssd1 vssd1 vccd1 vccd1 hold125/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout271_A _17417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout369_A _21777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13036__A _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14978__B1 _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21852_ _21853_/CLK _21852_/D vssd1 vssd1 vccd1 vccd1 hold321/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19905__A1 _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20803_ _20802_/A _20931_/B _20801_/X vssd1 vssd1 vccd1 vccd1 _20804_/B sky130_fd_sc_hd__o21bai_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19905__B2 _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12453__A1 _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21783_ _21821_/CLK _21783_/D vssd1 vssd1 vccd1 vccd1 _21783_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20515__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17916__B1 _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout536_A _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__B2 _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20734_ _21261_/A _21311_/B _20732_/Y _20857_/A vssd1 vssd1 vccd1 vccd1 _20736_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_9_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16195__A2 _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17392__A1 _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_93_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20665_ _20788_/A _20665_/B _20665_/C vssd1 vssd1 vccd1 vccd1 _20667_/A sky130_fd_sc_hd__or3_1
XFILLER_0_45_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20596_ _20597_/A _20597_/B vssd1 vssd1 vccd1 vccd1 _20596_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_34_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18281__B _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21217_ _21215_/Y _21217_/B vssd1 vssd1 vccd1 vccd1 _21218_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_143_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21148_ _21067_/A _21067_/B _21068_/X vssd1 vssd1 vccd1 vccd1 _21182_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__13469__B1 _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout540 _12637_/A vssd1 vssd1 vccd1 vccd1 _12751_/B sky130_fd_sc_hd__buf_4
Xfanout551 _21733_/Q vssd1 vssd1 vccd1 vccd1 _14936_/D sky130_fd_sc_hd__clkbuf_8
XANTENNA__15426__A _15426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout562 _14463_/D vssd1 vssd1 vccd1 vccd1 _13975_/B sky130_fd_sc_hd__buf_4
XANTENNA__20689__D _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13970_ hold133/X _13969_/X fanout2/X vssd1 vssd1 vccd1 vccd1 _21867_/D sky130_fd_sc_hd__mux2_1
X_21079_ _21291_/A _21286_/B _21296_/B _21293_/A vssd1 vssd1 vccd1 vccd1 _21083_/C
+ sky130_fd_sc_hd__a22o_1
Xfanout573 _14133_/D vssd1 vssd1 vccd1 vccd1 _13822_/B sky130_fd_sc_hd__buf_4
Xfanout584 _21726_/Q vssd1 vssd1 vccd1 vccd1 _13985_/A sky130_fd_sc_hd__buf_4
Xfanout595 _21720_/D vssd1 vssd1 vccd1 vccd1 _21412_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__21400__B1 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ _12921_/A _12921_/B _12921_/C vssd1 vssd1 vccd1 vccd1 _12924_/B sky130_fd_sc_hd__nand3_4
XANTENNA__17063__D _17086_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18737__A _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11165__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15640_ _15640_/A _15803_/B _15641_/B vssd1 vssd1 vccd1 vccd1 _15764_/A sky130_fd_sc_hd__or3b_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17641__A _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ _12853_/A _12853_/B vssd1 vssd1 vccd1 vccd1 _12966_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_38_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_96_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _11801_/A _11800_/Y _11776_/X _11777_/Y vssd1 vssd1 vccd1 vccd1 _11805_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_139_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15571_ _14508_/A _16084_/C _15954_/D _15838_/D vssd1 vssd1 vccd1 vccd1 _15575_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12783_ _12783_/A _12783_/B vssd1 vssd1 vccd1 vccd1 _12792_/A sky130_fd_sc_hd__nor2_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12785__A _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16257__A fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17310_ _17310_/A _17310_/B vssd1 vssd1 vccd1 vccd1 _17313_/A sky130_fd_sc_hd__xnor2_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19372__A2 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14522_ _14521_/B _14521_/C _14521_/A vssd1 vssd1 vccd1 vccd1 _14524_/B sky130_fd_sc_hd__a21o_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ _11734_/A _11734_/B _11734_/C vssd1 vssd1 vccd1 vccd1 _11736_/B sky130_fd_sc_hd__nand3_2
X_18290_ _18290_/A _18290_/B vssd1 vssd1 vccd1 vccd1 _18292_/B sky130_fd_sc_hd__xnor2_2
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17241_ _17240_/B _17240_/C _17240_/A vssd1 vssd1 vccd1 vccd1 _17243_/B sky130_fd_sc_hd__a21o_1
X_14453_ _14453_/A _14453_/B vssd1 vssd1 vccd1 vccd1 _14592_/A sky130_fd_sc_hd__or2_2
XANTENNA__19568__A _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11665_ _11665_/A vssd1 vssd1 vccd1 vccd1 _11666_/B sky130_fd_sc_hd__inv_2
XFILLER_0_138_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19124__A2 _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13404_ _14463_/D _13997_/C _13404_/C _13404_/D vssd1 vssd1 vccd1 vccd1 _13405_/B
+ sky130_fd_sc_hd__nand4_1
X_14384_ _14384_/A _15892_/B _14384_/C _14384_/D vssd1 vssd1 vccd1 vccd1 _14385_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_64_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17172_ _20770_/B _21331_/B vssd1 vssd1 vccd1 vccd1 _17172_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_36_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11596_ _12020_/A _12326_/D _12403_/A _12511_/A vssd1 vssd1 vccd1 vccd1 _11596_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_109_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16123_ _16123_/A vssd1 vssd1 vccd1 vccd1 _16123_/Y sky130_fd_sc_hd__inv_2
X_13335_ _13335_/A _13335_/B _13335_/C vssd1 vssd1 vccd1 vccd1 _13338_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_51_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14505__A _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16054_ _16054_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16055_/B sky130_fd_sc_hd__nand2_1
X_13266_ _13266_/A _13266_/B vssd1 vssd1 vccd1 vccd1 _13266_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11707__B1 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17238__D _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15005_ _15004_/B _15004_/C _15004_/A vssd1 vssd1 vccd1 vccd1 _15006_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_121_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12217_ _12217_/A _12217_/B _12217_/C vssd1 vssd1 vccd1 vccd1 _12217_/X sky130_fd_sc_hd__or3_1
XANTENNA__12670__D _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18635__A1 _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13197_ _13196_/A _13196_/B _13196_/C vssd1 vssd1 vccd1 vccd1 _13199_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_20_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19813_ _19813_/A _19813_/B vssd1 vssd1 vccd1 vccd1 _19814_/B sky130_fd_sc_hd__nor2_1
XANTENNA__17843__C1 _19030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ _12148_/A _12148_/B _12148_/C vssd1 vssd1 vccd1 vccd1 _12195_/A sky130_fd_sc_hd__nand3_1
XANTENNA__20242__A _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20734__A1_N _21261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15336__A _15336_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19744_ _19606_/A _19606_/C _19606_/B vssd1 vssd1 vccd1 vccd1 _19758_/A sky130_fd_sc_hd__a21bo_1
X_16956_ _16956_/A _16956_/B _16956_/C vssd1 vssd1 vccd1 vccd1 _16956_/Y sky130_fd_sc_hd__nand3_1
X_12079_ _12079_/A _12079_/B vssd1 vssd1 vccd1 vccd1 _12083_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__18399__B1 _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14672__A2 _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15907_ _15907_/A _15907_/B _15907_/C vssd1 vssd1 vccd1 vccd1 _15909_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_95_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19675_ _19673_/Y _19675_/B vssd1 vssd1 vccd1 vccd1 _19678_/A sky130_fd_sc_hd__nand2b_1
X_16887_ _16888_/B vssd1 vssd1 vccd1 vccd1 _16887_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_78_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18626_ _18626_/A _18626_/B vssd1 vssd1 vccd1 vccd1 _18628_/B sky130_fd_sc_hd__or2_1
XFILLER_0_56_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15838_ _15702_/D _15838_/B _16314_/D _15838_/D vssd1 vssd1 vccd1 vccd1 _15971_/A
+ sky130_fd_sc_hd__and4b_2
XANTENNA__17610__A2 _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18557_ _18429_/D _18430_/B _18555_/X _18709_/B vssd1 vssd1 vccd1 vccd1 _18559_/A
+ sky130_fd_sc_hd__a211o_1
X_15769_ _15769_/A _15769_/B vssd1 vssd1 vccd1 vccd1 _15772_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17508_ _17629_/A _17508_/B vssd1 vssd1 vccd1 vccd1 _17510_/B sky130_fd_sc_hd__and2_1
XFILLER_0_118_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18488_ _18489_/B _18489_/A vssd1 vssd1 vccd1 vccd1 _18632_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_145_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21170__A2 _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12845__D _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_14 _11335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17439_ _17439_/A _17439_/B vssd1 vssd1 vccd1 vccd1 _17441_/B sky130_fd_sc_hd__xnor2_2
XANTENNA_25 _11339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_36 _11430_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_47 hold247/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_58 hold270/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20450_ _20450_/A _20450_/B _20450_/C vssd1 vssd1 vccd1 vccd1 _20450_/X sky130_fd_sc_hd__or3_4
XANTENNA_69 hold268/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19109_ _19430_/A _19951_/B _19753_/B _19751_/C vssd1 vssd1 vccd1 vccd1 _19276_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_67_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20381_ _20381_/A _20381_/B vssd1 vssd1 vccd1 vccd1 _21146_/B sky130_fd_sc_hd__and2_1
XANTENNA__14415__A _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout117_A _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20136__B _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22051_ _22063_/CLK _22051_/D vssd1 vssd1 vccd1 vccd1 hold247/A sky130_fd_sc_hd__dfxtp_4
XFILLER_0_2_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17726__A _21795_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19644__C _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21002_ _20871_/X _20873_/X _21000_/Y _21001_/X vssd1 vssd1 vccd1 vccd1 _21005_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__16987__D _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout486_A _21747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15246__A _15246_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21904_ _21938_/CLK hold138/X vssd1 vssd1 vccd1 vccd1 hold137/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21835_ _21837_/CLK _21835_/D vssd1 vssd1 vccd1 vccd1 _21835_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12977__A2 _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21766_ _21767_/CLK _21766_/D vssd1 vssd1 vccd1 vccd1 _21766_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_77_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15412__C _15933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20717_ _20845_/D _21291_/B _20717_/C _20717_/D vssd1 vssd1 vccd1 vccd1 _20843_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_19_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21697_ _22080_/CLK _21697_/D vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13926__A1 _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11450_ _11123_/A t1y[0] t0x[0] _21724_/D vssd1 vssd1 vccd1 vccd1 _11450_/X sky130_fd_sc_hd__a22o_1
XANTENNA__13926__B2 _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20648_ hold276/X _20647_/X fanout2/X vssd1 vssd1 vccd1 vccd1 _21911_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11949__A _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ _11124_/A hold242/X fanout45/X hold199/X vssd1 vssd1 vccd1 vccd1 _11381_/X
+ sky130_fd_sc_hd__a22o_1
X_20579_ _20578_/B _20578_/C _20578_/A vssd1 vssd1 vccd1 vccd1 _20579_/X sky130_fd_sc_hd__o21a_1
X_13120_ _14936_/D _21776_/Q _13258_/D _14306_/A vssd1 vssd1 vccd1 vccd1 _13121_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12771__C _12771_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20046__B _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13051_ _13051_/A _13051_/B _13051_/C vssd1 vssd1 vccd1 vccd1 _13054_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_108_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17636__A _18010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16540__A _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14979__B _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ _12003_/A _12003_/B vssd1 vssd1 vccd1 vccd1 _12002_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_121_1240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21158__A _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14698__C _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16810_ _16810_/A _16810_/B _16810_/C vssd1 vssd1 vccd1 vccd1 _16823_/A sky130_fd_sc_hd__nand3_1
XANTENNA__14060__A _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17790_ _17790_/A _17790_/B vssd1 vssd1 vccd1 vccd1 _17799_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout370 _12402_/B vssd1 vssd1 vccd1 vccd1 _13573_/D sky130_fd_sc_hd__buf_4
Xfanout381 _21773_/Q vssd1 vssd1 vccd1 vccd1 _12858_/C sky130_fd_sc_hd__buf_4
Xfanout392 _15892_/B vssd1 vssd1 vccd1 vccd1 _14212_/B sky130_fd_sc_hd__clkbuf_8
X_16741_ _16741_/A _16741_/B _16741_/C vssd1 vssd1 vccd1 vccd1 _16754_/A sky130_fd_sc_hd__nand3_4
X_13953_ _13972_/B _13952_/B _13952_/C _13952_/D vssd1 vssd1 vccd1 vccd1 _13953_/X
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14995__A _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13862__B1 _14663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18467__A _19092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17053__B1 _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12904_ _12904_/A _12904_/B vssd1 vssd1 vccd1 vccd1 _12924_/A sky130_fd_sc_hd__xnor2_2
X_19460_ _19460_/A _19460_/B vssd1 vssd1 vccd1 vccd1 _19461_/B sky130_fd_sc_hd__xor2_2
X_16672_ _16672_/A _16672_/B _16672_/C vssd1 vssd1 vccd1 vccd1 _16676_/A sky130_fd_sc_hd__nand3_4
X_13884_ _13884_/A _13884_/B _13884_/C vssd1 vssd1 vccd1 vccd1 _13884_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_9_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18411_ _18411_/A _18411_/B vssd1 vssd1 vccd1 vccd1 _18414_/C sky130_fd_sc_hd__xnor2_1
X_15623_ _15753_/B _15621_/X _15483_/Y _15486_/Y vssd1 vssd1 vccd1 vccd1 _15624_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_97_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19391_ _19692_/A _20148_/C _19392_/C _19543_/A vssd1 vssd1 vccd1 vccd1 _19393_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ _12721_/A _12834_/A _12731_/B _12969_/A _12834_/Y vssd1 vssd1 vccd1 vccd1
+ _12837_/C sky130_fd_sc_hd__o32ai_4
XFILLER_0_154_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13404__A _14463_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18342_ _18343_/A _18343_/B vssd1 vssd1 vccd1 vccd1 _18478_/B sky130_fd_sc_hd__and2_1
XFILLER_0_69_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15554_ _15554_/A _15669_/B vssd1 vssd1 vccd1 vccd1 _15556_/B sky130_fd_sc_hd__or2_1
XFILLER_0_115_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16159__A2 _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ _12766_/A _12766_/B _12766_/C vssd1 vssd1 vccd1 vccd1 _12766_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_130_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10979__A1 _10978_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18553__B1 _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14505_ _16203_/D _15695_/A _14817_/C _14817_/D vssd1 vssd1 vccd1 vccd1 _14508_/D
+ sky130_fd_sc_hd__nand4_1
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18273_ _18273_/A _18273_/B vssd1 vssd1 vccd1 vccd1 _18275_/B sky130_fd_sc_hd__xnor2_1
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11717_ _11718_/A _11718_/B vssd1 vssd1 vccd1 vccd1 _12336_/B sky130_fd_sc_hd__nand2_1
X_15485_ _15315_/A _15315_/B _15313_/Y vssd1 vssd1 vccd1 vccd1 _15487_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_2_3__f_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12697_ _12716_/B _12697_/B _12697_/C _12697_/D vssd1 vssd1 vccd1 vccd1 _12697_/Y
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17224_ _17433_/A _17417_/A _19951_/A _17324_/D vssd1 vssd1 vccd1 vccd1 _17224_/X
+ sky130_fd_sc_hd__and4_1
X_14436_ _14273_/A _14273_/C _14270_/Y vssd1 vssd1 vccd1 vccd1 _14438_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_86_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11648_ _11648_/A _11648_/B vssd1 vssd1 vccd1 vccd1 _11649_/B sky130_fd_sc_hd__nor2_1
XANTENNA__21340__B _21340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15976__D _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11859__A _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17155_ _17120_/X _17136_/Y _17154_/X _17118_/Y _17110_/X vssd1 vssd1 vccd1 vccd1
+ _17159_/B sky130_fd_sc_hd__a2111o_1
XANTENNA__18856__A1 _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14367_ _14367_/A _16286_/A _14367_/C _14513_/A vssd1 vssd1 vccd1 vccd1 _14513_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_3_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18856__B2 _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11579_ _11579_/A _11579_/B vssd1 vssd1 vccd1 vccd1 _11585_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_13_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16106_ _16196_/B _21784_/Q _16104_/Y _16212_/A vssd1 vssd1 vccd1 vccd1 _16108_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16867__B1 _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13318_ _13318_/A _13318_/B vssd1 vssd1 vccd1 vccd1 _13338_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_52_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14298_ _12291_/B _14296_/Y _14297_/X vssd1 vssd1 vccd1 vccd1 _14298_/X sky130_fd_sc_hd__a21o_1
X_17086_ _17146_/A _17146_/B _17086_/C _17123_/C vssd1 vssd1 vccd1 vccd1 _17089_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_12_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16037_ _16036_/A _15906_/B _15907_/A vssd1 vssd1 vccd1 vccd1 _16038_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_122_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13249_ _13249_/A _13249_/B vssd1 vssd1 vccd1 vccd1 _13252_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_58_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20415__A1 _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20415__B2 _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17988_ _17989_/A _17989_/B vssd1 vssd1 vccd1 vccd1 _17988_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_74_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19727_ _19847_/A _19592_/X _19847_/B _19844_/C vssd1 vssd1 vccd1 vccd1 _19740_/A
+ sky130_fd_sc_hd__o211ai_1
X_16939_ _16989_/C _17146_/C vssd1 vssd1 vccd1 vccd1 _16984_/A sky130_fd_sc_hd__nand2_1
XANTENNA__20179__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19658_ _19658_/A _19658_/B vssd1 vssd1 vccd1 vccd1 _19659_/B sky130_fd_sc_hd__and2_1
XFILLER_0_95_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18609_ _18608_/B _18608_/C _18608_/A vssd1 vssd1 vccd1 vccd1 _18609_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_149_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19589_ _19439_/A _20247_/C _19723_/B _19723_/C vssd1 vssd1 vccd1 vccd1 _19589_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11533__S _11545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21620_ _21906_/CLK _21620_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[83] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_47_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21143__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18544__B1 _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11092__A0 _11048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21551_ mstream_o[14] hold8/X _21562_/S vssd1 vssd1 vccd1 vccd1 _22078_/D sky130_fd_sc_hd__mux2_1
XANTENNA__11631__A2 _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout234_A _17924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20502_ _20499_/Y _20500_/X _20355_/C _20355_/Y vssd1 vssd1 vccd1 vccd1 _20502_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20792__D _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21482_ hold161/X sstream_i[59] _21507_/S vssd1 vssd1 vccd1 vccd1 _22009_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_15_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16570__A2 _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20433_ _20558_/A _21283_/A _21171_/A _20433_/D vssd1 vssd1 vccd1 vccd1 _20558_/B
+ sky130_fd_sc_hd__and4b_1
XANTENNA_fanout401_A _21769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11395__A1 _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20364_ _20185_/A _20185_/B _20183_/Y vssd1 vssd1 vccd1 vccd1 _20366_/B sky130_fd_sc_hd__o21ai_1
X_22103_ _22105_/CLK _22103_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[39] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20295_ _20295_/A _20449_/A _20295_/C vssd1 vssd1 vccd1 vccd1 _20449_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_105_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12344__B1 _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22034_ _22038_/CLK _22034_/D vssd1 vssd1 vccd1 vccd1 hold235/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17606__D _18894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14636__A2 _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19390__B _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12647__A1 _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10950_ _10950_/A _10950_/B vssd1 vssd1 vccd1 vccd1 _10950_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_98_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16519__B _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10881_ _10885_/B _10881_/B vssd1 vssd1 vccd1 vccd1 _10881_/X sky130_fd_sc_hd__and2_2
XFILLER_0_151_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11443__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12620_ _12619_/A _13269_/C _12991_/D _13556_/A vssd1 vssd1 vccd1 vccd1 _12620_/Y
+ sky130_fd_sc_hd__a22oi_1
X_21818_ _21821_/CLK _21818_/D vssd1 vssd1 vccd1 vccd1 _21818_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_109_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11083__A0 _10959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18734__B _19053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ _13157_/A _13017_/A _12897_/C _12897_/D vssd1 vssd1 vccd1 vccd1 _12551_/X
+ sky130_fd_sc_hd__and4_1
X_21749_ _22038_/CLK _21749_/D vssd1 vssd1 vccd1 vccd1 _21749_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_108_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11502_ _11502_/A1 t2x[17] v1z[17] fanout20/X _11501_/X vssd1 vssd1 vccd1 vccd1 _11502_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15270_ _15270_/A _15270_/B vssd1 vssd1 vccd1 vccd1 _15286_/A sky130_fd_sc_hd__xor2_2
X_12482_ _12379_/B _12379_/Y _12479_/Y _12480_/X vssd1 vssd1 vccd1 vccd1 _12484_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14221_ _14062_/A _14062_/B _14062_/C vssd1 vssd1 vccd1 vccd1 _14222_/C sky130_fd_sc_hd__a21bo_1
X_11433_ hold272/A fanout28/X _11432_/X vssd1 vssd1 vccd1 vccd1 _11433_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11679__A _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18172__D _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14055__A _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11386__A1 _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14152_ _14031_/A _14030_/B _14028_/X vssd1 vssd1 vccd1 vccd1 _14162_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_151_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11364_ hold192/X fanout29/X _11363_/X vssd1 vssd1 vccd1 vccd1 _11364_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16313__A2 _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14324__A1 _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13103_ _13243_/A _13103_/B vssd1 vssd1 vccd1 vccd1 _13104_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_0_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14083_ _14713_/A _14557_/D _15234_/C _14572_/A vssd1 vssd1 vccd1 vccd1 _14083_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14324__B2 _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18960_ _18960_/A _18960_/B vssd1 vssd1 vccd1 vccd1 _18969_/A sky130_fd_sc_hd__xor2_2
X_11295_ fanout58/X v0z[17] fanout18/X _11294_/X vssd1 vssd1 vccd1 vccd1 _11295_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14875__A2 _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ _13173_/C _15076_/A _15076_/B _13034_/D vssd1 vssd1 vccd1 vccd1 _13169_/A
+ sky130_fd_sc_hd__nand4_2
X_17911_ _17910_/B _17910_/C _17910_/A vssd1 vssd1 vccd1 vccd1 _17912_/B sky130_fd_sc_hd__a21o_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19263__A1 _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18891_ _19051_/A _19382_/B _19051_/C _20317_/D vssd1 vssd1 vccd1 vccd1 _18894_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11689__A2 _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12886__B2 _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17842_ _17825_/A _17825_/B _17823_/X vssd1 vssd1 vccd1 vccd1 _17966_/A sky130_fd_sc_hd__a21bo_2
XFILLER_0_100_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14088__B1 hold319/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18909__B _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13118__B _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17773_ _17891_/B _17772_/C _17772_/A vssd1 vssd1 vccd1 vccd1 _17773_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12638__A1 _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14985_ _14984_/B _14984_/C _14984_/A vssd1 vssd1 vccd1 vccd1 _14985_/X sky130_fd_sc_hd__a21o_1
XANTENNA__20520__A _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12638__B2 _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19512_ _19512_/A _19512_/B _19512_/C vssd1 vssd1 vccd1 vccd1 _19514_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_89_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16724_ _17141_/A _17146_/B _17526_/B _17223_/A vssd1 vssd1 vccd1 vccd1 _16727_/A
+ sky130_fd_sc_hd__nand4_1
X_13936_ _13936_/A _13936_/B _13936_/C vssd1 vssd1 vccd1 vccd1 _13939_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_156_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11310__A1 _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19443_ _19440_/X _19441_/Y _19291_/A _19291_/B vssd1 vssd1 vccd1 vccd1 _19444_/B
+ sky130_fd_sc_hd__a211oi_1
X_16655_ _16633_/X _16635_/Y _16653_/A _16653_/Y vssd1 vssd1 vccd1 vccd1 _16657_/D
+ sky130_fd_sc_hd__o211a_1
X_13867_ _13867_/A _16273_/A _13867_/C _13867_/D vssd1 vssd1 vccd1 vccd1 _13867_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11861__A2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13236__A2_N _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15606_ _15605_/B _15605_/C _15605_/A vssd1 vssd1 vccd1 vccd1 _15606_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11580__C _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19374_ _21278_/A _19373_/X _19372_/X vssd1 vssd1 vccd1 vccd1 _19376_/A sky130_fd_sc_hd__a21bo_1
X_12818_ _12818_/A _12818_/B _12818_/C vssd1 vssd1 vccd1 vccd1 _12947_/B sky130_fd_sc_hd__or3_1
X_16586_ _16586_/A _16586_/B vssd1 vssd1 vccd1 vccd1 _16599_/A sky130_fd_sc_hd__nand2_2
X_13798_ _13795_/X _13796_/Y _13643_/C _13642_/Y vssd1 vssd1 vccd1 vccd1 _13800_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_85_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11074__A0 _10892_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18325_ _18326_/A _18326_/B vssd1 vssd1 vccd1 vccd1 _18325_/X sky130_fd_sc_hd__and2_1
XFILLER_0_45_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15537_ _15663_/A vssd1 vssd1 vccd1 vccd1 _15539_/D sky130_fd_sc_hd__inv_2
XFILLER_0_127_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ _12837_/A _12747_/X _12630_/B _12631_/Y vssd1 vssd1 vccd1 vccd1 _12808_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12973__A _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16445__A _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18256_ _19185_/D _19008_/D _19199_/C _19199_/D vssd1 vssd1 vccd1 vccd1 _18402_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_71_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15468_ _15465_/X _15466_/Y _15327_/Y _15332_/A vssd1 vssd1 vccd1 vccd1 _15469_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_115_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17207_ _17520_/A _17520_/B _17417_/C _17417_/D vssd1 vssd1 vccd1 vccd1 _17207_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_5_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11589__A _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14419_ _14419_/A _14419_/B vssd1 vssd1 vccd1 vccd1 _14422_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_114_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18468__A1_N _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15760__B1 _10950_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18187_ _18787_/B _18773_/B _19546_/D _18787_/A vssd1 vssd1 vccd1 vccd1 _18187_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_53_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15399_ _15399_/A _15541_/B vssd1 vssd1 vccd1 vccd1 _15402_/A sky130_fd_sc_hd__or2_1
XANTENNA__11377__A1 _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17138_ _17133_/A _17132_/C _17132_/B vssd1 vssd1 vccd1 vccd1 _17138_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_40_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16304__A2 _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17501__A1 _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17069_ _17069_/A _17069_/B vssd1 vssd1 vccd1 vccd1 _17071_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_988 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20080_ _19796_/A _19941_/A _19943_/B vssd1 vssd1 vccd1 vccd1 _20080_/X sky130_fd_sc_hd__a21o_1
XANTENNA__15508__B _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20939__A2 _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11755__C _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17280__A3 _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout184_A _17666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15524__A _16036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17032__A1_N _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20982_ _20983_/A _20983_/B vssd1 vssd1 vccd1 vccd1 _20984_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11301__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout351_A hold241/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13044__A _14712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21261__A _21261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18554__B _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21603_ _21888_/CLK _21603_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[66] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_36_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout616_A _21717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21534_ hold268/X sstream_i[111] _21536_/S vssd1 vssd1 vccd1 vccd1 _22061_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17740__A1 _18010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17740__B2 _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19666__A _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21465_ hold210/X sstream_i[42] _21494_/S vssd1 vssd1 vccd1 vccd1 _21992_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_105_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11368__A1 _17086_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14306__C _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20416_ _20416_/A _20416_/B _20924_/A _21305_/A vssd1 vssd1 vccd1 vccd1 _20552_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21396_ _21720_/D _21396_/B vssd1 vssd1 vccd1 vccd1 _21396_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_114_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16802__B _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12107__B _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20347_ _20344_/X _20345_/Y _20199_/Y _20201_/X vssd1 vssd1 vccd1 vccd1 _20348_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_105_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout97_A _21843_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11080_ _10941_/X hold7/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21675_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_41_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20278_ _20279_/A _20279_/B vssd1 vssd1 vccd1 vccd1 _20486_/B sky130_fd_sc_hd__or2_1
XANTENNA__13864__D _14663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22017_ _22020_/CLK _22017_/D vssd1 vssd1 vccd1 vccd1 hold192/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11540__A1 _11089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14770_ _14936_/D _15698_/B vssd1 vssd1 vccd1 vccd1 _14771_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13293__A1 _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11982_ _11982_/A _11982_/B vssd1 vssd1 vccd1 vccd1 _12286_/A sky130_fd_sc_hd__and2_1
XANTENNA__13293__B2 _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13721_ _13875_/B _14516_/A _14365_/C _13877_/A vssd1 vssd1 vccd1 vccd1 _13724_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15153__B _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10933_ _10926_/A _10926_/B _10931_/Y _10923_/B vssd1 vssd1 vccd1 vccd1 _10934_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16440_ hold232/X _16439_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _21885_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13045__A1 _14712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10864_ _10864_/A _10873_/A vssd1 vssd1 vccd1 vccd1 _10864_/Y sky130_fd_sc_hd__nand2_1
X_13652_ _13652_/A _13652_/B _13652_/C _13652_/D vssd1 vssd1 vccd1 vccd1 _13652_/Y
+ sky130_fd_sc_hd__nor4_4
XANTENNA__16886__A1_N _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13045__B2 _14712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11056__A0 _11055_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18464__B _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19183__A1_N _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21171__A _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12603_ hold74/X _12602_/X fanout3/X vssd1 vssd1 vccd1 vccd1 hold75/A sky130_fd_sc_hd__mux2_1
XFILLER_0_52_1171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16371_ _16371_/A _21755_/Q vssd1 vssd1 vccd1 vccd1 _16372_/B sky130_fd_sc_hd__nand2_1
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13583_ _13450_/X _13453_/Y _13581_/Y _13582_/X vssd1 vssd1 vccd1 vccd1 _13583_/X
+ sky130_fd_sc_hd__a211o_2
X_10795_ _20838_/B vssd1 vssd1 vccd1 vccd1 _21199_/B sky130_fd_sc_hd__inv_2
XFILLER_0_26_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19279__C _19751_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18110_ _19008_/D _21791_/Q _19199_/C _19199_/D vssd1 vssd1 vccd1 vccd1 _18253_/A
+ sky130_fd_sc_hd__and4_1
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15322_ _15322_/A _15450_/B vssd1 vssd1 vccd1 vccd1 _15324_/B sky130_fd_sc_hd__or2_1
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19090_ _19090_/A _19090_/B vssd1 vssd1 vccd1 vccd1 _19099_/A sky130_fd_sc_hd__xnor2_1
X_12534_ _12877_/A _12642_/A _13155_/C _13155_/D vssd1 vssd1 vccd1 vccd1 _12534_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18041_ _18164_/A _18040_/C _18040_/A vssd1 vssd1 vccd1 vccd1 _18042_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_151_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15253_ _15253_/A _15253_/B vssd1 vssd1 vccd1 vccd1 _15290_/A sky130_fd_sc_hd__and2_1
XFILLER_0_81_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12465_ _12465_/A _12465_/B _12465_/C vssd1 vssd1 vccd1 vccd1 _12468_/A sky130_fd_sc_hd__nand3_2
XANTENNA__11359__A1 _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14204_ _14203_/B _14203_/C _14203_/A vssd1 vssd1 vccd1 vccd1 _14204_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11416_ _11415_/X _17670_/B _11446_/S vssd1 vssd1 vccd1 vccd1 _21810_/D sky130_fd_sc_hd__mux2_1
X_15184_ _15331_/B _15182_/Y _14956_/X _14958_/Y vssd1 vssd1 vccd1 vccd1 _15185_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12396_ _13525_/A _13258_/C _13258_/D _12312_/A vssd1 vssd1 vccd1 vccd1 _12399_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14135_ _14321_/A _14135_/B vssd1 vssd1 vccd1 vccd1 _14136_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11347_ _21407_/S v0z[30] fanout20/X _11346_/X vssd1 vssd1 vccd1 vccd1 _11347_/X
+ sky130_fd_sc_hd__a31o_2
XANTENNA__17096__A _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19992_ _21291_/A _20416_/B _21296_/A _20416_/A vssd1 vssd1 vccd1 vccd1 _19995_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14066_ _14066_/A _14209_/A _14066_/C vssd1 vssd1 vccd1 vccd1 _14209_/B sky130_fd_sc_hd__nand3_1
XANTENNA__12859__A1 _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11278_ _11493_/A1 t1x[13] v2z[13] _11501_/B2 _11277_/X vssd1 vssd1 vccd1 vccd1 _11278_/X
+ sky130_fd_sc_hd__a221o_2
X_18943_ _19084_/B _18942_/C _18942_/A vssd1 vssd1 vccd1 vccd1 _18944_/C sky130_fd_sc_hd__a21o_1
XANTENNA__12859__B2 _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11348__S _11348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13017_ _13017_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _13020_/A sky130_fd_sc_hd__and2_1
X_18874_ _18874_/A _18874_/B _19028_/B vssd1 vssd1 vccd1 vccd1 _18876_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_20_1126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11531__A1 _11089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17825_ _17825_/A _17825_/B vssd1 vssd1 vccd1 vccd1 _17828_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__21346__A _21349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17543__B _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
X_17756_ _17664_/A _17663_/B _17661_/X vssd1 vssd1 vccd1 vccd1 _17772_/A sky130_fd_sc_hd__a21o_1
X_14968_ _14968_/A _14968_/B vssd1 vssd1 vccd1 vccd1 _14970_/B sky130_fd_sc_hd__xnor2_1
X_16707_ _16705_/A _16705_/Y _16706_/Y _16675_/X vssd1 vssd1 vccd1 vccd1 _16712_/B
+ sky130_fd_sc_hd__a211o_2
X_13919_ _13919_/A _13919_/B vssd1 vssd1 vccd1 vccd1 _13939_/A sky130_fd_sc_hd__xor2_1
XANTENNA__11295__B1 _11294_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17687_ _17683_/X _17685_/Y _17570_/B _17570_/Y vssd1 vssd1 vccd1 vccd1 _17689_/D
+ sky130_fd_sc_hd__o211a_1
X_14899_ _14900_/B _14900_/A vssd1 vssd1 vccd1 vccd1 _14899_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_76_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19426_ _19426_/A _19426_/B vssd1 vssd1 vccd1 vccd1 _19453_/A sky130_fd_sc_hd__and2_2
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16638_ _17146_/A _18166_/A _17434_/B _17146_/B vssd1 vssd1 vccd1 vccd1 _16639_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19357_ _19356_/B _19356_/C _19356_/A vssd1 vssd1 vccd1 vccd1 _19358_/C sky130_fd_sc_hd__a21o_1
X_16569_ _17621_/C _17300_/C _17520_/D _17504_/C vssd1 vssd1 vccd1 vccd1 _16569_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_31_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16175__A _16284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11598__A1 _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18308_ _18305_/Y _18306_/X _18183_/B _18183_/Y vssd1 vssd1 vccd1 vccd1 _18308_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11598__B2 _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16606__C _17557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19288_ _19439_/A _20242_/D vssd1 vssd1 vccd1 vccd1 _19289_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14536__A1 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13311__B _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18239_ _18389_/A _18239_/B vssd1 vssd1 vccd1 vccd1 _18241_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_5_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20128__C _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21250_ _11550_/A _21248_/Y _21249_/X vssd1 vssd1 vccd1 vccd1 _21250_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_41_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18278__A2 _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20201_ _20202_/A _20202_/B vssd1 vssd1 vccd1 vccd1 _20201_/X sky130_fd_sc_hd__and2_1
XANTENNA__20085__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21181_ _21182_/A _21182_/B vssd1 vssd1 vccd1 vccd1 _21181_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_13_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20132_ _20416_/B _20273_/A _20270_/C _20416_/A vssd1 vssd1 vccd1 vccd1 _20136_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout399_A _21770_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20063_ _19837_/A _19838_/X _20216_/A _20062_/X vssd1 vssd1 vccd1 vccd1 _20216_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11522__A1 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17789__A1 _17670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21256__A _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout566_A _12403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16461__A1 _16743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_307 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_318 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_329 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20965_ _21293_/A _21286_/B _21296_/B _21199_/A vssd1 vssd1 vccd1 vccd1 _20969_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20896_ _20896_/A _20896_/B vssd1 vssd1 vccd1 vccd1 _20898_/B sky130_fd_sc_hd__or2_1
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12786__B1 _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19702__A2 _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout12_A _11446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21517_ hold237/X sstream_i[94] _21528_/S vssd1 vssd1 vccd1 vccd1 _22044_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_145_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_clk_i _21806_/CLK vssd1 vssd1 vccd1 vccd1 _21809_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16813__A _16813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12250_ _12245_/X _12248_/X _12217_/X _12244_/Y vssd1 vssd1 vccd1 vccd1 _12250_/X
+ sky130_fd_sc_hd__o211a_1
X_21448_ hold293/X sstream_i[25] _21489_/S vssd1 vssd1 vccd1 vccd1 _21975_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_82_1131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11210__A0 _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11201_ _14077_/B _11200_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21750_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_31_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21273__A1 _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21273__B2 _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12181_ _12268_/A _12246_/C vssd1 vssd1 vccd1 vccd1 _12183_/B sky130_fd_sc_hd__and2_1
X_21379_ _14449_/B _19322_/Y _21420_/S vssd1 vssd1 vccd1 vccd1 _21379_/X sky130_fd_sc_hd__mux2_1
XANTENNA__13875__C _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_1186 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17554__A1_N _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11132_ _12269_/C _11131_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21727_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13594__D _14212_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11168__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20989__B _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15940_ _15940_/A _15940_/B _15940_/C vssd1 vssd1 vccd1 vccd1 _15941_/C sky130_fd_sc_hd__nand3_1
X_11063_ _11063_/A _11063_/B vssd1 vssd1 vccd1 vccd1 _11063_/X sky130_fd_sc_hd__xor2_4
XANTENNA__11513__A1 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15871_ _15952_/B _15868_/Y _15687_/B _15689_/B vssd1 vssd1 vccd1 vccd1 _15871_/X
+ sky130_fd_sc_hd__a211o_1
X_17610_ _19337_/D _20797_/A _21258_/A _18851_/C vssd1 vssd1 vccd1 vccd1 _17611_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11692__A _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14822_ _14818_/X _14820_/Y _14662_/X _14665_/X vssd1 vssd1 vccd1 vccd1 _14823_/B
+ sky130_fd_sc_hd__a211o_1
X_18590_ _18590_/A _18590_/B vssd1 vssd1 vccd1 vccd1 _18592_/B sky130_fd_sc_hd__xnor2_1
XTAP_3830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21328__A2 _11553_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17541_ _17446_/A _17445_/B _17445_/A vssd1 vssd1 vccd1 vccd1 _17548_/A sky130_fd_sc_hd__o21ba_1
XTAP_3863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14753_ _14754_/A _14754_/B vssd1 vssd1 vccd1 vccd1 _14753_/Y sky130_fd_sc_hd__nor2_1
XTAP_3874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11965_ _11872_/Y _11873_/X _11899_/B _11892_/D vssd1 vssd1 vccd1 vccd1 _11965_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XFILLER_0_58_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11842__D _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12300__B _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16204__B2 _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13704_ _13858_/B _13858_/C _13402_/D _14936_/D vssd1 vssd1 vccd1 vccd1 _13707_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10916_ _10916_/A _10924_/A vssd1 vssd1 vccd1 vccd1 _10919_/A sky130_fd_sc_hd__or2_2
X_17472_ _17360_/C _17362_/A _17470_/X _17471_/X vssd1 vssd1 vccd1 vccd1 _17474_/A
+ sky130_fd_sc_hd__o211a_1
X_14684_ _14684_/A _14809_/A _14684_/C vssd1 vssd1 vccd1 vccd1 _14809_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_6_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11896_ _11830_/Y _11893_/X _11892_/X _11872_/Y vssd1 vssd1 vccd1 vccd1 _11901_/B
+ sky130_fd_sc_hd__a211o_1
X_19211_ _19037_/X _19211_/B vssd1 vssd1 vccd1 vccd1 _19213_/B sky130_fd_sc_hd__and2b_1
X_16423_ _16423_/A _16423_/B vssd1 vssd1 vccd1 vccd1 _16433_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13635_ _13635_/A _13635_/B _13635_/C vssd1 vssd1 vccd1 vccd1 _13638_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_132_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10847_ hold315/A hold122/A vssd1 vssd1 vccd1 vccd1 _11063_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_132_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14508__A _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19142_ _19139_/Y _19140_/X _18979_/B _18979_/Y vssd1 vssd1 vccd1 vccd1 _19143_/C
+ sky130_fd_sc_hd__a211o_1
X_16354_ _16354_/A _16354_/B vssd1 vssd1 vccd1 vccd1 _16356_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13566_ _13567_/A _13567_/B vssd1 vssd1 vccd1 vccd1 _13690_/B sky130_fd_sc_hd__or2_1
XFILLER_0_87_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15305_ _15305_/A _15305_/B vssd1 vssd1 vccd1 vccd1 _15307_/B sky130_fd_sc_hd__or2_1
X_19073_ _19073_/A _19073_/B _19073_/C vssd1 vssd1 vccd1 vccd1 _19076_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12517_ _12517_/A _12517_/B vssd1 vssd1 vccd1 vccd1 _12519_/B sky130_fd_sc_hd__xor2_2
X_16285_ _16286_/A _16286_/B _16286_/C _16286_/D vssd1 vssd1 vccd1 vccd1 _16287_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15715__B1 _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13497_ _13496_/A _13496_/B _13496_/C _13496_/D vssd1 vssd1 vccd1 vccd1 _13497_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_48_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17180__A2 _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18024_ _17883_/B _17884_/Y _18107_/A _18023_/X vssd1 vssd1 vccd1 vccd1 _18107_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_35_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15236_ _15233_/Y _15377_/A _15375_/A _15368_/D vssd1 vssd1 vccd1 vccd1 _15377_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_140_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12448_ _12449_/A _12449_/B vssd1 vssd1 vccd1 vccd1 _12544_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_124_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11201__A0 _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13741__A2 _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15167_ _15167_/A _15167_/B vssd1 vssd1 vccd1 vccd1 _15185_/A sky130_fd_sc_hd__xnor2_1
X_12379_ _12379_/A _12379_/B _12379_/C vssd1 vssd1 vccd1 vccd1 _12379_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_1_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14118_ _14117_/B _14117_/C _14117_/A vssd1 vssd1 vccd1 vccd1 _14118_/Y sky130_fd_sc_hd__o21ai_1
X_15098_ _15375_/A _15098_/B _15098_/C _15238_/A vssd1 vssd1 vccd1 vccd1 _15238_/B
+ sky130_fd_sc_hd__nand4_4
XANTENNA__19753__B _19753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19975_ _19871_/X _19874_/X _19973_/X _20110_/B vssd1 vssd1 vccd1 vccd1 _20098_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_120_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11078__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14049_ _13884_/B _13884_/Y _14132_/A _14048_/Y vssd1 vssd1 vccd1 vccd1 _14132_/B
+ sky130_fd_sc_hd__a211oi_2
X_18926_ _18793_/A _18792_/B _18790_/X vssd1 vssd1 vccd1 vccd1 _18942_/A sky130_fd_sc_hd__a21o_1
XANTENNA__20775__B1 _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18857_ _19008_/D _18857_/B _19181_/B _19185_/B vssd1 vssd1 vccd1 vccd1 _18859_/D
+ sky130_fd_sc_hd__and4_1
XFILLER_0_119_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20411__C _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17808_ _17804_/X _17806_/Y _17684_/B _17684_/Y vssd1 vssd1 vccd1 vccd1 _17810_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18788_ _18789_/A _18789_/B _18789_/C _18947_/A vssd1 vssd1 vccd1 vccd1 _18790_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11268__A0 _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12848__D _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17739_ _18010_/A _17874_/A _17739_/C _17739_/D vssd1 vssd1 vccd1 vccd1 _17870_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20750_ _20750_/A vssd1 vssd1 vccd1 vccd1 _20750_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_148_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17720__C _19051_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19409_ _20101_/A _20101_/B _19906_/C vssd1 vssd1 vccd1 vccd1 _19409_/X sky130_fd_sc_hd__and3_1
XANTENNA__15521__B _15521_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20681_ _20681_/A _20681_/B vssd1 vssd1 vccd1 vccd1 _20683_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_58_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout147_A _19092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11440__A0 _11439_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1096 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout314_A _21792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21302_ _21146_/X _21183_/B _20788_/A _21034_/B vssd1 vssd1 vccd1 vccd1 _21303_/B
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17448__B _17557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21233_ _21234_/A _21234_/B vssd1 vssd1 vccd1 vccd1 _21255_/A sky130_fd_sc_hd__nand2b_1
Xhold220 hold220/A vssd1 vssd1 vccd1 vccd1 hold220/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold231 hold231/A vssd1 vssd1 vccd1 vccd1 hold231/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 hold314/A vssd1 vssd1 vccd1 vccd1 hold242/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 hold253/A vssd1 vssd1 vccd1 vccd1 hold253/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold264 hold264/A vssd1 vssd1 vccd1 vccd1 hold264/X sky130_fd_sc_hd__dlygate4sd3_1
X_21164_ _21164_/A vssd1 vssd1 vccd1 vccd1 _21178_/A sky130_fd_sc_hd__inv_2
Xhold275 hold275/A vssd1 vssd1 vccd1 vccd1 hold275/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 hold286/A vssd1 vssd1 vccd1 vccd1 hold286/X sky130_fd_sc_hd__buf_4
Xhold297 hold297/A vssd1 vssd1 vccd1 vccd1 hold297/X sky130_fd_sc_hd__dlygate4sd3_1
X_20115_ _20116_/A _20116_/B vssd1 vssd1 vccd1 vccd1 _20115_/X sky130_fd_sc_hd__and2_1
X_21095_ _21095_/A _21095_/B vssd1 vssd1 vccd1 vccd1 _21116_/A sky130_fd_sc_hd__xor2_2
XANTENNA__12299__A2 _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18279__B _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20046_ _20845_/D _20721_/D _20733_/C _20606_/D vssd1 vssd1 vccd1 vccd1 _20188_/A
+ sky130_fd_sc_hd__and4_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17183__B _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20230__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11259__B1 _11258_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_104 mstream_o[115] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18187__A1 _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_115 sstream_i[68] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_126 v0z[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18295__A _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21997_ _22021_/CLK _21997_/D vssd1 vssd1 vccd1 vccd1 hold153/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_137 v1z[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18187__B2 _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_148 v1z[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20975__D _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11750_ _11750_/A _11750_/B _11750_/C vssd1 vssd1 vccd1 vccd1 _11753_/B sky130_fd_sc_hd__nand3_4
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20948_ _20946_/X _20948_/B vssd1 vssd1 vccd1 vccd1 _20949_/B sky130_fd_sc_hd__and2b_1
XANTENNA_159 v2z[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16527__B _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11681_ _12109_/C _12750_/A _11680_/C _11705_/A vssd1 vssd1 vccd1 vccd1 _11682_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14328__A _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20879_ _20880_/B _20880_/C vssd1 vssd1 vccd1 vccd1 _20881_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_37_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13420_ _13417_/Y _13569_/A _13867_/A _13573_/D vssd1 vssd1 vccd1 vccd1 _13569_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_14_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19687__A1 fanout96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13589__D _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20991__C _20991_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11431__A0 _11430_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13351_ _13348_/X _13349_/Y _13209_/C _13208_/Y vssd1 vssd1 vccd1 vccd1 _13353_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14762__S fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12302_ _12302_/A _12402_/B _12302_/C _12302_/D vssd1 vssd1 vccd1 vccd1 _12305_/B
+ sky130_fd_sc_hd__and4_1
X_16070_ _16070_/A _16070_/B _16070_/C vssd1 vssd1 vccd1 vccd1 _16071_/A sky130_fd_sc_hd__and3_1
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13282_ _13166_/B _13168_/A _13280_/Y _13281_/X vssd1 vssd1 vccd1 vccd1 _13373_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15021_ _16196_/A _15791_/A _16196_/B _16371_/A vssd1 vssd1 vccd1 vccd1 _15024_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11687__A _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13723__A2 _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14920__A1 _12291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12233_ _12228_/A _12228_/B _12228_/C vssd1 vssd1 vccd1 vccd1 _12234_/C sky130_fd_sc_hd__a21oi_1
XANTENNA__19854__A _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18111__A1 _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18111__B2 _21791_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12164_ _12165_/A _12165_/B vssd1 vssd1 vccd1 vccd1 _12175_/A sky130_fd_sc_hd__nor2_1
XANTENNA__14998__A _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11115_ _10950_/Y hold28/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21709_/D sky130_fd_sc_hd__mux2_1
X_16972_ _16971_/B _16971_/C _16971_/A vssd1 vssd1 vccd1 vccd1 _16973_/C sky130_fd_sc_hd__a21bo_1
X_12095_ _12094_/A _12512_/A _12214_/C _12094_/B vssd1 vssd1 vccd1 vccd1 _12096_/B
+ sky130_fd_sc_hd__a22o_1
X_19760_ _19758_/B _19758_/C _19758_/A vssd1 vssd1 vccd1 vccd1 _19760_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15923_ _15923_/A _15923_/B vssd1 vssd1 vccd1 vccd1 _15925_/B sky130_fd_sc_hd__xor2_1
X_18711_ _18873_/A _19493_/D _19199_/C _19199_/D vssd1 vssd1 vccd1 vccd1 _18713_/D
+ sky130_fd_sc_hd__nand4_1
X_11046_ _11045_/X hold72/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21653_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17093__B _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19691_ _21199_/A _19692_/B _20416_/A _19691_/D vssd1 vssd1 vccd1 vccd1 _19691_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__15228__A2 _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18642_ _18641_/B _18784_/B _18641_/A vssd1 vssd1 vccd1 vccd1 _18643_/B sky130_fd_sc_hd__a21o_1
X_15854_ _15972_/A _15978_/B _16084_/A _15854_/D vssd1 vssd1 vccd1 vccd1 _15972_/B
+ sky130_fd_sc_hd__and4b_1
XANTENNA__12311__A _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14805_ _14806_/A _14806_/B vssd1 vssd1 vccd1 vccd1 _14924_/A sky130_fd_sc_hd__and2b_1
X_18573_ _18572_/B _18572_/C _18572_/A vssd1 vssd1 vccd1 vccd1 _18573_/X sky130_fd_sc_hd__o21a_1
XTAP_3660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15785_ _15653_/C _16424_/A _15911_/C _16399_/A vssd1 vssd1 vccd1 vccd1 _15788_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12997_ _12997_/A _12997_/B _12997_/C vssd1 vssd1 vccd1 vccd1 _13000_/A sky130_fd_sc_hd__nand3_1
XTAP_3671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17524_ _17524_/A _17524_/B vssd1 vssd1 vccd1 vccd1 _17534_/A sky130_fd_sc_hd__and2_1
XFILLER_0_59_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14736_ _14576_/A _14576_/B _14574_/X vssd1 vssd1 vccd1 vccd1 _14738_/B sky130_fd_sc_hd__a21oi_4
XANTENNA__21343__B _21343_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ _11948_/A _11948_/B vssd1 vssd1 vccd1 vccd1 _11956_/A sky130_fd_sc_hd__nor2_1
XTAP_2970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16437__B _16437_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17455_ _17455_/A _17455_/B _17455_/C vssd1 vssd1 vccd1 vccd1 _17458_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_74_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14667_ _14504_/X _14507_/X _14664_/X _14666_/Y vssd1 vssd1 vccd1 vccd1 _14667_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11879_ _11879_/A _11948_/A vssd1 vssd1 vccd1 vccd1 _11881_/B sky130_fd_sc_hd__or2_1
XFILLER_0_131_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16406_ _16406_/A _16406_/B vssd1 vssd1 vccd1 vccd1 _16407_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_156_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13618_ _13618_/A _13618_/B vssd1 vssd1 vccd1 vccd1 _13638_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__20334__A1_N _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17386_ _17386_/A _17386_/B vssd1 vssd1 vccd1 vccd1 _17388_/A sky130_fd_sc_hd__nand2_1
X_14598_ _14599_/A _14599_/B vssd1 vssd1 vccd1 vccd1 _14608_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_43_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18652__B _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19125_ _21824_/Q _21171_/B vssd1 vssd1 vccd1 vccd1 _19126_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_70_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11422__A0 _11421_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16337_ _16337_/A _16337_/B _16337_/C vssd1 vssd1 vccd1 vccd1 _16337_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_15_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13549_ _13669_/B _13546_/X _13430_/X _13433_/Y vssd1 vssd1 vccd1 vccd1 _13549_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_82_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19056_ _19686_/B _19529_/B _19227_/C _19227_/D vssd1 vssd1 vccd1 vccd1 _19056_/X
+ sky130_fd_sc_hd__and4_1
X_16268_ _16377_/A _16268_/B vssd1 vssd1 vccd1 vccd1 _16269_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18007_ _18008_/A _18769_/B _17895_/X _17894_/X _18767_/B vssd1 vssd1 vccd1 vccd1
+ _18012_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_51_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15219_ _15218_/B _15361_/B _15218_/A vssd1 vssd1 vccd1 vccd1 _15220_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11597__A _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16199_ _16374_/A _16404_/B _16199_/C _16199_/D vssd1 vssd1 vccd1 vccd1 _16309_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_10_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19850__A1 _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_878 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19958_ _19958_/A _19958_/B _19958_/C vssd1 vssd1 vccd1 vccd1 _19961_/C sky130_fd_sc_hd__and3_1
XFILLER_0_77_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14701__A _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18909_ _19535_/A _19695_/A _20103_/A _19906_/A vssd1 vssd1 vccd1 vccd1 _19065_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__19602__A1 _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19889_ _20838_/B _21278_/A _20265_/D _20975_/D vssd1 vssd1 vccd1 vccd1 _19891_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11536__S _11545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17434__D _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21920_ _21923_/CLK _21920_/D vssd1 vssd1 vccd1 vccd1 hold193/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12221__A _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14978__A1 _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13036__B _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21851_ _21853_/CLK _21851_/D vssd1 vssd1 vccd1 vccd1 hold325/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__14978__B2 _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout264_A _19531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20802_ _20802_/A _20931_/B _20801_/X vssd1 vssd1 vccd1 vccd1 _20999_/A sky130_fd_sc_hd__or3b_2
XANTENNA__19905__A2 _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21782_ _21821_/CLK _21782_/D vssd1 vssd1 vccd1 vccd1 _21782_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17916__A1 _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12453__A2 _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17916__B2 _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20733_ _20863_/C _20991_/C _20733_/C _21305_/B vssd1 vssd1 vccd1 vccd1 _20857_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout431_A _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17392__A2 _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout529_A _21738_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20664_ _21034_/A _20664_/B vssd1 vssd1 vccd1 vccd1 _20665_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11413__A0 _11412_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20595_ _20465_/A _20600_/A _20464_/B _20461_/B _20461_/A vssd1 vssd1 vccd1 vccd1
+ _20597_/B sky130_fd_sc_hd__o32ai_4
XFILLER_0_144_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16363__A _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_1222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21216_ _21216_/A _21216_/B vssd1 vssd1 vccd1 vccd1 _21217_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20987__B1 _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21147_ _20788_/A _21034_/B _21146_/X vssd1 vssd1 vccd1 vccd1 _21183_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13469__A1 _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12830__S fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13469__B2 _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout530 _12877_/A vssd1 vssd1 vccd1 vccd1 _12443_/A sky130_fd_sc_hd__buf_4
Xfanout541 _13858_/A vssd1 vssd1 vccd1 vccd1 _12637_/A sky130_fd_sc_hd__buf_4
Xfanout552 _12530_/A vssd1 vssd1 vccd1 vccd1 _12619_/A sky130_fd_sc_hd__buf_4
XANTENNA__15426__B _15426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21078_ _21077_/A _21077_/B _21077_/C vssd1 vssd1 vccd1 vccd1 _21122_/B sky130_fd_sc_hd__a21oi_1
Xfanout563 _12403_/A vssd1 vssd1 vccd1 vccd1 _14463_/D sky130_fd_sc_hd__clkbuf_4
Xfanout574 _12268_/B vssd1 vssd1 vccd1 vccd1 _14133_/D sky130_fd_sc_hd__buf_4
XANTENNA__21400__A1 _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11446__S _11446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout585 _11447_/A1 vssd1 vssd1 vccd1 vccd1 _11124_/A sky130_fd_sc_hd__buf_4
Xfanout596 _21349_/A vssd1 vssd1 vccd1 vccd1 _21720_/D sky130_fd_sc_hd__buf_4
X_12920_ _12792_/A _12792_/C _12792_/B vssd1 vssd1 vccd1 vccd1 _12921_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__17604__B1 _18894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20029_ _20027_/X _20175_/B _19804_/D _19808_/B vssd1 vssd1 vccd1 vccd1 _20029_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_38_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11673__C _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_24_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21906_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18737__B _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12851_ _12851_/A _12851_/B vssd1 vssd1 vccd1 vccd1 _12853_/B sky130_fd_sc_hd__or2_1
XANTENNA__17641__B _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11802_ _11801_/A _11800_/Y _11776_/X _11777_/Y vssd1 vssd1 vccd1 vccd1 _11802_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15570_ _15567_/X _15568_/Y _15426_/B _15426_/Y vssd1 vssd1 vccd1 vccd1 _15612_/B
+ sky130_fd_sc_hd__a211oi_2
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ _13173_/C _12781_/D _12779_/Y _12780_/X vssd1 vssd1 vccd1 vccd1 _12783_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11247__A3 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12785__B _12785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14521_ _14521_/A _14521_/B _14521_/C vssd1 vssd1 vccd1 vccd1 _14524_/A sky130_fd_sc_hd__nand3_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11733_ _11732_/B _11732_/C _11732_/A vssd1 vssd1 vccd1 vccd1 _11734_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_96_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14058__A _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18580__A1 _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17240_ _17240_/A _17240_/B _17240_/C vssd1 vssd1 vccd1 vccd1 _17243_/A sky130_fd_sc_hd__nand3_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15394__A1 _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14452_ _14321_/A _14320_/Y _14319_/B vssd1 vssd1 vccd1 vccd1 _14596_/A sky130_fd_sc_hd__a21o_1
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11664_ _11664_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11665_/A sky130_fd_sc_hd__and2_1
XFILLER_0_3_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19568__B _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11404__A0 _11403_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13403_ _14463_/D hold241/A _13404_/C _13404_/D vssd1 vssd1 vccd1 vccd1 _13405_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17171_ _17171_/A _17171_/B vssd1 vssd1 vccd1 vccd1 _21331_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_64_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14383_ _14212_/B _14384_/C _14384_/D _14384_/A vssd1 vssd1 vccd1 vccd1 _14385_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16273__A _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11595_ _11595_/A _11595_/B vssd1 vssd1 vccd1 vccd1 _11602_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16122_ _15944_/Y _15948_/B _16120_/A _16121_/Y vssd1 vssd1 vccd1 vccd1 _16123_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13334_ _13193_/A _13193_/C _13193_/B vssd1 vssd1 vccd1 vccd1 _13335_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14505__B _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15697__A2 _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16053_ _16054_/A _16054_/B vssd1 vssd1 vccd1 vccd1 _16226_/B sky130_fd_sc_hd__or2_1
XFILLER_0_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13265_ _13265_/A _13265_/B vssd1 vssd1 vccd1 vccd1 _13266_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11707__A1 _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15004_ _15004_/A _15004_/B _15004_/C vssd1 vssd1 vccd1 vccd1 _15006_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_122_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12216_ _12269_/A _12214_/C _12246_/C _12245_/B vssd1 vssd1 vccd1 vccd1 _12217_/C
+ sky130_fd_sc_hd__a22oi_2
X_13196_ _13196_/A _13196_/B _13196_/C vssd1 vssd1 vccd1 vccd1 _13199_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_20_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18635__A2 _19732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20523__A _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17843__B1 _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19812_ _19810_/D _20178_/B _10798_/Y _19650_/D vssd1 vssd1 vccd1 vccd1 _19813_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_12147_ _12141_/A _12141_/B _12141_/C vssd1 vssd1 vccd1 vccd1 _12148_/C sky130_fd_sc_hd__a21o_1
XANTENNA__20242__B _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19743_ _19743_/A _19743_/B _19743_/C vssd1 vssd1 vccd1 vccd1 _19743_/X sky130_fd_sc_hd__and3_1
X_16955_ _16890_/Y _16947_/X _16945_/Y _16946_/A vssd1 vssd1 vccd1 vccd1 _16956_/C
+ sky130_fd_sc_hd__a211o_1
X_12078_ _12079_/A _12079_/B vssd1 vssd1 vccd1 vccd1 _12078_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__18399__A1 _21791_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18399__B2 _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11356__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15906_ _16151_/A _15906_/B vssd1 vssd1 vccd1 vccd1 _15907_/C sky130_fd_sc_hd__xnor2_1
X_11029_ mstream_o[103] hold309/X _11039_/S vssd1 vssd1 vccd1 vccd1 hold310/A sky130_fd_sc_hd__mux2_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16886_ _17124_/C _16882_/X _16935_/A _16935_/B vssd1 vssd1 vccd1 vccd1 _16888_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_19674_ _19671_/X _19672_/Y _19512_/B _19514_/B vssd1 vssd1 vccd1 vccd1 _19675_/B
+ sky130_fd_sc_hd__o211ai_1
X_15837_ _15837_/A _15966_/A vssd1 vssd1 vccd1 vccd1 _15841_/A sky130_fd_sc_hd__or2_1
X_18625_ _18625_/A _18625_/B vssd1 vssd1 vccd1 vccd1 _18628_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_95_1196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12976__A _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15768_ _15768_/A _16177_/B vssd1 vssd1 vccd1 vccd1 _15769_/B sky130_fd_sc_hd__nand2_1
XANTENNA__21155__B1 _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18556_ _18553_/Y _18709_/A _19185_/D _19201_/B vssd1 vssd1 vccd1 vccd1 _18709_/B
+ sky130_fd_sc_hd__and4bb_1
XTAP_3490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14719_ _14418_/A _14418_/B _14715_/X _14716_/Y vssd1 vssd1 vccd1 vccd1 _14719_/Y
+ sky130_fd_sc_hd__o211ai_2
X_17507_ _17618_/B _17505_/X _17413_/C _17415_/A vssd1 vssd1 vccd1 vccd1 _17508_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_59_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18487_ _18487_/A _18487_/B vssd1 vssd1 vccd1 vccd1 _18489_/B sky130_fd_sc_hd__or2_1
XFILLER_0_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15699_ _15699_/A _15834_/B vssd1 vssd1 vccd1 vccd1 _15701_/A sky130_fd_sc_hd__or2_2
XFILLER_0_118_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17438_ _17439_/A _17439_/B vssd1 vssd1 vccd1 vccd1 _17536_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__15385__A1 _15386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_15 _11335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_26 _11343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_37 _11430_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_1180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_48 hold247/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17369_ _17369_/A _17369_/B vssd1 vssd1 vccd1 vccd1 _17479_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_43_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_59 hold270/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19108_ _19951_/B _19753_/B _19751_/C _19951_/A vssd1 vssd1 vccd1 vccd1 _19111_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20380_ _20380_/A _20381_/B vssd1 vssd1 vccd1 vccd1 _20788_/A sky130_fd_sc_hd__nor2_4
XANTENNA__14415__B _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16885__A1 _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19039_ _18876_/B _18878_/B _19037_/X _19038_/Y vssd1 vssd1 vccd1 vccd1 _19211_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22050_ _22063_/CLK _22050_/D vssd1 vssd1 vccd1 vccd1 hold290/A sky130_fd_sc_hd__dfxtp_4
XFILLER_0_140_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17726__B _19337_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12736__A2_N _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21001_ _20998_/Y _20999_/X _20865_/Y _20869_/A vssd1 vssd1 vccd1 vccd1 _21001_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19644__D _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14788__D _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout381_A _21773_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout479_A _14217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21394__B1 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21264__A _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21903_ _21938_/CLK hold218/X vssd1 vssd1 vccd1 vccd1 hold217/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11882__B1 _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16358__A _16359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19339__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21834_ _21837_/CLK _21834_/D vssd1 vssd1 vccd1 vccd1 _21834_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21765_ _21767_/CLK _21765_/D vssd1 vssd1 vccd1 vccd1 _21765_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_114_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20716_ _20845_/D _21291_/B _20717_/C _20717_/D vssd1 vssd1 vccd1 vccd1 _20718_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_148_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21696_ _22080_/CLK _21696_/D vssd1 vssd1 vccd1 vccd1 hold152/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13926__A2 _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20647_ hold112/X fanout8/X _20645_/X _11547_/X _20646_/Y vssd1 vssd1 vccd1 vccd1
+ _20647_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_19_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11380_ _11379_/X _17520_/B _11401_/S vssd1 vssd1 vccd1 vccd1 _21798_/D sky130_fd_sc_hd__mux2_1
XANTENNA__16325__B1 _16418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11949__B _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20578_ _20578_/A _20578_/B _20578_/C vssd1 vssd1 vccd1 vccd1 _20712_/B sky130_fd_sc_hd__nor3_4
XFILLER_0_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20046__C _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12771__D _21765_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17917__A _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13050_ _14087_/A _13913_/C _14077_/B _14089_/A vssd1 vssd1 vccd1 vccd1 _13051_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17636__B _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16540__B _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12001_ _12001_/A _12001_/B vssd1 vssd1 vccd1 vccd1 _12003_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__14979__C _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21158__B _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21651__RESET_B _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14698__D _14698_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15173__A1_N _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14060__B _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout360 hold333/X vssd1 vssd1 vccd1 vccd1 _14176_/C sky130_fd_sc_hd__buf_6
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout371 _21775_/Q vssd1 vssd1 vccd1 vccd1 _12402_/B sky130_fd_sc_hd__clkbuf_4
X_16740_ _16698_/A _16698_/B _16698_/C vssd1 vssd1 vccd1 vccd1 _16741_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout382 _21773_/Q vssd1 vssd1 vccd1 vccd1 _13269_/C sky130_fd_sc_hd__clkbuf_4
Xfanout393 _15892_/B vssd1 vssd1 vccd1 vccd1 _15632_/B sky130_fd_sc_hd__clkbuf_8
X_13952_ _13972_/B _13952_/B _13952_/C _13952_/D vssd1 vssd1 vccd1 vccd1 _13952_/Y
+ sky130_fd_sc_hd__nor4_4
XANTENNA__13862__A1 _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21385__B1 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14995__B _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13862__B2 _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17053__A1 _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18467__B _19092_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12903_ _12901_/X _12903_/B vssd1 vssd1 vccd1 vccd1 _12904_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__17053__B2 _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16671_ _16645_/A _16645_/B _16645_/C vssd1 vssd1 vccd1 vccd1 _16672_/C sky130_fd_sc_hd__a21o_1
X_13883_ _13883_/A _13883_/B _13883_/C vssd1 vssd1 vccd1 vccd1 _13884_/C sky130_fd_sc_hd__nand3_2
XANTENNA__16268__A _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15622_ _15483_/Y _15486_/Y _15753_/B _15621_/X vssd1 vssd1 vccd1 vccd1 _15622_/Y
+ sky130_fd_sc_hd__a211oi_2
X_18410_ _18411_/A _18411_/B vssd1 vssd1 vccd1 vccd1 _18410_/Y sky130_fd_sc_hd__nand2_1
X_19390_ _19906_/A _20146_/B _19692_/B _19705_/B vssd1 vssd1 vccd1 vccd1 _19543_/A
+ sky130_fd_sc_hd__nand4_2
X_12834_ _12834_/A _12834_/B vssd1 vssd1 vccd1 vccd1 _12834_/Y sky130_fd_sc_hd__nor2_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18341_ _18341_/A _18341_/B vssd1 vssd1 vccd1 vccd1 _18343_/B sky130_fd_sc_hd__xnor2_2
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15553_ _15669_/A _16396_/A _15808_/C _15553_/D vssd1 vssd1 vccd1 vccd1 _15669_/B
+ sky130_fd_sc_hd__and4b_1
XANTENNA__13404__B _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12765_ _12766_/A _12766_/B _12766_/C vssd1 vssd1 vccd1 vccd1 _12765_/X sky130_fd_sc_hd__a21o_4
XFILLER_0_90_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18553__A1 _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_336 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14504_ _16087_/A _15695_/A _14817_/C _14817_/D vssd1 vssd1 vccd1 vccd1 _14504_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__18553__B2 _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15900__A _16031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15367__A1 _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18272_ _18273_/A _18273_/B vssd1 vssd1 vccd1 vccd1 _18272_/X sky130_fd_sc_hd__or2_1
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ _11716_/A _11716_/B vssd1 vssd1 vccd1 vccd1 _11718_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__15367__B2 _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15484_ _15484_/A _15484_/B vssd1 vssd1 vccd1 vccd1 _15487_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12696_ _12716_/B _12697_/B _12697_/C _12697_/D vssd1 vssd1 vccd1 vccd1 _12696_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17223_ _17223_/A _19432_/A vssd1 vssd1 vccd1 vccd1 _17227_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14435_ _14435_/A _14435_/B vssd1 vssd1 vccd1 vccd1 _14438_/A sky130_fd_sc_hd__xor2_2
X_11647_ _12319_/C _12420_/D _12403_/A _12511_/A vssd1 vssd1 vccd1 vccd1 _11648_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_4_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14516__A _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17154_ _17120_/X _17136_/Y _17137_/Y _17153_/X vssd1 vssd1 vccd1 vccd1 _17154_/X
+ sky130_fd_sc_hd__o22a_1
X_14366_ _14367_/A _16286_/A _14367_/C _14513_/A vssd1 vssd1 vccd1 vccd1 _14368_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11859__B _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18856__A2 _19181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11578_ _12619_/A _11577_/X _11576_/X vssd1 vssd1 vccd1 vccd1 _11579_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_141_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16105_ _16305_/B _16399_/A _16396_/B _16418_/B vssd1 vssd1 vccd1 vccd1 _16212_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_123_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16867__A1 _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13317_ _13318_/A _13318_/B vssd1 vssd1 vccd1 vccd1 _13451_/B sky130_fd_sc_hd__nand2_2
XANTENNA__16867__B2 _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17085_ _17066_/A _17066_/C _17066_/B vssd1 vssd1 vccd1 vccd1 _17091_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_126_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14297_ _21725_/D hold118/X _10881_/X fanout6/X vssd1 vssd1 vccd1 vccd1 _14297_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16036_ _16036_/A _16036_/B vssd1 vssd1 vccd1 vccd1 _16038_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13248_ _13249_/A _13249_/B vssd1 vssd1 vccd1 vccd1 _13248_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_58_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21349__A _21349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11875__A _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20415__A2 _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13179_ _13179_/A _13179_/B vssd1 vssd1 vccd1 vccd1 _13199_/A sky130_fd_sc_hd__xor2_2
X_17987_ _17987_/A _17987_/B vssd1 vssd1 vccd1 vccd1 _17989_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11086__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19726_ _19847_/A _19592_/X _19847_/B _19844_/C vssd1 vssd1 vccd1 vccd1 _19726_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__21376__A0 _14296_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16938_ _17029_/A _17029_/B _17124_/C _17145_/B vssd1 vssd1 vccd1 vccd1 _16938_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_79_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19657_ _19658_/A _19658_/B vssd1 vssd1 vccd1 vccd1 _19659_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_79_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16869_ _17013_/C _16868_/X _16867_/X vssd1 vssd1 vccd1 vccd1 _16871_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_133_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18608_ _18608_/A _18608_/B _18608_/C vssd1 vssd1 vccd1 vccd1 _18608_/Y sky130_fd_sc_hd__nand3_2
X_19588_ _19587_/A _19587_/B _20247_/D vssd1 vssd1 vccd1 vccd1 _19723_/C sky130_fd_sc_hd__o21a_2
XFILLER_0_133_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18539_ hold94/X fanout8/X _18537_/Y _11550_/A _18538_/Y vssd1 vssd1 vccd1 vccd1
+ _18539_/X sky130_fd_sc_hd__a221o_1
XANTENNA__19489__A _19650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18544__A1 _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18544__B2 _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15358__A1 _12291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21550_ mstream_o[13] hold31/X _21562_/S vssd1 vssd1 vccd1 vccd1 _22077_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_47_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20501_ _20355_/C _20355_/Y _20499_/Y _20500_/X vssd1 vssd1 vccd1 vccd1 _20501_/Y
+ sky130_fd_sc_hd__a211oi_4
X_21481_ hold178/X sstream_i[58] _21481_/S vssd1 vssd1 vccd1 vccd1 _22008_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13419__A2_N _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20432_ _21171_/A _21153_/B _20430_/Y _20558_/A vssd1 vssd1 vccd1 vccd1 _20434_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_71_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20363_ _20363_/A _20363_/B vssd1 vssd1 vccd1 vccd1 _20366_/A sky130_fd_sc_hd__and2_1
XFILLER_0_28_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16976__A2_N _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22102_ _22105_/CLK _22102_/D _11089_/A vssd1 vssd1 vccd1 vccd1 mstream_o[38] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_28_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20294_ _20294_/A _20294_/B _20294_/C vssd1 vssd1 vccd1 vccd1 _20295_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_101_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout596_A _21349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12344__A1 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22033_ _22038_/CLK _22033_/D vssd1 vssd1 vccd1 vccd1 hold246/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16086__A2 _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12647__A2 _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10880_ _10880_/A _10880_/B _10878_/Y vssd1 vssd1 vccd1 vccd1 _10881_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_156_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21817_ _21817_/CLK _21817_/D vssd1 vssd1 vccd1 vccd1 _21817_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ _13013_/A _12899_/B vssd1 vssd1 vccd1 vccd1 _12554_/A sky130_fd_sc_hd__nand2_1
X_21748_ _22005_/CLK _21748_/D vssd1 vssd1 vccd1 vccd1 _21748_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_66_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11501_ _11507_/A1 t1y[17] t0x[17] _11501_/B2 vssd1 vssd1 vccd1 vccd1 _11501_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_53_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12481_ _12379_/B _12379_/Y _12479_/Y _12480_/X vssd1 vssd1 vccd1 vccd1 _12481_/Y
+ sky130_fd_sc_hd__a211oi_1
X_21679_ _21682_/CLK _21679_/D vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_151_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14220_ _14220_/A _14220_/B _14220_/C vssd1 vssd1 vccd1 vccd1 _14222_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_151_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11432_ _11447_/A1 hold119/A fanout48/X hold178/A vssd1 vssd1 vccd1 vccd1 _11432_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20772__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11679__B _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14055__B _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14151_ _14148_/X _14149_/Y _13985_/D _13986_/B vssd1 vssd1 vccd1 vccd1 _14168_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_81_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11363_ _11124_/A hold230/X _11126_/B hold196/X vssd1 vssd1 vccd1 vccd1 _11363_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13102_ _13102_/A _13102_/B _13102_/C vssd1 vssd1 vccd1 vccd1 _13103_/B sky130_fd_sc_hd__or3_1
XANTENNA__21169__A _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14082_ _14713_/B _15098_/B vssd1 vssd1 vccd1 vccd1 _14086_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14324__A2 _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11294_ _11493_/A1 t1x[17] v2z[17] _11507_/B2 _11293_/X vssd1 vssd1 vccd1 vccd1 _11294_/X
+ sky130_fd_sc_hd__a221o_2
X_13033_ _14716_/A _13034_/D _12906_/X _12907_/X _14384_/C vssd1 vssd1 vccd1 vccd1
+ _13038_/A sky130_fd_sc_hd__a32o_1
X_17910_ _17910_/A _17910_/B _17910_/C vssd1 vssd1 vccd1 vccd1 _17912_/A sky130_fd_sc_hd__nand3_2
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18890_ _18889_/B _18889_/C _18889_/A vssd1 vssd1 vccd1 vccd1 _18987_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__12886__A2 _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17841_ _17594_/A _17595_/A _17837_/X _17839_/X vssd1 vssd1 vccd1 vccd1 _17841_/Y
+ sky130_fd_sc_hd__o31ai_4
XANTENNA__14088__A1 _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18909__C _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14984_ _14984_/A _14984_/B _14984_/C vssd1 vssd1 vccd1 vccd1 _14984_/Y sky130_fd_sc_hd__nand3_1
X_17772_ _17772_/A _17891_/B _17772_/C vssd1 vssd1 vccd1 vccd1 _17772_/Y sky130_fd_sc_hd__nand3_4
Xfanout190 _18498_/B vssd1 vssd1 vccd1 vccd1 _19123_/B sky130_fd_sc_hd__buf_4
XANTENNA__12638__A2 _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20520__B _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19511_ _19510_/B _19661_/B _19510_/A vssd1 vssd1 vccd1 vccd1 _19512_/C sky130_fd_sc_hd__a21o_1
X_13935_ _13784_/A _13784_/C _13784_/B vssd1 vssd1 vccd1 vccd1 _13936_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_88_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16723_ _16723_/A _16723_/B vssd1 vssd1 vccd1 vccd1 _16792_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_88_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19971__B1 _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16654_ _16653_/A _16653_/Y _16633_/X _16635_/Y vssd1 vssd1 vccd1 vccd1 _16657_/C
+ sky130_fd_sc_hd__a211oi_4
X_19442_ _19291_/A _19291_/B _19440_/X _19441_/Y vssd1 vssd1 vccd1 vccd1 _19444_/A
+ sky130_fd_sc_hd__o211a_1
X_13866_ _13867_/A _16273_/A _13867_/C _13867_/D vssd1 vssd1 vccd1 vccd1 _13866_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_92_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15605_ _15605_/A _15605_/B _15605_/C vssd1 vssd1 vccd1 vccd1 _15693_/B sky130_fd_sc_hd__or3_2
XFILLER_0_92_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12817_ _12816_/A _12816_/B _12816_/C vssd1 vssd1 vccd1 vccd1 _12818_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16585_ _17178_/A _16583_/Y _16532_/A _16534_/B vssd1 vssd1 vccd1 vccd1 _16657_/B
+ sky130_fd_sc_hd__o211a_1
X_19373_ _19529_/B _19373_/B _20265_/D vssd1 vssd1 vccd1 vccd1 _19373_/X sky130_fd_sc_hd__and3_1
XFILLER_0_69_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13797_ _13643_/C _13642_/Y _13795_/X _13796_/Y vssd1 vssd1 vccd1 vccd1 _13800_/C
+ sky130_fd_sc_hd__o211a_2
XANTENNA__11580__D _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14134__A2_N _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15536_ _15791_/A _15916_/B _16424_/A _16040_/C vssd1 vssd1 vccd1 vccd1 _15663_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_85_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18324_ _18324_/A _18324_/B vssd1 vssd1 vccd1 vccd1 _18326_/B sky130_fd_sc_hd__xor2_1
XANTENNA__21530__A0 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ _12630_/B _12631_/Y _12837_/A _12747_/X vssd1 vssd1 vccd1 vccd1 _12837_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_139_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16445__B _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18255_ _19185_/D _19199_/C _19199_/D _19008_/D vssd1 vssd1 vccd1 vccd1 _18255_/Y
+ sky130_fd_sc_hd__a22oi_1
X_15467_ _15327_/Y _15332_/A _15465_/X _15466_/Y vssd1 vssd1 vccd1 vccd1 _15469_/B
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_115_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12679_ _12679_/A _12679_/B _12679_/C vssd1 vssd1 vccd1 vccd1 _12681_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13150__A _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17206_ _17619_/A _17206_/B vssd1 vssd1 vccd1 vccd1 _17210_/A sky130_fd_sc_hd__nand2_1
X_14418_ _14418_/A _14418_/B vssd1 vssd1 vccd1 vccd1 _14419_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_115_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15760__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18186_ _18062_/A _18061_/B _18061_/A vssd1 vssd1 vccd1 vccd1 _18193_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__11589__B _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15398_ _16305_/B _16369_/A _15398_/C _15398_/D vssd1 vssd1 vccd1 vccd1 _15541_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__15760__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17137_ _17134_/Y _17135_/X _17130_/B vssd1 vssd1 vccd1 vccd1 _17137_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_123_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14349_ _14176_/C _14348_/X _14347_/X vssd1 vssd1 vccd1 vccd1 _14351_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__17557__A _17557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17501__A2 _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15512__A1 _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17068_ _17068_/A _17068_/B _17068_/C vssd1 vssd1 vccd1 vccd1 _17071_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_111_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16019_ _15756_/A _16016_/B _16016_/C vssd1 vssd1 vccd1 vccd1 _16019_/X sky130_fd_sc_hd__o21ba_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15508__C _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20133__D _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11755__D _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13826__A1 _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17723__C _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13826__B2 _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17280__A4 _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19709_ _19708_/B _19708_/C _19708_/A vssd1 vssd1 vccd1 vccd1 _19711_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_100_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20981_ _20981_/A _20981_/B vssd1 vssd1 vccd1 vccd1 _20983_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout177_A _21826_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13325__A _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_1206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13044__B _14712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout344_A _14477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16636__A _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21602_ _21888_/CLK _21602_/D _11041_/A vssd1 vssd1 vccd1 vccd1 mstream_o[65] sky130_fd_sc_hd__dfrtp_4
XANTENNA__18554__C _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21521__A0 hold239/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21261__B _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12262__B1 _21727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16528__B1 _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21533_ hold306/X sstream_i[110] _21536_/S vssd1 vssd1 vccd1 vccd1 _22060_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_7_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout511_A _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout609_A _21718_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17740__A2 _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19666__B _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21464_ hold199/X sstream_i[41] _21494_/S vssd1 vssd1 vccd1 vccd1 _21991_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20415_ _20416_/B _20924_/A _21305_/A _20416_/A vssd1 vssd1 vccd1 vccd1 _20419_/C
+ sky130_fd_sc_hd__a22o_1
X_21395_ hold38/X fanout40/X _21393_/Y _21394_/Y vssd1 vssd1 vccd1 vccd1 _21939_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16371__A _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12107__C _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20346_ _20199_/Y _20201_/X _20344_/X _20345_/Y vssd1 vssd1 vccd1 vccd1 _20498_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_101_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16521__D _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20277_ _20277_/A _20277_/B vssd1 vssd1 vccd1 vccd1 _20279_/B sky130_fd_sc_hd__xor2_1
X_22016_ _22016_/CLK _22016_/D vssd1 vssd1 vccd1 vccd1 hold176/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11981_ _11971_/A _11971_/B _11971_/C vssd1 vssd1 vccd1 vccd1 _11982_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13293__A2 _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13720_ _13720_/A _13720_/B vssd1 vssd1 vccd1 vccd1 _13729_/A sky130_fd_sc_hd__or2_1
X_10932_ _10923_/B _10925_/Y _10931_/Y vssd1 vssd1 vccd1 vccd1 _10940_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__15153__C _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13651_ _13648_/X _13649_/Y _13496_/C _13495_/Y vssd1 vssd1 vccd1 vccd1 _13652_/D
+ sky130_fd_sc_hd__a211oi_2
X_10863_ hold133/A hold115/A vssd1 vssd1 vccd1 vccd1 _10873_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_156_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13045__A2 _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12602_ _21725_/D hold125/A _11051_/Y fanout6/X _12601_/Y vssd1 vssd1 vccd1 vccd1
+ _12602_/X sky130_fd_sc_hd__a221o_1
X_16370_ _16370_/A _16370_/B vssd1 vssd1 vccd1 vccd1 _16373_/A sky130_fd_sc_hd__xor2_1
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21171__B _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13582_ _13581_/A _13581_/B _13568_/X vssd1 vssd1 vccd1 vccd1 _13582_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_94_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10794_ _16286_/A vssd1 vssd1 vccd1 vccd1 _10794_/Y sky130_fd_sc_hd__inv_2
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15321_ _15318_/Y _15450_/A _15838_/D _15978_/B vssd1 vssd1 vccd1 vccd1 _15450_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_87_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19279__D _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12533_ _12637_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _12537_/A sky130_fd_sc_hd__nand2_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18040_ _18040_/A _18164_/A _18040_/C vssd1 vssd1 vccd1 vccd1 _18164_/B sky130_fd_sc_hd__nand3_2
X_15252_ _15252_/A _15252_/B vssd1 vssd1 vccd1 vccd1 _15292_/A sky130_fd_sc_hd__xnor2_1
X_12464_ _12463_/A _12463_/B _12463_/C vssd1 vssd1 vccd1 vccd1 _12465_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_136_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14203_ _14203_/A _14203_/B _14203_/C vssd1 vssd1 vccd1 vccd1 _14203_/X sky130_fd_sc_hd__and3_1
XFILLER_0_2_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11415_ hold235/A fanout28/X _11414_/X vssd1 vssd1 vccd1 vccd1 _11415_/X sky130_fd_sc_hd__a21o_1
X_15183_ _14956_/X _14958_/Y _15331_/B _15182_/Y vssd1 vssd1 vccd1 vccd1 _15296_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12395_ _11667_/B _11666_/A _11666_/B _12317_/A _12314_/X vssd1 vssd1 vccd1 vccd1
+ _12484_/A sky130_fd_sc_hd__a41o_1
XFILLER_0_151_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14134_ _14133_/D _16406_/B _16374_/B _13983_/B vssd1 vssd1 vccd1 vccd1 _14135_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_11346_ _11544_/A1 t1x[30] v2z[30] _11543_/B2 _11345_/X vssd1 vssd1 vccd1 vccd1 _11346_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__17096__B _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19991_ _19991_/A _19991_/B vssd1 vssd1 vccd1 vccd1 _20000_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14065_ _14064_/A _14064_/B _14064_/C vssd1 vssd1 vccd1 vccd1 _14066_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_24_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18942_ _18942_/A _19084_/B _18942_/C vssd1 vssd1 vccd1 vccd1 _18944_/B sky130_fd_sc_hd__nand3_2
X_11277_ _11325_/A1 t2y[13] t0y[13] _11498_/A1 vssd1 vssd1 vccd1 vccd1 _11277_/X sky130_fd_sc_hd__a22o_1
XANTENNA__12859__A2 _13269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13016_ _13016_/A _13016_/B vssd1 vssd1 vccd1 vccd1 _13025_/A sky130_fd_sc_hd__xor2_1
X_18873_ _18873_/A _21847_/Q _18873_/C _19028_/A vssd1 vssd1 vccd1 vccd1 _19028_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17824_ _17824_/A _17824_/B vssd1 vssd1 vccd1 vccd1 _17825_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_20_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__21346__B _21346_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17543__C _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14967_ _14967_/A _14967_/B vssd1 vssd1 vccd1 vccd1 _14968_/B sky130_fd_sc_hd__xnor2_1
X_17755_ _17852_/A _17753_/Y _17630_/B _17630_/Y vssd1 vssd1 vccd1 vccd1 _17815_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__18747__A1 _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20003__B1 _19868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16706_ _16676_/A _16676_/B _16676_/C vssd1 vssd1 vccd1 vccd1 _16706_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_57_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13918_ _13916_/X _13918_/B vssd1 vssd1 vccd1 vccd1 _13919_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_57_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14898_ _14747_/A _14747_/B _14745_/Y vssd1 vssd1 vccd1 vccd1 _14900_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_89_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17686_ _17570_/B _17570_/Y _17683_/X _17685_/Y vssd1 vssd1 vccd1 vccd1 _17689_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_49_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19425_ _19424_/B _19424_/C _19406_/X vssd1 vssd1 vccd1 vccd1 _19426_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_58_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13849_ _13689_/Y _13692_/X _13847_/Y _13848_/X vssd1 vssd1 vccd1 vccd1 _13973_/A
+ sky130_fd_sc_hd__a211oi_2
X_16637_ _17145_/A _17433_/A vssd1 vssd1 vccd1 vccd1 _16639_/B sky130_fd_sc_hd__and2_1
XANTENNA__14233__A1 _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14233__B2 _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19356_ _19356_/A _19356_/B _19356_/C vssd1 vssd1 vccd1 vccd1 _19358_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_91_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16568_ _17636_/B _17490_/A vssd1 vssd1 vccd1 vccd1 _16572_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11598__A2 _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18307_ _18183_/B _18183_/Y _18305_/Y _18306_/X vssd1 vssd1 vccd1 vccd1 _18307_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_155_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15519_ _15519_/A _15519_/B vssd1 vssd1 vccd1 vccd1 _15521_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__16606__D _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16499_ _17277_/A _17739_/C _17739_/D _17387_/A vssd1 vssd1 vccd1 vccd1 _16549_/A
+ sky130_fd_sc_hd__and4_1
X_19287_ _20247_/C _19117_/X _19286_/X vssd1 vssd1 vccd1 vccd1 _19289_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18238_ _18386_/B _18235_/X _18095_/B _18095_/Y vssd1 vssd1 vccd1 vccd1 _18239_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__20128__D _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13311__C _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18169_ _18169_/A _18169_/B vssd1 vssd1 vccd1 vccd1 _18179_/A sky130_fd_sc_hd__and2_1
XFILLER_0_142_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20200_ _20200_/A _20200_/B vssd1 vssd1 vccd1 vccd1 _20202_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_123_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21180_ _21259_/A _21180_/B vssd1 vssd1 vccd1 vccd1 _21182_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11539__S _11545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20131_ _20131_/A _20330_/B vssd1 vssd1 vccd1 vccd1 _20142_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_110_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20062_ _20167_/B _20060_/X _19919_/X _19921_/Y vssd1 vssd1 vccd1 vccd1 _20062_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout294_A _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21256__B _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20793__A1 _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout461_A _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout559_A _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_308 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_319 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20964_ _20964_/A _20964_/B vssd1 vssd1 vccd1 vccd1 _21012_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20895_ _20895_/A _20895_/B vssd1 vssd1 vccd1 vccd1 _20898_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11038__A1 hold277/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12786__A1 _12785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12786__B2 _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17174__B1 _11553_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18581__A _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18910__A1 _19379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21516_ hold236/X sstream_i[93] _21528_/S vssd1 vssd1 vccd1 vccd1 _22043_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12538__A1 _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16813__B _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21447_ hold296/X sstream_i[24] _21489_/S vssd1 vssd1 vccd1 vccd1 _21974_/D sky130_fd_sc_hd__mux2_1
XANTENNA__20335__B _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11200_ hold130/X fanout22/X _11199_/X vssd1 vssd1 vccd1 vccd1 _11200_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_82_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21273__A2 _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12180_ _12269_/A _12245_/B _12512_/A _12214_/C vssd1 vssd1 vccd1 vccd1 _12183_/A
+ sky130_fd_sc_hd__nand4_2
X_21378_ hold57/X _21381_/B vssd1 vssd1 vccd1 vccd1 _21378_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__13875__D _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11449__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11131_ hold213/X fanout23/X _11130_/X vssd1 vssd1 vccd1 vccd1 _11131_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_82_1198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20329_ _20329_/A _20329_/B vssd1 vssd1 vccd1 vccd1 _20340_/A sky130_fd_sc_hd__or2_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20989__C _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18426__B1 _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11062_ _11061_/X hold40/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21660_/D sky130_fd_sc_hd__mux2_1
X_15870_ _15870_/A vssd1 vssd1 vccd1 vccd1 _15870_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16988__B1 _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14821_ _14662_/X _14665_/X _14818_/X _14820_/Y vssd1 vssd1 vccd1 vccd1 _14821_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11692__B _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14752_ _14592_/A _14592_/B _14590_/Y vssd1 vssd1 vccd1 vccd1 _14754_/B sky130_fd_sc_hd__a21boi_4
XANTENNA__11277__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17540_ _21802_/Q _19432_/A _17436_/B _17434_/X vssd1 vssd1 vccd1 vccd1 _17550_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_3864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11964_ _11964_/A _11964_/B _11969_/C _11964_/D vssd1 vssd1 vccd1 vccd1 _11964_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12300__C _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13703_ _13819_/A _13702_/C _13702_/A vssd1 vssd1 vccd1 vccd1 _13804_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_86_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10915_ hold205/A hold89/A vssd1 vssd1 vccd1 vccd1 _10924_/A sky130_fd_sc_hd__and2_1
XFILLER_0_86_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17471_ _17487_/B _17470_/B _17468_/Y _17469_/X vssd1 vssd1 vccd1 vccd1 _17471_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_129_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14683_ _14682_/A _14682_/B _14682_/C vssd1 vssd1 vccd1 vccd1 _14684_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11895_ _11872_/Y _11892_/X _11893_/X _11830_/Y vssd1 vssd1 vccd1 vccd1 _11901_/A
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_128_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11029__A1 hold309/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19210_ _19363_/B _19210_/B vssd1 vssd1 vccd1 vccd1 _19213_/A sky130_fd_sc_hd__nand2b_1
X_16422_ _16422_/A _16422_/B vssd1 vssd1 vccd1 vccd1 _16423_/B sky130_fd_sc_hd__xnor2_1
X_13634_ _13480_/A _13480_/C _13480_/B vssd1 vssd1 vccd1 vccd1 _13635_/C sky130_fd_sc_hd__a21bo_1
X_10846_ hold315/A hold122/A _10845_/X vssd1 vssd1 vccd1 vccd1 _11065_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15963__B2 _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16353_ _16354_/A _16354_/B vssd1 vssd1 vccd1 vccd1 _16353_/X sky130_fd_sc_hd__or2_1
XANTENNA__13974__B1 _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19141_ _18979_/B _18979_/Y _19139_/Y _19140_/X vssd1 vssd1 vccd1 vccd1 _19143_/B
+ sky130_fd_sc_hd__o211ai_4
X_13565_ _13565_/A _13565_/B vssd1 vssd1 vccd1 vccd1 _13567_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_109_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15304_ _15306_/A _15437_/B vssd1 vssd1 vccd1 vccd1 _15307_/A sky130_fd_sc_hd__or2_1
XFILLER_0_82_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19072_ _19071_/B _19235_/B _19071_/A vssd1 vssd1 vccd1 vccd1 _19073_/C sky130_fd_sc_hd__a21o_1
X_12516_ _12517_/A _12517_/B vssd1 vssd1 vccd1 vccd1 _12629_/A sky130_fd_sc_hd__nand2_1
X_16284_ _16284_/A _16284_/B vssd1 vssd1 vccd1 vccd1 _16286_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_82_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13496_ _13496_/A _13496_/B _13496_/C _13496_/D vssd1 vssd1 vccd1 vccd1 _13496_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_87_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18405__A1_N _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12529__A1 _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15235_ _15375_/A _15368_/D _15233_/Y _15377_/A vssd1 vssd1 vccd1 vccd1 _15237_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_81_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18023_ _18020_/X _18021_/Y _17910_/B _17912_/A vssd1 vssd1 vccd1 vccd1 _18023_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12529__B2 _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12447_ _12447_/A _12447_/B vssd1 vssd1 vccd1 vccd1 _12449_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_140_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15166_ _15166_/A _15166_/B vssd1 vssd1 vccd1 vccd1 _15167_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_10_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12378_ _12375_/X _12376_/Y _11776_/C _11775_/Y vssd1 vssd1 vccd1 vccd1 _12379_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11359__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14117_ _14117_/A _14117_/B _14117_/C vssd1 vssd1 vccd1 vccd1 _14280_/B sky130_fd_sc_hd__or3_1
XFILLER_0_50_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11329_ _11349_/A1 t2y[26] t0y[26] _11089_/B vssd1 vssd1 vccd1 vccd1 _11329_/X sky130_fd_sc_hd__a22o_1
X_15097_ _15375_/A _15098_/B _15098_/C _15238_/A vssd1 vssd1 vccd1 vccd1 _15097_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19974_ _20650_/A _20242_/C _19974_/C _20110_/A vssd1 vssd1 vccd1 vccd1 _20110_/B
+ sky130_fd_sc_hd__nand4_2
X_14048_ _14174_/B _14046_/Y _13906_/X _13943_/A vssd1 vssd1 vccd1 vccd1 _14048_/Y
+ sky130_fd_sc_hd__a211oi_2
X_18925_ _18925_/A _18925_/B vssd1 vssd1 vccd1 vccd1 _18944_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18856_ _19008_/D _19181_/B _19185_/B _18857_/B vssd1 vssd1 vccd1 vccd1 _18859_/C
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__20775__A1 _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_98_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17807_ _17684_/B _17684_/Y _17804_/X _17806_/Y vssd1 vssd1 vccd1 vccd1 _17810_/B
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__20411__D _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18787_ _18787_/A _18787_/B _21040_/A _19866_/C vssd1 vssd1 vccd1 vccd1 _18947_/A
+ sky130_fd_sc_hd__nand4_2
X_15999_ _15999_/A _15999_/B _15999_/C _15999_/D vssd1 vssd1 vccd1 vccd1 _15999_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_55_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17738_ _18010_/A _18769_/B _17638_/X _17637_/X _18767_/B vssd1 vssd1 vccd1 vccd1
+ _17743_/A sky130_fd_sc_hd__a32o_1
XANTENNA__20527__A1 _20249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17669_ _17669_/A _17669_/B vssd1 vssd1 vccd1 vccd1 _17678_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17720__D _18894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19408_ _20101_/B _19906_/C _19906_/D _20101_/A vssd1 vssd1 vccd1 vccd1 _19408_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20680_ _20681_/A _20681_/B vssd1 vssd1 vccd1 vccd1 _20872_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_46_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13313__A1_N _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19339_ _18849_/B _20178_/B _21261_/B _18851_/C vssd1 vssd1 vccd1 vccd1 _19340_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_70_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11123__A _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11440__A1 _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21301_ _21301_/A _21816_/Q vssd1 vssd1 vccd1 vccd1 _21303_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17448__C _17924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout307_A _21794_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21232_ _21232_/A _21232_/B vssd1 vssd1 vccd1 vccd1 _21234_/B sky130_fd_sc_hd__or2_1
Xhold210 hold210/A vssd1 vssd1 vccd1 vccd1 hold210/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold221 hold221/A vssd1 vssd1 vccd1 vccd1 hold221/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold232 hold232/A vssd1 vssd1 vccd1 vccd1 hold232/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold243 hold243/A vssd1 vssd1 vccd1 vccd1 hold243/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20463__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold254 hold254/A vssd1 vssd1 vccd1 vccd1 hold254/X sky130_fd_sc_hd__dlygate4sd3_1
X_21163_ _21163_/A _21163_/B vssd1 vssd1 vccd1 vccd1 _21164_/A sky130_fd_sc_hd__xor2_1
Xhold265 hold265/A vssd1 vssd1 vccd1 vccd1 hold265/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 hold276/A vssd1 vssd1 vccd1 vccd1 hold276/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 hold287/A vssd1 vssd1 vccd1 vccd1 hold287/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold298 hold298/A vssd1 vssd1 vccd1 vccd1 hold298/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__21267__A _21267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20114_ _20114_/A _20114_/B vssd1 vssd1 vccd1 vccd1 _20116_/B sky130_fd_sc_hd__xor2_2
X_21094_ _21095_/B vssd1 vssd1 vccd1 vccd1 _21094_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_102_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18279__C _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20045_ _20845_/D _20733_/C _20606_/D _20721_/D vssd1 vssd1 vccd1 vccd1 _20045_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11259__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_105 _21800_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_116 sstream_i[69] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21996_ _22021_/CLK _21996_/D vssd1 vssd1 vccd1 vccd1 hold198/A sky130_fd_sc_hd__dfxtp_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18295__B _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18187__A2 _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_127 v0z[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_138 v1z[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16198__A1 _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20947_ _20946_/B _20946_/C _20946_/A vssd1 vssd1 vccd1 vccd1 _20948_/B sky130_fd_sc_hd__a21o_1
XANTENNA_149 v1z[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ _12109_/C _12750_/A _11680_/C _11705_/A vssd1 vssd1 vccd1 vccd1 _11705_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20878_ _20877_/B _20877_/C _20877_/A vssd1 vssd1 vccd1 vccd1 _20880_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_49_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14328__B _15174_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13350_ _13209_/C _13208_/Y _13348_/X _13349_/Y vssd1 vssd1 vccd1 vccd1 _13353_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11431__A1 _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ _12511_/A _12858_/C _12991_/D _12402_/A vssd1 vssd1 vccd1 vccd1 _12302_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13281_ _13280_/A _13280_/B _13266_/Y vssd1 vssd1 vccd1 vccd1 _13281_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_84_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15020_ _15791_/A _16196_/B _16371_/A _16196_/A vssd1 vssd1 vccd1 vccd1 _15024_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12232_ _12232_/A _12232_/B vssd1 vssd1 vccd1 vccd1 _12234_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11687__B _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15159__B _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14920__A2 _14918_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13174__A2_N _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19854__B _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11195__A0 _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18111__A2 _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12163_ _12154_/A _12154_/B _12156_/X vssd1 vssd1 vccd1 vccd1 _12165_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14998__B _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11114_ _10946_/Y hold43/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21708_/D sky130_fd_sc_hd__mux2_1
X_16971_ _16971_/A _16971_/B _16971_/C vssd1 vssd1 vccd1 vccd1 _17018_/A sky130_fd_sc_hd__nand3_1
X_12094_ _12094_/A _12094_/B _12512_/A _12214_/C vssd1 vssd1 vccd1 vccd1 _12094_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_120_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18710_ _18873_/A _19199_/C _19199_/D _19493_/D vssd1 vssd1 vccd1 vccd1 _18713_/C
+ sky130_fd_sc_hd__a22o_1
X_15922_ _15923_/A _15923_/B vssd1 vssd1 vccd1 vccd1 _16114_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__18189__C _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11045_ _11045_/A _11045_/B vssd1 vssd1 vccd1 vccd1 _11045_/X sky130_fd_sc_hd__xor2_4
XANTENNA__17093__C _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19690_ _19692_/B _19692_/C _20416_/B _19535_/A vssd1 vssd1 vccd1 vccd1 _19695_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18641_ _18641_/A _18641_/B _18784_/B vssd1 vssd1 vccd1 vccd1 _18641_/X sky130_fd_sc_hd__and3_1
X_15853_ _16084_/A _15978_/B _15851_/Y _15972_/A vssd1 vssd1 vccd1 vccd1 _15855_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__18486__A _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__B _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14804_ _14804_/A _14804_/B vssd1 vssd1 vccd1 vccd1 _14806_/B sky130_fd_sc_hd__xnor2_1
X_18572_ _18572_/A _18572_/B _18572_/C vssd1 vssd1 vccd1 vccd1 _18572_/X sky130_fd_sc_hd__or3_1
XFILLER_0_8_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15784_ _15784_/A _15784_/B vssd1 vssd1 vccd1 vccd1 _15823_/A sky130_fd_sc_hd__nand2_1
XTAP_3650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12996_ _13128_/B _12995_/C _12995_/A vssd1 vssd1 vccd1 vccd1 _12997_/C sky130_fd_sc_hd__a21o_1
XTAP_3661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17523_ _17619_/A _17636_/B _17522_/C _17522_/D vssd1 vssd1 vccd1 vccd1 _17524_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14735_ _14735_/A _14735_/B vssd1 vssd1 vccd1 vccd1 _14738_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_8_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11947_ _12426_/B _12302_/A _11876_/Y _11878_/B vssd1 vssd1 vccd1 vccd1 _11948_/B
+ sky130_fd_sc_hd__a22oi_1
XTAP_3694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14666_ _15695_/A _15022_/B _14666_/C _14666_/D vssd1 vssd1 vccd1 vccd1 _14666_/Y
+ sky130_fd_sc_hd__nand4_1
XTAP_2993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17454_ _17453_/A _17453_/B _17453_/C vssd1 vssd1 vccd1 vccd1 _17455_/C sky130_fd_sc_hd__a21o_1
X_11878_ _11879_/A _11878_/B _12426_/B _12302_/A vssd1 vssd1 vccd1 vccd1 _11948_/A
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_55_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11746__A1_N _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16405_ _16372_/A _16294_/A _16294_/B _16296_/Y vssd1 vssd1 vccd1 vccd1 _16407_/A
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_129_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13617_ _13618_/A _13618_/B vssd1 vssd1 vccd1 vccd1 _13758_/B sky130_fd_sc_hd__and2b_1
X_10829_ hold206/A hold223/A vssd1 vssd1 vccd1 vccd1 _10830_/B sky130_fd_sc_hd__or2_1
X_14597_ _14443_/A _14443_/B _14441_/Y vssd1 vssd1 vccd1 vccd1 _14599_/B sky130_fd_sc_hd__a21oi_1
X_17385_ _17282_/A _20797_/A _21258_/A _17277_/A vssd1 vssd1 vccd1 vccd1 _17386_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19124_ _19123_/A _19123_/B _20247_/D vssd1 vssd1 vccd1 vccd1 _19126_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_54_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11422__A1 _21311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16336_ _16337_/A _16337_/B _16337_/C vssd1 vssd1 vccd1 vccd1 _16388_/B sky130_fd_sc_hd__a21o_1
X_13548_ _13548_/A vssd1 vssd1 vccd1 vccd1 _13548_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_6_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16267_ _16414_/B _16266_/X _16265_/X vssd1 vssd1 vccd1 vccd1 _16269_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_124_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19055_ _19382_/A _19057_/C _19057_/D _19529_/B vssd1 vssd1 vccd1 vccd1 _19060_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13479_ _13478_/A _13478_/B _13478_/C vssd1 vssd1 vccd1 vccd1 _13480_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_124_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15218_ _15218_/A _15218_/B _15361_/B vssd1 vssd1 vccd1 vccd1 _15218_/X sky130_fd_sc_hd__and3_1
X_18006_ _18006_/A _18006_/B vssd1 vssd1 vccd1 vccd1 _18014_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11597__B _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16198_ _16374_/A _16404_/B _16199_/C _16199_/D vssd1 vssd1 vccd1 vccd1 _16200_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__11186__A0 _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15149_ _15013_/X _15050_/X _15147_/X _15148_/X vssd1 vssd1 vccd1 vccd1 _15151_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_50_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19957_ _19956_/B _20087_/B _20091_/A vssd1 vssd1 vccd1 vccd1 _19958_/C sky130_fd_sc_hd__a21o_1
XANTENNA__14675__A1 _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18908_ _19535_/A _20103_/A _19068_/C _19695_/A vssd1 vssd1 vccd1 vccd1 _18911_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11489__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19602__A2 _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19888_ _19883_/Y _19885_/X _19743_/X _19763_/X vssd1 vssd1 vccd1 vccd1 _19923_/B
+ sky130_fd_sc_hd__a211oi_1
X_18839_ _18839_/A _18839_/B vssd1 vssd1 vccd1 vccd1 _18839_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12221__B _12242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_5_clk_i _21806_/CLK vssd1 vssd1 vccd1 vccd1 _21803_/CLK sky130_fd_sc_hd__clkbuf_16
X_21850_ _21853_/CLK _21850_/D vssd1 vssd1 vccd1 vccd1 hold329/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__14978__A2 _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20801_ _20801_/A _20801_/B vssd1 vssd1 vccd1 vccd1 _20801_/X sky130_fd_sc_hd__or2_1
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21781_ _21821_/CLK _21781_/D vssd1 vssd1 vccd1 vccd1 hold241/A sky130_fd_sc_hd__dfxtp_2
XANTENNA__11110__A0 _10919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17916__A2 _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20732_ _20735_/D vssd1 vssd1 vccd1 vccd1 _20732_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_77_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20663_ _20918_/A _20664_/B vssd1 vssd1 vccd1 vccd1 _20788_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_19_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout424_A _12771_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11413__A1 _20991_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20594_ _20594_/A _20594_/B vssd1 vssd1 vccd1 vccd1 _20597_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__18190__A2_N _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19955__A _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11177__A0 _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21215_ _21216_/A _21216_/B vssd1 vssd1 vccd1 vccd1 _21215_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_143_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20987__A1 _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20987__B2 _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21146_ _21034_/B _21146_/B vssd1 vssd1 vccd1 vccd1 _21146_/X sky130_fd_sc_hd__and2b_1
XANTENNA__13469__A2 _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout520 _14024_/B vssd1 vssd1 vccd1 vccd1 _13017_/A sky130_fd_sc_hd__buf_4
Xfanout531 _13864_/B vssd1 vssd1 vccd1 vccd1 _12877_/A sky130_fd_sc_hd__clkbuf_4
Xfanout542 _21735_/Q vssd1 vssd1 vccd1 vccd1 _13858_/A sky130_fd_sc_hd__clkbuf_8
X_21077_ _21077_/A _21077_/B _21077_/C vssd1 vssd1 vccd1 vccd1 _21232_/A sky130_fd_sc_hd__and3_1
Xfanout553 _13554_/B vssd1 vssd1 vccd1 vccd1 _12530_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout72_A _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout564 _12621_/C vssd1 vssd1 vccd1 vccd1 _12403_/A sky130_fd_sc_hd__buf_4
Xfanout575 _21728_/Q vssd1 vssd1 vccd1 vccd1 _12268_/B sky130_fd_sc_hd__buf_4
XANTENNA__17604__A1 _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout586 _21718_/D vssd1 vssd1 vccd1 vccd1 _11447_/A1 sky130_fd_sc_hd__buf_4
Xfanout597 _11122_/A vssd1 vssd1 vccd1 vccd1 _21349_/A sky130_fd_sc_hd__buf_4
XANTENNA__17604__B2 _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20028_ _20025_/Y _20175_/A _20178_/D _20841_/B vssd1 vssd1 vccd1 vccd1 _20175_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_38_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12850_ _12984_/B _12850_/B vssd1 vssd1 vccd1 vccd1 _12853_/A sky130_fd_sc_hd__or2_1
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11801_ _11801_/A _11801_/B _11801_/C vssd1 vssd1 vccd1 vccd1 _11801_/X sky130_fd_sc_hd__or3_2
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ _12779_/Y _12780_/X _13173_/C _12781_/D vssd1 vssd1 vccd1 vccd1 _12783_/A
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__11101__A0 _10852_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21979_ _22013_/CLK _21979_/D vssd1 vssd1 vccd1 vccd1 hold175/A sky130_fd_sc_hd__dfxtp_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14520_ _14519_/B _14671_/B _14519_/A vssd1 vssd1 vccd1 vccd1 _14521_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_95_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12785__C _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11732_ _11732_/A _11732_/B _11732_/C vssd1 vssd1 vccd1 vccd1 _11744_/A sky130_fd_sc_hd__nand3_1
XANTENNA__15918__A1 _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14058__B _14218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18580__A2 _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14451_ hold243/X _14450_/X fanout3/X vssd1 vssd1 vccd1 vccd1 _21870_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11663_ _11664_/A _11664_/B vssd1 vssd1 vccd1 vccd1 _11666_/A sky130_fd_sc_hd__or2_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16554__A _21825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13402_ _13554_/B _13556_/A _13858_/C _13402_/D vssd1 vssd1 vccd1 vccd1 _13404_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_153_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17170_ _16962_/X _17164_/X _17169_/X vssd1 vssd1 vccd1 vccd1 _17171_/B sky130_fd_sc_hd__a21o_2
XANTENNA__11404__A1 _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14382_ _14240_/A _14239_/B _14237_/X vssd1 vssd1 vccd1 vccd1 _14398_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11594_ _11610_/A _11610_/B _11610_/C vssd1 vssd1 vccd1 vccd1 _11833_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_24_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16121_ _16119_/B _16119_/C _16119_/A vssd1 vssd1 vccd1 vccd1 _16121_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__16273__B _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13333_ _13332_/B _13332_/C _13332_/A vssd1 vssd1 vccd1 vccd1 _13335_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16052_ _16052_/A _16052_/B vssd1 vssd1 vccd1 vccd1 _16054_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_49_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13264_ _13411_/B _13263_/B _13263_/C vssd1 vssd1 vccd1 vccd1 _13265_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__11168__A0 _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15003_ _15000_/Y _15001_/X _14878_/D _14878_/Y vssd1 vssd1 vccd1 vccd1 _15004_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__11707__A2 _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12215_ _12268_/A _12246_/D vssd1 vssd1 vccd1 vccd1 _12217_/B sky130_fd_sc_hd__nand2_1
X_13195_ _13056_/A _13056_/C _13056_/B vssd1 vssd1 vccd1 vccd1 _13196_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__18635__A3 _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20523__B _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19811_ _19813_/A vssd1 vssd1 vccd1 vccd1 _20041_/A sky130_fd_sc_hd__inv_2
X_12146_ _12146_/A _12146_/B vssd1 vssd1 vccd1 vccd1 _12148_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20242__C _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13418__A _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19742_ _19743_/A _19743_/B _19743_/C vssd1 vssd1 vccd1 vccd1 _19742_/Y sky130_fd_sc_hd__a21oi_1
X_16954_ _16954_/A _16954_/B vssd1 vssd1 vccd1 vccd1 _16956_/B sky130_fd_sc_hd__xnor2_1
X_12077_ _12077_/A _12077_/B vssd1 vssd1 vccd1 vccd1 _12079_/B sky130_fd_sc_hd__xor2_1
XANTENNA__12668__B1 _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18399__A2 _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15905_ _15905_/A _15905_/B vssd1 vssd1 vccd1 vccd1 _15906_/B sky130_fd_sc_hd__nand2_2
X_11028_ mstream_o[102] hold275/X _11039_/S vssd1 vssd1 vccd1 vccd1 _21639_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_155_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19673_ _19512_/B _19514_/B _19671_/X _19672_/Y vssd1 vssd1 vccd1 vccd1 _19673_/Y
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__11340__A0 _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16885_ _17124_/C _16882_/X _16884_/X vssd1 vssd1 vccd1 vccd1 _16935_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18624_ _18624_/A _19089_/B _18624_/C _18624_/D vssd1 vssd1 vccd1 vccd1 _18625_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__18647__C _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15836_ _15835_/B _15836_/B vssd1 vssd1 vccd1 vccd1 _15966_/A sky130_fd_sc_hd__and2b_1
XANTENNA__13681__A2_N _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12976__B _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18555_ _19185_/D _19201_/B _18553_/Y _18709_/A vssd1 vssd1 vccd1 vccd1 _18555_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_63_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15767_ _15767_/A _15767_/B vssd1 vssd1 vccd1 vccd1 _15769_/A sky130_fd_sc_hd__nor2_1
XTAP_3480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21155__A1 _21841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12979_ _13975_/B _14018_/C vssd1 vssd1 vccd1 vccd1 _12983_/A sky130_fd_sc_hd__nand2_1
XTAP_3491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21155__B2 _21267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17506_ _17413_/C _17415_/A _17618_/B _17505_/X vssd1 vssd1 vccd1 vccd1 _17629_/A
+ sky130_fd_sc_hd__a211o_1
X_14718_ _14418_/A _14418_/B _14715_/X _14716_/Y vssd1 vssd1 vccd1 vccd1 _14718_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12840__B1 _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18486_ _20088_/A _19703_/C _18486_/C _18486_/D vssd1 vssd1 vccd1 vccd1 _18487_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_74_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15698_ _15838_/D _15698_/B _15698_/C _15698_/D vssd1 vssd1 vccd1 vccd1 _15834_/B
+ sky130_fd_sc_hd__and4_1
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17437_ _17437_/A _17437_/B vssd1 vssd1 vccd1 vccd1 _17439_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14649_ _14649_/A _14649_/B vssd1 vssd1 vccd1 vccd1 _14650_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_28_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_16 _11335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16464__A _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_27 _11343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_38 _11436_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_49 hold247/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17368_ _17369_/A _17369_/B vssd1 vssd1 vccd1 vccd1 _17590_/A sky130_fd_sc_hd__and2_1
XFILLER_0_32_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_938 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19107_ _19587_/B _20242_/C _18957_/X _18958_/X _20242_/D vssd1 vssd1 vccd1 vccd1
+ _19112_/A sky130_fd_sc_hd__a32o_1
X_16319_ _16319_/A _16319_/B vssd1 vssd1 vccd1 vccd1 _16321_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17299_ _17296_/A _17297_/Y _17190_/Y _17193_/X vssd1 vssd1 vccd1 vccd1 _17360_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_43_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19038_ _19037_/B _19037_/C _19037_/A vssd1 vssd1 vccd1 vccd1 _19038_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11159__A0 _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20714__A _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14712__A _14712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17726__C _19692_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20433__B _21283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21000_ _20865_/Y _20869_/A _20998_/Y _20999_/X vssd1 vssd1 vccd1 vccd1 _21000_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_10_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15309__A1_N _21735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_37_clk_i_A clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout374_A _21775_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21394__A1 _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11331__B1 _11330_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21902_ _21934_/CLK hold253/X vssd1 vssd1 vccd1 vccd1 hold252/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__21264__B _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19015__A _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__A1 _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__B2 _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16270__B1 _21755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19339__B2 _18851_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21833_ _21837_/CLK _21833_/D vssd1 vssd1 vccd1 vccd1 _21833_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_78_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout541_A _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout639_A _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18011__A1 _18010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21764_ _21767_/CLK _21764_/D vssd1 vssd1 vccd1 vccd1 _21764_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20715_ _20843_/A vssd1 vssd1 vccd1 vccd1 _20717_/D sky130_fd_sc_hd__inv_2
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16374__A _16374_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21695_ _22080_/CLK _21695_/D vssd1 vssd1 vccd1 vccd1 hold49/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20608__B _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20646_ _21142_/A _21404_/B vssd1 vssd1 vccd1 vccd1 _20646_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_34_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16325__A1 _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16325__B2 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11949__C _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20577_ _20574_/X _20575_/Y _20441_/B _20442_/Y vssd1 vssd1 vccd1 vccd1 _20578_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20046__D _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17917__B _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12843__A2_N _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12898__B1 _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12000_ _11992_/A _11994_/B _11992_/B vssd1 vssd1 vccd1 vccd1 _12003_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__14979__D _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11570__B1 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21129_ _21129_/A _21129_/B vssd1 vssd1 vccd1 vccd1 _21131_/B sky130_fd_sc_hd__or2_1
Xfanout350 _16377_/A vssd1 vssd1 vccd1 vccd1 _15913_/B sky130_fd_sc_hd__buf_2
XANTENNA__14060__C _14873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout361 _16369_/A vssd1 vssd1 vccd1 vccd1 _15022_/B sky130_fd_sc_hd__clkbuf_4
Xfanout372 _21775_/Q vssd1 vssd1 vccd1 vccd1 _15808_/C sky130_fd_sc_hd__buf_4
Xfanout383 _16173_/A vssd1 vssd1 vccd1 vccd1 _14516_/A sky130_fd_sc_hd__clkbuf_8
X_13951_ _13948_/X _13949_/Y _13800_/C _13799_/Y vssd1 vssd1 vccd1 vccd1 _13952_/D
+ sky130_fd_sc_hd__a211oi_2
Xfanout394 _21771_/Q vssd1 vssd1 vccd1 vccd1 _15892_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__21385__A1 _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13862__A2 _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12902_ _13032_/B _12900_/X _12780_/X _12783_/A vssd1 vssd1 vccd1 vccd1 _12903_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__17053__A2 _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18467__C _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13882_ _13883_/A _13883_/B _13883_/C vssd1 vssd1 vccd1 vccd1 _13884_/B sky130_fd_sc_hd__a21o_2
X_16670_ _16669_/B _16669_/C _16669_/A vssd1 vssd1 vccd1 vccd1 _16672_/B sky130_fd_sc_hd__a21bo_1
X_15621_ _15753_/A _15619_/X _15445_/Y _15448_/Y vssd1 vssd1 vccd1 vccd1 _15621_/X
+ sky130_fd_sc_hd__o211a_1
X_12833_ _12834_/A _12834_/B vssd1 vssd1 vccd1 vccd1 _12969_/A sky130_fd_sc_hd__and2_2
XFILLER_0_9_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11192__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18340_ _18341_/B _18341_/A vssd1 vssd1 vccd1 vccd1 _18478_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_68_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15552_ _15808_/C _16396_/A _15550_/Y _15669_/A vssd1 vssd1 vccd1 vccd1 _15554_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_115_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12764_ _12764_/A _12764_/B vssd1 vssd1 vccd1 vccd1 _12766_/C sky130_fd_sc_hd__xnor2_2
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_495 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21190__A _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18553__A2 _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19750__A1 _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14503_ _16203_/D _14354_/C _14817_/D _15695_/A vssd1 vssd1 vccd1 vccd1 _14508_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19750__B2 _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11715_ _11716_/A _11716_/B vssd1 vssd1 vccd1 vccd1 _12336_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15483_ _15484_/B _15484_/A vssd1 vssd1 vccd1 vccd1 _15483_/Y sky130_fd_sc_hd__nand2b_1
X_18271_ _18703_/A _19013_/C vssd1 vssd1 vccd1 vccd1 _18273_/B sky130_fd_sc_hd__nand2_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ _12692_/X _12693_/Y _12583_/C _12582_/Y vssd1 vssd1 vccd1 vccd1 _12697_/D
+ sky130_fd_sc_hd__a211o_2
XANTENNA__16284__A _16284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13378__A1 _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17222_ _16604_/A _16603_/A _16603_/B vssd1 vssd1 vccd1 vccd1 _17229_/A sky130_fd_sc_hd__o21ba_1
X_14434_ _14434_/A _14434_/B vssd1 vssd1 vccd1 vccd1 _14435_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_25_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11646_ _12319_/C _12403_/A _12511_/A _12420_/D vssd1 vssd1 vccd1 vccd1 _11648_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__14516__B _14828_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14365_ _14365_/A _14516_/A _14365_/C _14365_/D vssd1 vssd1 vccd1 vccd1 _14513_/A
+ sky130_fd_sc_hd__nand4_2
X_17153_ _17130_/B _17134_/Y _17135_/X _17152_/Y vssd1 vssd1 vccd1 vccd1 _17153_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_123_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11577_ _12020_/A _12326_/D _14621_/D vssd1 vssd1 vccd1 vccd1 _11577_/X sky130_fd_sc_hd__and3_1
XANTENNA__11859__C _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16104_ _16107_/D vssd1 vssd1 vccd1 vccd1 _16104_/Y sky130_fd_sc_hd__inv_2
X_13316_ _13316_/A _13316_/B vssd1 vssd1 vccd1 vccd1 _13318_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_24_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17084_ _17071_/A _17071_/C _17071_/B vssd1 vssd1 vccd1 vccd1 _17101_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_123_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14296_ _14601_/C _14296_/B vssd1 vssd1 vccd1 vccd1 _14296_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_40_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16035_ _16035_/A _16035_/B vssd1 vssd1 vccd1 vccd1 _16036_/B sky130_fd_sc_hd__nand2_1
X_13247_ _13400_/A _13247_/B vssd1 vssd1 vccd1 vccd1 _13249_/B sky130_fd_sc_hd__nor2_1
XANTENNA__21349__B _21349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13178_ _13179_/A _13179_/B vssd1 vssd1 vccd1 vccd1 _13304_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11875__B _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12129_ _12130_/A _12130_/B vssd1 vssd1 vccd1 vccd1 _12129_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_97_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17986_ _18121_/A _18127_/B vssd1 vssd1 vccd1 vccd1 _17987_/B sky130_fd_sc_hd__nor2_1
X_19725_ _19291_/A _19291_/B _19722_/X _19723_/Y vssd1 vssd1 vccd1 vccd1 _19844_/C
+ sky130_fd_sc_hd__o211ai_2
X_16937_ _16937_/A _16937_/B vssd1 vssd1 vccd1 vccd1 _16943_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__21376__A1 _19169_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11864__A1 _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19656_ _19656_/A _19656_/B vssd1 vssd1 vccd1 vccd1 _19658_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16868_ _16868_/A _17129_/B _16968_/C vssd1 vssd1 vccd1 vccd1 _16868_/X sky130_fd_sc_hd__and3_1
XANTENNA__11864__B2 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18607_ _18608_/A _18608_/B _18608_/C vssd1 vssd1 vccd1 vccd1 _18607_/X sky130_fd_sc_hd__and3_1
X_15819_ _15642_/Y _15644_/Y _15817_/A _15818_/Y vssd1 vssd1 vccd1 vccd1 _15819_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_133_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19587_ _19587_/A _19587_/B _21056_/B vssd1 vssd1 vccd1 vccd1 _19723_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_87_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16799_ _16727_/A _16727_/C _16727_/B vssd1 vssd1 vccd1 vccd1 _16800_/C sky130_fd_sc_hd__a21o_1
X_18538_ _21142_/A _21364_/B vssd1 vssd1 vccd1 vccd1 _18538_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_133_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19489__B _20841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18544__A2 _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15358__A2 _15356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18469_ _18466_/Y _18626_/A _19535_/A _18624_/A vssd1 vssd1 vccd1 vccd1 _18626_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_74_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13611__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20500_ _20499_/A _20499_/B _20499_/C _20499_/D vssd1 vssd1 vccd1 vccd1 _20500_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_145_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21480_ hold207/X sstream_i[57] _21481_/S vssd1 vssd1 vccd1 vccd1 _22007_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20431_ _21056_/A _21169_/A _21264_/B _21046_/B vssd1 vssd1 vccd1 vccd1 _20558_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_99_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout122_A _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21938_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_43_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20362_ _20359_/Y _20360_/X _20214_/X _20217_/Y vssd1 vssd1 vccd1 vccd1 _20363_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22101_ _22105_/CLK _22101_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[37] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20293_ _20294_/A _20294_/B _20294_/C vssd1 vssd1 vccd1 vccd1 _20449_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_140_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22032_ _22038_/CLK _22032_/D vssd1 vssd1 vccd1 vccd1 hold281/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12344__A2 _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout491_A _21746_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11552__B1 _21329_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_38_clk_i clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21837_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__18849__A _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout589_A _11549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19009__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20975__A_N _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20147__A2_N _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__A0 _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12897__A _21743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16369__A _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18584__A _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21816_ _21816_/CLK _21816_/D vssd1 vssd1 vccd1 vccd1 _21816_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__11607__A1 _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout35_A _21490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21747_ _22005_/CLK _21747_/D vssd1 vssd1 vccd1 vccd1 _21747_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14617__A _14774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11500_ _11499_/X _19238_/C _11521_/S vssd1 vssd1 vccd1 vccd1 _21838_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18113__A1_N _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12480_ _12479_/A _12479_/B _12479_/C _12479_/D vssd1 vssd1 vccd1 vccd1 _12480_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_65_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21678_ _21939_/CLK _21678_/D vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout1_A fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11431_ _11430_/X _21264_/B _11470_/S vssd1 vssd1 vccd1 vccd1 _21815_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_11_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12152__A2_N _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20629_ _20628_/A _20628_/B _20627_/C _20627_/D vssd1 vssd1 vccd1 vccd1 _20629_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_105_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12137__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11679__C _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14055__C _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14150_ _13985_/D _13986_/B _14148_/X _14149_/Y vssd1 vssd1 vccd1 vccd1 _14301_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12782__A2_N _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11362_ _11361_/X _17145_/B _11401_/S vssd1 vssd1 vccd1 vccd1 _21792_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_22_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13101_ _13102_/A _13102_/B _13102_/C vssd1 vssd1 vccd1 vccd1 _13243_/A sky130_fd_sc_hd__o21ai_2
X_14081_ _14081_/A _14081_/B vssd1 vssd1 vccd1 vccd1 _14101_/A sky130_fd_sc_hd__xnor2_2
X_11293_ _11325_/A1 t2y[17] t0y[17] _11498_/A1 vssd1 vssd1 vccd1 vccd1 _11293_/X sky130_fd_sc_hd__a22o_1
X_13032_ _13032_/A _13032_/B vssd1 vssd1 vccd1 vccd1 _13040_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_120_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17840_ _17594_/A _17595_/A _17837_/X _17839_/X vssd1 vssd1 vccd1 vccd1 _17969_/A
+ sky130_fd_sc_hd__o31a_2
XFILLER_0_28_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14088__A2 hold313/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17771_ _17891_/A _17770_/C _17770_/A vssd1 vssd1 vccd1 vccd1 _17772_/C sky130_fd_sc_hd__a21o_1
X_14983_ _14982_/B _15075_/B _15218_/A vssd1 vssd1 vccd1 vccd1 _14984_/C sky130_fd_sc_hd__a21o_1
Xfanout180 _21826_/Q vssd1 vssd1 vccd1 vccd1 _17443_/D sky130_fd_sc_hd__buf_4
XANTENNA__18909__D _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 _17557_/B vssd1 vssd1 vccd1 vccd1 _18498_/B sky130_fd_sc_hd__clkbuf_4
X_19510_ _19510_/A _19510_/B _19661_/B vssd1 vssd1 vccd1 vccd1 _19512_/B sky130_fd_sc_hd__nand3_2
XANTENNA__20520__C _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16722_ _16721_/B _16721_/C _16721_/A vssd1 vssd1 vccd1 vccd1 _16723_/B sky130_fd_sc_hd__a21oi_1
X_13934_ _13933_/B _13933_/C _13933_/A vssd1 vssd1 vccd1 vccd1 _13936_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_135_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19441_ _19441_/A _19441_/B _19441_/C vssd1 vssd1 vccd1 vccd1 _19441_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__19971__A1 _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16653_ _16653_/A _16653_/B _16653_/C vssd1 vssd1 vccd1 vccd1 _16653_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__19971__B2 _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13865_ _13867_/A _16273_/A _13867_/C _13867_/D vssd1 vssd1 vccd1 vccd1 _13865_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15604_ _15601_/Y _15602_/X _15463_/X _15465_/X vssd1 vssd1 vccd1 vccd1 _15605_/C
+ sky130_fd_sc_hd__o211a_1
X_19372_ _19529_/B _21278_/A _20265_/D _19531_/A vssd1 vssd1 vccd1 vccd1 _19372_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12816_ _12816_/A _12816_/B _12816_/C vssd1 vssd1 vccd1 vccd1 _12818_/B sky130_fd_sc_hd__and3_1
X_16584_ _16532_/A _16534_/B _17178_/A _16583_/Y vssd1 vssd1 vccd1 vccd1 _17178_/B
+ sky130_fd_sc_hd__a211oi_4
X_13796_ _13795_/A _13795_/B _13795_/C _13795_/D vssd1 vssd1 vccd1 vccd1 _13796_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18323_ _18324_/A _18324_/B vssd1 vssd1 vccd1 vccd1 _18323_/X sky130_fd_sc_hd__and2_1
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15535_ _15916_/B _16424_/A _16418_/A _15791_/A vssd1 vssd1 vccd1 vccd1 _15539_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ _12744_/Y _12745_/X _12652_/X _12655_/Y vssd1 vssd1 vccd1 vccd1 _12747_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12973__C _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18254_ _19185_/D _19223_/B _18130_/X _18131_/X _18732_/C vssd1 vssd1 vccd1 vccd1
+ _18261_/A sky130_fd_sc_hd__a32oi_2
XFILLER_0_60_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15466_ _15462_/Y _15464_/X _15323_/X _15325_/Y vssd1 vssd1 vccd1 vccd1 _15466_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_127_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12678_ _12567_/A _12567_/C _12567_/B vssd1 vssd1 vccd1 vccd1 _12679_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_72_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17205_ _17281_/B _17205_/B vssd1 vssd1 vccd1 vccd1 _17215_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_5_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14417_ _14572_/B _14251_/B _14572_/A vssd1 vssd1 vccd1 vccd1 _14418_/B sky130_fd_sc_hd__mux2_4
XANTENNA__13150__B _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11629_ _12229_/A _12155_/B _12751_/B _12637_/B vssd1 vssd1 vccd1 vccd1 _11683_/A
+ sky130_fd_sc_hd__nand4_2
X_18185_ _18185_/A _18185_/B vssd1 vssd1 vccd1 vccd1 _18195_/A sky130_fd_sc_hd__or2_1
X_15397_ _16305_/B _16369_/A _15398_/C _15398_/D vssd1 vssd1 vccd1 vccd1 _15399_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_128_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12047__A _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17136_ _17130_/B _17135_/X _17134_/Y vssd1 vssd1 vccd1 vccd1 _17136_/Y sky130_fd_sc_hd__a21boi_1
X_14348_ _14659_/A _15435_/A _15112_/D vssd1 vssd1 vccd1 vccd1 _14348_/X sky130_fd_sc_hd__and3_1
XANTENNA__17557__B _17557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14279_ _14279_/A _14279_/B vssd1 vssd1 vccd1 vccd1 _14282_/A sky130_fd_sc_hd__or2_2
X_17067_ _17066_/B _17066_/C _17066_/A vssd1 vssd1 vccd1 vccd1 _17068_/C sky130_fd_sc_hd__a21bo_1
X_16018_ _15625_/A _15622_/Y _15624_/B vssd1 vssd1 vccd1 vccd1 _16018_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17969_ _17969_/A _18243_/A vssd1 vssd1 vccd1 vccd1 _17970_/B sky130_fd_sc_hd__nand2_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13826__A2 _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17723__D _19053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15093__A _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19708_ _19708_/A _19708_/B _19708_/C vssd1 vssd1 vccd1 vccd1 _19711_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20980_ _20849_/A _20848_/A _20848_/B _20844_/B _20844_/A vssd1 vssd1 vccd1 vccd1
+ _20981_/B sky130_fd_sc_hd__o32ai_4
XFILLER_0_79_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13325__B _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19639_ _19499_/A _19499_/B _19502_/A vssd1 vssd1 vccd1 vccd1 _19782_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_149_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14787__B1 _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13044__C _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16636__B _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21601_ _21888_/CLK _21601_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[64] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16528__A1 _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18554__D _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16528__B2 _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout337_A _21784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21532_ hold262/X sstream_i[109] _21536_/S vssd1 vssd1 vccd1 vccd1 _22059_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14539__B1 _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21463_ hold183/X sstream_i[40] _21494_/S vssd1 vssd1 vccd1 vccd1 _21990_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_141_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout504_A _21743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13762__A1 _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20414_ _20414_/A _20603_/B vssd1 vssd1 vccd1 vccd1 _20425_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21394_ _21720_/D _15210_/B _21381_/B vssd1 vssd1 vccd1 vccd1 _21394_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__16371__B _21755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12107__D _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20345_ _20341_/Y _20343_/X _20195_/X _20197_/Y vssd1 vssd1 vccd1 vccd1 _20345_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_3_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20276_ _20277_/A _20277_/B vssd1 vssd1 vccd1 vccd1 _20486_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__18579__A _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22015_ _22016_/CLK _22015_/D vssd1 vssd1 vccd1 vccd1 hold197/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_105_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11980_ _12388_/B _11980_/B vssd1 vssd1 vccd1 vccd1 _12294_/B sky130_fd_sc_hd__and2b_1
XANTENNA__12420__A _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ _10931_/A _10931_/B vssd1 vssd1 vccd1 vccd1 _10931_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__17930__B _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15153__D _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13650_ _13496_/C _13495_/Y _13648_/X _13649_/Y vssd1 vssd1 vccd1 vccd1 _13652_/C
+ sky130_fd_sc_hd__o211a_2
X_10862_ hold133/A hold115/A vssd1 vssd1 vccd1 vccd1 _10864_/A sky130_fd_sc_hd__or2_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12601_ fanout9/X _21340_/B vssd1 vssd1 vccd1 vccd1 _12601_/Y sky130_fd_sc_hd__nor2_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13581_ _13581_/A _13581_/B _13568_/X vssd1 vssd1 vccd1 vccd1 _13581_/Y sky130_fd_sc_hd__nor3b_4
XANTENNA__18052__A1_N _19692_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10793_ _16203_/D vssd1 vssd1 vccd1 vccd1 _16314_/B sky130_fd_sc_hd__inv_2
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11470__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15320_ _15838_/D _15978_/B _15318_/Y _15450_/A vssd1 vssd1 vccd1 vccd1 _15322_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_94_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12532_ _12532_/A _12532_/B vssd1 vssd1 vccd1 vccd1 _12542_/A sky130_fd_sc_hd__and2_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_6_clk_i_A _21806_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__22071__RESET_B fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15251_ _15252_/A _15252_/B vssd1 vssd1 vccd1 vccd1 _15251_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_0_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12463_ _12463_/A _12463_/B _12463_/C vssd1 vssd1 vccd1 vccd1 _12465_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_136_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14202_ _14201_/A _14201_/B _14201_/C vssd1 vssd1 vccd1 vccd1 _14203_/C sky130_fd_sc_hd__a21o_1
X_11414_ _11447_/A1 hold267/A fanout47/X hold166/A vssd1 vssd1 vccd1 vccd1 _11414_/X
+ sky130_fd_sc_hd__a22o_1
X_15182_ _15179_/X _15180_/Y _14954_/B _14956_/B vssd1 vssd1 vccd1 vccd1 _15182_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_50_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12394_ hold206/X _12393_/X fanout3/X vssd1 vssd1 vccd1 vccd1 _21855_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18697__A1_N _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14133_ _13381_/C _16406_/B _16314_/D _14133_/D vssd1 vssd1 vccd1 vccd1 _14321_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_50_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11345_ _11349_/A1 t2y[30] t0y[30] _11089_/B vssd1 vssd1 vccd1 vccd1 _11345_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14082__A _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19990_ _20975_/D _20671_/B vssd1 vssd1 vccd1 vccd1 _19991_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_120_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14064_ _14064_/A _14064_/B _14064_/C vssd1 vssd1 vccd1 vccd1 _14209_/A sky130_fd_sc_hd__nand3_1
X_18941_ _19084_/A _18940_/C _18940_/A vssd1 vssd1 vccd1 vccd1 _18942_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_123_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11276_ _12319_/C _11275_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21770_/D sky130_fd_sc_hd__mux2_1
XANTENNA__20812__A _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21579__A1 _11066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13015_ _13152_/C _13013_/X _13014_/X vssd1 vssd1 vccd1 vccd1 _13016_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_123_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18872_ _18873_/A _19199_/D _18873_/C _19028_/A vssd1 vssd1 vccd1 vccd1 _18874_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_990 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17823_ _17824_/A _17824_/B vssd1 vssd1 vccd1 vccd1 _17823_/X sky130_fd_sc_hd__or2_1
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17754_ _17630_/B _17630_/Y _17852_/A _17753_/Y vssd1 vssd1 vccd1 vccd1 _17852_/B
+ sky130_fd_sc_hd__o211ai_4
X_14966_ _14967_/A _14967_/B vssd1 vssd1 vccd1 vccd1 _14966_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__20003__A1 _20562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18747__A2 _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16705_ _16705_/A _16705_/B _16705_/C vssd1 vssd1 vccd1 vccd1 _16705_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__20003__B2 _20689_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20607__A2_N _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13917_ _13916_/B _14073_/B _13916_/A vssd1 vssd1 vccd1 vccd1 _13918_/B sky130_fd_sc_hd__a21o_1
X_17685_ _17684_/B _17684_/C _17684_/A vssd1 vssd1 vccd1 vccd1 _17685_/Y sky130_fd_sc_hd__a21oi_2
X_14897_ _14897_/A _14897_/B vssd1 vssd1 vccd1 vccd1 _14900_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_58_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19424_ _19406_/X _19424_/B _19424_/C vssd1 vssd1 vccd1 vccd1 _19426_/A sky130_fd_sc_hd__nand3b_2
X_16636_ _17146_/A _17146_/B _18166_/A _17434_/B vssd1 vssd1 vccd1 vccd1 _16639_/A
+ sky130_fd_sc_hd__nand4_1
X_13848_ _13845_/Y _13846_/X _13685_/A _13686_/Y vssd1 vssd1 vccd1 vccd1 _13848_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14233__A2 _15091_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19355_ _19354_/B _19504_/B _19354_/A vssd1 vssd1 vccd1 vccd1 _19356_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13441__B1 _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16567_ _16566_/B _16566_/C _16566_/A vssd1 vssd1 vccd1 vccd1 _16582_/A sky130_fd_sc_hd__a21bo_1
X_13779_ _13779_/A _13779_/B _13779_/C vssd1 vssd1 vccd1 vccd1 _13782_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11380__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18306_ _18305_/A _18305_/B _18292_/Y vssd1 vssd1 vccd1 vccd1 _18306_/X sky130_fd_sc_hd__o21ba_1
XFILLER_0_57_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15518_ _15518_/A _15518_/B vssd1 vssd1 vccd1 vccd1 _15519_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19286_ _19587_/B _20249_/B _20247_/C _19587_/A vssd1 vssd1 vccd1 vccd1 _19286_/X
+ sky130_fd_sc_hd__a22o_1
X_16498_ _17277_/A _17739_/C _17739_/D _17387_/A vssd1 vssd1 vccd1 vccd1 _16498_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18237_ _18386_/B _18235_/X _18095_/B _18095_/Y vssd1 vssd1 vccd1 vccd1 _18240_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15449_ _15449_/A _15449_/B vssd1 vssd1 vccd1 vccd1 _15469_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_5_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13311__D _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16472__A _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18168_ _19373_/B _18769_/B _18167_/C _18167_/D vssd1 vssd1 vccd1 vccd1 _18169_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17119_ _17106_/A _17106_/C _17106_/B vssd1 vssd1 vccd1 vccd1 _17120_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_141_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18099_ _18241_/A _18099_/B vssd1 vssd1 vccd1 vccd1 _18100_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_29_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20179__A1_N _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20130_ _20838_/B _20671_/B _20130_/C _20330_/A vssd1 vssd1 vccd1 vccd1 _20330_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_111_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_96_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21723__RESET_B fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_99_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20061_ _19919_/X _19921_/Y _20167_/B _20060_/X vssd1 vssd1 vccd1 vccd1 _20216_/A
+ sky130_fd_sc_hd__a211oi_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20793__A2 _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout287_A _21798_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_309 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20963_ _20960_/X _20961_/Y _20790_/B _20830_/Y vssd1 vssd1 vccd1 vccd1 _20964_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_136_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout454_A hold313/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15551__A _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20894_ _20895_/A _20895_/B vssd1 vssd1 vccd1 vccd1 _20894_/X sky130_fd_sc_hd__or2_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout621_A _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12786__A2 _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18581__B _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21515_ hold245/X sstream_i[92] _21528_/S vssd1 vssd1 vccd1 vccd1 _22042_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_17_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18910__A2 _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16813__C _17063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12538__A2 _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21446_ hold291/X sstream_i[23] _21489_/S vssd1 vssd1 vccd1 vccd1 _21973_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_1107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20335__C _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21377_ hold118/X _21376_/X _21403_/S vssd1 vssd1 vccd1 vccd1 _21933_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_32_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11130_ hold224/X _11126_/A _11126_/B hold197/X vssd1 vssd1 vccd1 vccd1 _11130_/X
+ sky130_fd_sc_hd__a22o_1
X_20328_ _20328_/A _20328_/B vssd1 vssd1 vccd1 vccd1 _20348_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_101_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11061_ _11061_/A _11061_/B vssd1 vssd1 vccd1 vccd1 _11061_/X sky130_fd_sc_hd__xor2_4
XANTENNA__18426__A1 _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20989__D _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18426__B2 _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20259_ _20260_/B _20260_/C _20260_/A vssd1 vssd1 vccd1 vccd1 _20259_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__18102__A _19636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16988__A1 _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16988__B2 _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14820_ _16203_/D _15022_/B _14820_/C _14820_/D vssd1 vssd1 vccd1 vccd1 _14820_/Y
+ sky130_fd_sc_hd__nand4_1
XANTENNA__11692__C _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15660__A1 _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14751_ _14751_/A _14751_/B vssd1 vssd1 vccd1 vccd1 _14754_/A sky130_fd_sc_hd__xnor2_4
XTAP_3854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11963_ _11969_/C _11964_/D vssd1 vssd1 vccd1 vccd1 _12027_/B sky130_fd_sc_hd__nor2_1
XTAP_3865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18248__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13702_ _13702_/A _13819_/A _13702_/C vssd1 vssd1 vccd1 vccd1 _13819_/B sky130_fd_sc_hd__nor3_1
XANTENNA__12300__D _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10914_ hold205/A hold89/A vssd1 vssd1 vccd1 vccd1 _10916_/A sky130_fd_sc_hd__nor2_1
X_17470_ _17487_/B _17470_/B _17468_/Y _17469_/X vssd1 vssd1 vccd1 vccd1 _17470_/X
+ sky130_fd_sc_hd__or4bb_4
X_14682_ _14682_/A _14682_/B _14682_/C vssd1 vssd1 vccd1 vccd1 _14809_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11894_ _11872_/Y _11892_/X _11893_/X _11830_/Y vssd1 vssd1 vccd1 vccd1 _11894_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_86_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16421_ _16421_/A _16421_/B vssd1 vssd1 vccd1 vccd1 _16422_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13633_ _13632_/B _13632_/C _13632_/A vssd1 vssd1 vccd1 vccd1 _13635_/B sky130_fd_sc_hd__a21o_1
X_10845_ hold315/A hold122/A hold219/A hold58/A vssd1 vssd1 vccd1 vccd1 _10845_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19868__A _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14077__A _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18772__A _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19140_ _19139_/B _19139_/C _19139_/A vssd1 vssd1 vccd1 vccd1 _19140_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_67_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16352_ _16352_/A _16352_/B vssd1 vssd1 vccd1 vccd1 _16354_/B sky130_fd_sc_hd__and2_1
XANTENNA__13974__A1 _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13564_ _13565_/A _13565_/B vssd1 vssd1 vccd1 vccd1 _13690_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_27_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11985__B1 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15303_ _15439_/D _15698_/B _15303_/C _15303_/D vssd1 vssd1 vccd1 vccd1 _15437_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__21402__S _21407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19071_ _19071_/A _19071_/B _19235_/B vssd1 vssd1 vccd1 vccd1 _19073_/B sky130_fd_sc_hd__nand3_1
X_12515_ _12515_/A _12515_/B vssd1 vssd1 vccd1 vccd1 _12517_/B sky130_fd_sc_hd__xnor2_2
X_16283_ _16283_/A vssd1 vssd1 vccd1 vccd1 _16286_/C sky130_fd_sc_hd__inv_2
X_13495_ _13496_/A _13496_/B _13496_/C _13496_/D vssd1 vssd1 vccd1 vccd1 _13495_/Y
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_48_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21249__B1 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18022_ _17910_/B _17912_/A _18020_/X _18021_/Y vssd1 vssd1 vccd1 vccd1 _18107_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12529__A2 _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15234_ _15373_/A _15373_/B _15234_/C _16286_/B vssd1 vssd1 vccd1 vccd1 _15377_/A
+ sky130_fd_sc_hd__and4_1
X_12446_ _12444_/X _12446_/B vssd1 vssd1 vccd1 vccd1 _12447_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_112_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15165_ _15166_/A _15166_/B vssd1 vssd1 vccd1 vccd1 _15165_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12377_ _11776_/C _11775_/Y _12375_/X _12376_/Y vssd1 vssd1 vccd1 vccd1 _12379_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__12325__A _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14116_ _14113_/X _14114_/X _13952_/C _13952_/Y vssd1 vssd1 vccd1 vccd1 _14117_/C
+ sky130_fd_sc_hd__a211oi_1
X_11328_ _14635_/D _11327_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21783_/D sky130_fd_sc_hd__mux2_1
X_15096_ _15373_/A _15373_/B _15368_/D _15234_/C vssd1 vssd1 vccd1 vccd1 _15238_/A
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_61_1239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19973_ _20650_/A _20242_/C _19974_/C _20110_/A vssd1 vssd1 vccd1 vccd1 _19973_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20542__A _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10960__A1 _10959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18924_ _19007_/A _18922_/Y _18758_/B _18758_/Y vssd1 vssd1 vccd1 vccd1 _18983_/B
+ sky130_fd_sc_hd__o211a_1
X_14047_ _13906_/X _13943_/A _14174_/B _14046_/Y vssd1 vssd1 vccd1 vccd1 _14132_/A
+ sky130_fd_sc_hd__o211a_1
X_11259_ fanout59/X v0z[8] fanout19/X _11258_/X vssd1 vssd1 vccd1 vccd1 _11259_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__14540__A _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12979__B _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18855_ _18855_/A _18855_/B vssd1 vssd1 vccd1 vccd1 _18863_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_98_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20775__A2 _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17806_ _17805_/B _17805_/C _17805_/A vssd1 vssd1 vccd1 vccd1 _17806_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18786_ _18787_/B _21040_/A _19866_/C _18787_/A vssd1 vssd1 vccd1 vccd1 _18789_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15998_ _16134_/A _15996_/C _15996_/A vssd1 vssd1 vccd1 vccd1 _15999_/D sky130_fd_sc_hd__a21oi_1
XANTENNA__21373__A _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17737_ _17737_/A _17737_/B vssd1 vssd1 vccd1 vccd1 _17746_/A sky130_fd_sc_hd__or2_1
X_14949_ _15838_/D _15702_/D _15717_/C _15976_/D vssd1 vssd1 vccd1 vccd1 _15169_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17668_ _17915_/A _19439_/A _17665_/Y _17666_/X vssd1 vssd1 vccd1 vccd1 _17669_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_19407_ _19285_/A _19284_/B _19282_/X vssd1 vssd1 vccd1 vccd1 _19422_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_148_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16619_ _17146_/A _17146_/B _17334_/B _18166_/A vssd1 vssd1 vccd1 vccd1 _16622_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_134_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17599_ _19636_/A _17599_/B vssd1 vssd1 vccd1 vccd1 _17599_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19338_ _19340_/A vssd1 vssd1 vccd1 vccd1 _19501_/A sky130_fd_sc_hd__inv_2
XANTENNA__16092__A_N _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20717__A _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19269_ _19406_/A _19268_/C _19268_/A vssd1 vssd1 vccd1 vccd1 _19271_/C sky130_fd_sc_hd__a21o_1
XANTENNA__17729__C _18851_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21300_ _21300_/A _21300_/B vssd1 vssd1 vccd1 vccd1 _21310_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17448__D _17670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14390__A1 _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21231_ _21231_/A _21231_/B vssd1 vssd1 vccd1 vccd1 _21234_/A sky130_fd_sc_hd__xor2_2
Xhold200 hold200/A vssd1 vssd1 vccd1 vccd1 hold200/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold211 hold211/A vssd1 vssd1 vccd1 vccd1 hold211/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout202_A _21817_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold222 hold222/A vssd1 vssd1 vccd1 vccd1 hold222/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold233 hold233/A vssd1 vssd1 vccd1 vccd1 hold233/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 hold318/A vssd1 vssd1 vccd1 vccd1 hold244/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21162_ _21162_/A _21162_/B vssd1 vssd1 vccd1 vccd1 _21163_/B sky130_fd_sc_hd__nand2_1
Xhold255 hold255/A vssd1 vssd1 vccd1 vccd1 hold255/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20463__B2 _18008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10951__A1 _10950_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold266 hold266/A vssd1 vssd1 vccd1 vccd1 hold266/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold277 hold277/A vssd1 vssd1 vccd1 vccd1 hold277/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 hold288/A vssd1 vssd1 vccd1 vccd1 hold288/X sky130_fd_sc_hd__buf_4
X_20113_ _20114_/A _20114_/B vssd1 vssd1 vccd1 vccd1 _20258_/B sky130_fd_sc_hd__or2_1
Xhold299 hold299/A vssd1 vssd1 vccd1 vccd1 hold299/X sky130_fd_sc_hd__buf_4
XFILLER_0_102_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21093_ _21093_/A _21093_/B vssd1 vssd1 vccd1 vccd1 _21095_/B sky130_fd_sc_hd__or2_2
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15890__A1 _12291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20044_ _19891_/A _19893_/B _19891_/B vssd1 vssd1 vccd1 vccd1 _20049_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__18279__D _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout571_A _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18857__A _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17092__B1 _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21283__A _21283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21995_ _22021_/CLK _21995_/D vssd1 vssd1 vccd1 vccd1 hold170/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__16377__A _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_106 sstream_i[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15281__A _15281_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_117 sstream_i[70] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_128 v1z[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18295__C _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20946_ _20946_/A _20946_/B _20946_/C vssd1 vssd1 vccd1 vccd1 _20946_/X sky130_fd_sc_hd__and3_1
XANTENNA_139 v1z[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16198__A2 _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold247_A hold247/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19688__A _19823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20877_ _20877_/A _20877_/B _20877_/C vssd1 vssd1 vccd1 vccd1 _20880_/B sky130_fd_sc_hd__nor3_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12300_ _12511_/A _12402_/A _12858_/C _12991_/D vssd1 vssd1 vccd1 vccd1 _12302_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13280_ _13280_/A _13280_/B _13266_/Y vssd1 vssd1 vccd1 vccd1 _13280_/Y sky130_fd_sc_hd__nor3b_4
XFILLER_0_106_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12231_ _12232_/A _12232_/B vssd1 vssd1 vccd1 vccd1 _12238_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_122_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21429_ hold231/X sstream_i[6] _21489_/S vssd1 vssd1 vccd1 vccd1 _21956_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_121_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15159__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12145__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20454__A1 _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20454__B2 _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ _14698_/A _12269_/D vssd1 vssd1 vccd1 vccd1 _12165_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10942__A1 _10941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11984__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ _10941_/X hold54/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21707_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_130_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16970_ _17141_/A _16968_/C _17013_/C _17141_/B vssd1 vssd1 vccd1 vccd1 _16971_/C
+ sky130_fd_sc_hd__a22o_1
X_12093_ _12093_/A _12093_/B _12093_/C vssd1 vssd1 vccd1 vccd1 _12100_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_21_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15921_ _15921_/A _15921_/B vssd1 vssd1 vccd1 vccd1 _15923_/B sky130_fd_sc_hd__or2_1
X_11044_ _11043_/X hold59/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21652_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_21_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18189__D _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13892__B1 _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17093__D _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18767__A _19535_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11195__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18640_ _18789_/A _18640_/B _18640_/C _18784_/A vssd1 vssd1 vccd1 vccd1 _18784_/B
+ sky130_fd_sc_hd__nand4_1
X_15852_ _16196_/A _16196_/B _16396_/B _16418_/B vssd1 vssd1 vccd1 vccd1 _15972_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__18486__B _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14803_ _14804_/A _14804_/B vssd1 vssd1 vccd1 vccd1 _14925_/B sky130_fd_sc_hd__and2b_1
X_18571_ _18572_/A _18572_/B _18572_/C vssd1 vssd1 vccd1 vccd1 _18571_/Y sky130_fd_sc_hd__nor3_1
X_15783_ _15907_/A _15782_/B _15782_/C vssd1 vssd1 vccd1 vccd1 _15784_/B sky130_fd_sc_hd__o21ai_2
XTAP_3640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12995_ _12995_/A _13128_/B _12995_/C vssd1 vssd1 vccd1 vccd1 _12997_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17522_ _17619_/A _17636_/B _17522_/C _17522_/D vssd1 vssd1 vccd1 vccd1 _17524_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_3673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14734_ _14734_/A _14734_/B vssd1 vssd1 vccd1 vccd1 _14735_/B sky130_fd_sc_hd__and2_2
XTAP_3684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11946_ _11964_/A _11964_/B vssd1 vssd1 vccd1 vccd1 _12027_/A sky130_fd_sc_hd__nor2_1
XTAP_3695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_143_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17453_ _17453_/A _17453_/B _17453_/C vssd1 vssd1 vccd1 vccd1 _17455_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_131_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14665_ _15695_/A _15022_/B _14666_/C _14666_/D vssd1 vssd1 vccd1 vccd1 _14665_/X
+ sky130_fd_sc_hd__and4_1
XTAP_2983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11877_ _12020_/A _12511_/A _12402_/A _12326_/D vssd1 vssd1 vccd1 vccd1 _11878_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16404_ _16404_/A _16404_/B vssd1 vssd1 vccd1 vccd1 _16408_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11224__A _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13616_ _13616_/A _13616_/B vssd1 vssd1 vccd1 vccd1 _13618_/B sky130_fd_sc_hd__xnor2_2
X_17384_ _21792_/Q _17493_/A _20797_/A _21258_/A vssd1 vssd1 vccd1 vccd1 _17386_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10828_ hold206/A hold223/A vssd1 vssd1 vccd1 vccd1 _10828_/Y sky130_fd_sc_hd__nor2_1
X_14596_ _14596_/A _14596_/B vssd1 vssd1 vccd1 vccd1 _14599_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16734__B _16734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19123_ _19123_/A _19123_/B _20247_/D vssd1 vssd1 vccd1 vccd1 _19445_/B sky130_fd_sc_hd__and3_1
XFILLER_0_138_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16335_ _16335_/A _16335_/B vssd1 vssd1 vccd1 vccd1 _16337_/C sky130_fd_sc_hd__xor2_1
X_13547_ _13430_/X _13433_/Y _13669_/B _13546_/X vssd1 vssd1 vccd1 vccd1 _13548_/A
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__18652__D _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19054_ _19054_/A _19054_/B vssd1 vssd1 vccd1 vccd1 _19064_/A sky130_fd_sc_hd__xor2_1
X_16266_ _16391_/A _16414_/A _16266_/C vssd1 vssd1 vccd1 vccd1 _16266_/X sky130_fd_sc_hd__and3_1
XFILLER_0_113_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13478_ _13478_/A _13478_/B _13478_/C vssd1 vssd1 vccd1 vccd1 _13480_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_125_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18005_ _18005_/A _18005_/B vssd1 vssd1 vccd1 vccd1 _18020_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15217_ _15217_/A _16027_/B _15361_/A _15217_/D vssd1 vssd1 vccd1 vccd1 _15361_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_140_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12429_ _12427_/X _12429_/B vssd1 vssd1 vccd1 vccd1 _12430_/B sky130_fd_sc_hd__and2b_1
X_16197_ _16309_/A vssd1 vssd1 vccd1 vccd1 _16199_/D sky130_fd_sc_hd__inv_2
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15148_ _15147_/A _15147_/B _15298_/B _15146_/D vssd1 vssd1 vccd1 vccd1 _15148_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_22_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21087__B _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15079_ _15217_/A _16380_/B _15361_/A _15217_/D vssd1 vssd1 vccd1 vccd1 _15215_/B
+ sky130_fd_sc_hd__nand4_2
X_19956_ _20091_/A _19956_/B _20087_/B vssd1 vssd1 vccd1 vccd1 _19958_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13296__A2_N _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18907_ _19695_/A _20103_/A _18766_/X _18767_/X _19089_/B vssd1 vssd1 vccd1 vccd1
+ _18912_/A sky130_fd_sc_hd__a32o_1
X_19887_ _19923_/A vssd1 vssd1 vccd1 vccd1 _19887_/Y sky130_fd_sc_hd__inv_2
X_18838_ _18687_/A _18534_/Y _18687_/B vssd1 vssd1 vccd1 vccd1 _18838_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__12221__C _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18769_ _19695_/A _18769_/B vssd1 vssd1 vccd1 vccd1 _18770_/B sky130_fd_sc_hd__nand2_1
X_20800_ _21256_/A _21153_/B _20800_/C _20800_/D vssd1 vssd1 vccd1 vccd1 _20931_/B
+ sky130_fd_sc_hd__and4_1
X_21780_ _21809_/CLK _21780_/D vssd1 vssd1 vccd1 vccd1 hold326/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20731_ _20991_/C _21283_/B _21305_/B _20863_/C vssd1 vssd1 vccd1 vccd1 _20735_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout152_A _19092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16925__A _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20662_ _20662_/A _20662_/B vssd1 vssd1 vccd1 vccd1 _20664_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_133_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20593_ _20593_/A _20593_/B vssd1 vssd1 vccd1 vccd1 _20594_/B sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_33_clk_i_A clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout417_A _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19955__B _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16660__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21214_ _21214_/A _21214_/B vssd1 vssd1 vccd1 vccd1 _21216_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_44_1223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21278__A _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20987__A2 _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21145_ _21035_/A _21035_/B _21077_/B vssd1 vssd1 vccd1 vccd1 _21185_/A sky130_fd_sc_hd__o21ai_1
Xfanout510 _21742_/Q vssd1 vssd1 vccd1 vccd1 _16203_/D sky130_fd_sc_hd__buf_4
Xfanout521 _13877_/A vssd1 vssd1 vccd1 vccd1 _14024_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout532 _21737_/Q vssd1 vssd1 vccd1 vccd1 _13864_/B sky130_fd_sc_hd__buf_4
Xfanout543 _21735_/Q vssd1 vssd1 vccd1 vccd1 _15155_/C sky130_fd_sc_hd__clkbuf_8
X_21076_ _20920_/A _20920_/B _20960_/X vssd1 vssd1 vccd1 vccd1 _21077_/C sky130_fd_sc_hd__o21ai_1
XANTENNA__13874__B1 _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20910__A _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout554 _14774_/D vssd1 vssd1 vccd1 vccd1 _13554_/B sky130_fd_sc_hd__clkbuf_8
Xfanout565 _21730_/Q vssd1 vssd1 vccd1 vccd1 _12621_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__17065__B1 _17086_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout576 _21727_/Q vssd1 vssd1 vccd1 vccd1 _12269_/C sky130_fd_sc_hd__buf_4
X_20027_ _20178_/D _20841_/B _20025_/Y _20175_/A vssd1 vssd1 vccd1 vccd1 _20027_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__17604__A2 _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout587 _11549_/A vssd1 vssd1 vccd1 vccd1 _21718_/D sky130_fd_sc_hd__buf_6
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout598 _21723_/Q vssd1 vssd1 vccd1 vccd1 _11122_/A sky130_fd_sc_hd__buf_8
XANTENNA__13626__B1 _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ _11801_/A _11801_/B _11801_/C vssd1 vssd1 vccd1 vccd1 _11800_/Y sky130_fd_sc_hd__nor3_2
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ _12780_/A _12780_/B _13034_/D _14386_/B vssd1 vssd1 vccd1 vccd1 _12780_/X
+ sky130_fd_sc_hd__and4_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21978_ _22005_/CLK _21978_/D vssd1 vssd1 vccd1 vccd1 hold214/A sky130_fd_sc_hd__dfxtp_1
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12785__D _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11731_ _12458_/A _13155_/A _13155_/B _12357_/C vssd1 vssd1 vccd1 vccd1 _11732_/C
+ sky130_fd_sc_hd__a22o_1
X_20929_ _21842_/Q _21264_/B _20930_/C _20930_/D vssd1 vssd1 vccd1 vccd1 _20932_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_90_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16835__A _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14450_ _21725_/D hold57/X _10886_/Y fanout6/X _14449_/Y vssd1 vssd1 vccd1 vccd1
+ _14450_/X sky130_fd_sc_hd__a221o_1
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ _11662_/A _11662_/B vssd1 vssd1 vccd1 vccd1 _11664_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__16554__B _16734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13401_ _13554_/B _13858_/C _13402_/D _13556_/A vssd1 vssd1 vccd1 vccd1 _13404_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18868__A1 _19650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14381_ _14381_/A _14381_/B vssd1 vssd1 vccd1 vccd1 _14431_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_14_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11593_ _11593_/A _11593_/B vssd1 vssd1 vccd1 vccd1 _11610_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16120_ _16120_/A vssd1 vssd1 vccd1 vccd1 _16120_/Y sky130_fd_sc_hd__inv_2
XANTENNA__20563__A1_N _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13332_ _13332_/A _13332_/B _13332_/C vssd1 vssd1 vccd1 vccd1 _13335_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_52_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17540__A1 _21802_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16051_ _16052_/A _16052_/B vssd1 vssd1 vccd1 vccd1 _16226_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_121_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17666__A _17666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13263_ _13411_/B _13263_/B _13263_/C vssd1 vssd1 vccd1 vccd1 _13265_/A sky130_fd_sc_hd__and3_1
XFILLER_0_51_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15002_ _14878_/D _14878_/Y _15000_/Y _15001_/X vssd1 vssd1 vccd1 vccd1 _15004_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_20_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12214_ _12269_/A _12245_/B _12214_/C _12246_/C vssd1 vssd1 vccd1 vccd1 _12217_/A
+ sky130_fd_sc_hd__and4_1
X_13194_ _13193_/B _13193_/C _13193_/A vssd1 vssd1 vccd1 vccd1 _13196_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12145_ _12223_/A _12246_/D vssd1 vssd1 vccd1 vccd1 _12146_/B sky130_fd_sc_hd__nand2_1
X_19810_ _19650_/D _20178_/B _20721_/C _19810_/D vssd1 vssd1 vccd1 vccd1 _19813_/A
+ sky130_fd_sc_hd__and4b_1
XANTENNA__12117__B1 _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16953_ _16954_/B _16954_/A vssd1 vssd1 vccd1 vccd1 _16961_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_21_1020 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12076_ _12076_/A _12076_/B vssd1 vssd1 vccd1 vccd1 _12079_/A sky130_fd_sc_hd__nand2_1
X_19741_ _19595_/X _19608_/A _19608_/B _19597_/B vssd1 vssd1 vccd1 vccd1 _19743_/C
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13418__B _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12668__A1 _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18497__A _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12668__B2 _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15904_ _16034_/A _15904_/B _15904_/C vssd1 vssd1 vccd1 vccd1 _15905_/B sky130_fd_sc_hd__or3_1
X_11027_ mstream_o[101] hold247/X _11027_/S vssd1 vssd1 vccd1 vccd1 _21638_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_95_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19672_ _19671_/B _19671_/C _19660_/Y vssd1 vssd1 vccd1 vccd1 _19672_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_95_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16884_ _17029_/A _17019_/C _17124_/C _17029_/B vssd1 vssd1 vccd1 vccd1 _16884_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11340__A1 _11339_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18623_ _18624_/A _19089_/B _18624_/C _18624_/D vssd1 vssd1 vccd1 vccd1 _18625_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15835_ _15836_/B _15835_/B vssd1 vssd1 vccd1 vccd1 _15837_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_56_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18554_ _18849_/A _18849_/B _19199_/C _19199_/D vssd1 vssd1 vccd1 vccd1 _18709_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15766_ _15892_/A _15892_/B _16286_/B _16173_/B vssd1 vssd1 vccd1 vccd1 _15767_/B
+ sky130_fd_sc_hd__and4_1
XTAP_3470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12978_ _13102_/B _12978_/B vssd1 vssd1 vccd1 vccd1 _12988_/A sky130_fd_sc_hd__or2_1
XTAP_3481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21155__A2 _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17505_ _17504_/C _17741_/B _17618_/A _17503_/Y vssd1 vssd1 vccd1 vccd1 _17505_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_14717_ _14715_/X _14716_/Y _14418_/A _14418_/B vssd1 vssd1 vccd1 vccd1 _14717_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_87_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19009__A2_N _19185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18485_ _20088_/A _19703_/C _18486_/C _18486_/D vssd1 vssd1 vccd1 vccd1 _18487_/A
+ sky130_fd_sc_hd__a22oi_1
X_11929_ _11928_/A _11928_/C _11928_/B vssd1 vssd1 vccd1 vccd1 _11941_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_129_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15697_ _15838_/D _15698_/B _15698_/C _15698_/D vssd1 vssd1 vccd1 vccd1 _15699_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12840__B2 _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17436_ _17434_/X _17436_/B vssd1 vssd1 vccd1 vccd1 _17437_/B sky130_fd_sc_hd__and2b_1
X_14648_ _14649_/A _14649_/B vssd1 vssd1 vccd1 vccd1 _14648_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_131_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20267__A _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_17 _11335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16464__B _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_28 _11343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_39 _11436_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17367_ _17265_/A _17264_/B _17264_/A vssd1 vssd1 vccd1 vccd1 _17369_/B sky130_fd_sc_hd__o21bai_4
XANTENNA__10793__A _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14579_ _14579_/A _14579_/B vssd1 vssd1 vccd1 vccd1 _14580_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_43_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19106_ _19106_/A _19106_/B vssd1 vssd1 vccd1 vccd1 _19115_/A sky130_fd_sc_hd__nand2_1
X_16318_ _16319_/A _16319_/B vssd1 vssd1 vccd1 vccd1 _16318_/X sky130_fd_sc_hd__and2_1
XFILLER_0_125_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17298_ _17190_/Y _17193_/X _17296_/A _17297_/Y vssd1 vssd1 vccd1 vccd1 _17382_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19037_ _19037_/A _19037_/B _19037_/C vssd1 vssd1 vccd1 vccd1 _19037_/X sky130_fd_sc_hd__and3_1
X_16249_ _16098_/A _16098_/B _16099_/Y vssd1 vssd1 vccd1 vccd1 _16250_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_88_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16480__A _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20714__B _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20418__A1 _21842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15808__B _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14712__B _14712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17726__D _19691_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15096__A _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20433__C _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12108__B1 _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19939_ _19939_/A _19939_/B vssd1 vssd1 vccd1 vccd1 _19942_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21394__A2 _15210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21901_ _21942_/CLK _21901_/D vssd1 vssd1 vccd1 vccd1 hold188/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__19015__B _19181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11882__A2 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16270__A1 _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout367_A _15916_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16270__B2 _16380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21832_ _21837_/CLK _21832_/D vssd1 vssd1 vccd1 vccd1 _21832_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA__11095__A0 _11055_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18011__A2 _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21763_ _21963_/CLK _21763_/D vssd1 vssd1 vccd1 vccd1 _21763_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_66_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout534_A _21737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20714_ _20838_/B _20975_/D _21286_/B _21296_/B vssd1 vssd1 vccd1 vccd1 _20843_/A
+ sky130_fd_sc_hd__and4_1
X_21694_ _22080_/CLK _21694_/D vssd1 vssd1 vccd1 vccd1 hold82/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16374__B _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20645_ _20900_/A _20645_/B vssd1 vssd1 vccd1 vccd1 _20645_/X sky130_fd_sc_hd__xor2_2
XFILLER_0_18_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20608__C _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11398__A1 _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20576_ _20441_/B _20442_/Y _20574_/X _20575_/Y vssd1 vssd1 vccd1 vccd1 _20578_/B
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__16325__A2 _16396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11949__D _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12898__A1 _21743_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21822__CLK _21822_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12898__B2 _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21082__A1 _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11570__A1 _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11570__B2 _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21128_ _21238_/B _21130_/B vssd1 vssd1 vccd1 vccd1 _21131_/A sky130_fd_sc_hd__nand2_1
Xfanout340 _14635_/D vssd1 vssd1 vccd1 vccd1 _14155_/D sky130_fd_sc_hd__buf_4
Xfanout351 hold241/A vssd1 vssd1 vccd1 vccd1 _16377_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14060__D _14217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout362 _16273_/A vssd1 vssd1 vccd1 vccd1 _16369_/A sky130_fd_sc_hd__buf_4
Xfanout373 _21775_/Q vssd1 vssd1 vccd1 vccd1 _15933_/C sky130_fd_sc_hd__buf_2
X_13950_ _13800_/C _13799_/Y _13948_/X _13949_/Y vssd1 vssd1 vccd1 vccd1 _13952_/C
+ sky130_fd_sc_hd__o211a_2
X_21059_ _21059_/A _21059_/B vssd1 vssd1 vccd1 vccd1 _21061_/A sky130_fd_sc_hd__or2_1
Xfanout384 _16173_/A vssd1 vssd1 vccd1 vccd1 _15931_/A sky130_fd_sc_hd__buf_4
XANTENNA__18110__A _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21385__A2 _19636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18786__B1 _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout395 _12319_/C vssd1 vssd1 vccd1 vccd1 _13152_/C sky130_fd_sc_hd__buf_4
X_12901_ _12780_/X _12783_/A _13032_/B _12900_/X vssd1 vssd1 vccd1 vccd1 _12901_/X
+ sky130_fd_sc_hd__o211a_1
X_13881_ _13881_/A _13881_/B vssd1 vssd1 vccd1 vccd1 _13883_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_88_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18467__D _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11473__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15620_ _15445_/Y _15448_/Y _15753_/A _15619_/X vssd1 vssd1 vccd1 vccd1 _15753_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__13254__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ _12827_/A _12827_/B _12831_/X vssd1 vssd1 vccd1 vccd1 _12952_/A sky130_fd_sc_hd__o21ba_2
XFILLER_0_97_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11086__A0 _10978_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15551_ _15931_/A _15931_/B _16377_/B _16414_/B vssd1 vssd1 vccd1 vccd1 _15669_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_96_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12763_ _12764_/A _12764_/B vssd1 vssd1 vccd1 vccd1 _12763_/X sky130_fd_sc_hd__and2_1
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14502_ _14502_/A _14502_/B vssd1 vssd1 vccd1 vccd1 _14512_/A sky130_fd_sc_hd__xor2_2
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21190__B _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18270_ _18270_/A _18270_/B vssd1 vssd1 vccd1 vccd1 _18273_/A sky130_fd_sc_hd__xnor2_1
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19750__A2 _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11714_ _11714_/A _11714_/B vssd1 vssd1 vccd1 vccd1 _11716_/B sky130_fd_sc_hd__xnor2_2
X_15482_ _15347_/A _15347_/B _15344_/X vssd1 vssd1 vccd1 vccd1 _15484_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_1008 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12694_ _12583_/C _12582_/Y _12692_/X _12693_/Y vssd1 vssd1 vccd1 vccd1 _12697_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_139_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17221_ _16989_/C _17520_/A _16594_/B _16592_/X vssd1 vssd1 vccd1 vccd1 _17231_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14433_ _14434_/A _14434_/B vssd1 vssd1 vccd1 vccd1 _14433_/X sky130_fd_sc_hd__and2b_1
XANTENNA__13378__A2 _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11645_ _13012_/B _12402_/A vssd1 vssd1 vccd1 vccd1 _11649_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11389__A1 _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17152_ _17149_/X _17150_/Y _17151_/X vssd1 vssd1 vccd1 vccd1 _17152_/Y sky130_fd_sc_hd__a21oi_1
X_14364_ _14365_/A _14365_/C _21744_/Q _14516_/A vssd1 vssd1 vccd1 vccd1 _14367_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13420__C _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11576_ _14698_/A _12619_/A _14621_/D _13155_/D vssd1 vssd1 vccd1 vccd1 _11576_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18710__B1 _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11859__D _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16103_ _16399_/A _16396_/B _16418_/B _16305_/B vssd1 vssd1 vccd1 vccd1 _16107_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_123_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14327__A1 _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13315_ _13316_/A _13455_/B _13315_/C vssd1 vssd1 vccd1 vccd1 _13451_/A sky130_fd_sc_hd__or3_2
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17083_ _17078_/A _17078_/C _17078_/B vssd1 vssd1 vccd1 vccd1 _17083_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_4_clk_i _21806_/CLK vssd1 vssd1 vccd1 vccd1 _22021_/CLK sky130_fd_sc_hd__clkbuf_16
X_14295_ _14295_/A _14295_/B _14295_/C vssd1 vssd1 vccd1 vccd1 _14296_/B sky130_fd_sc_hd__and3_2
XANTENNA__14813__A _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16034_ _16034_/A _16034_/B _16150_/A vssd1 vssd1 vccd1 vccd1 _16035_/B sky130_fd_sc_hd__or3_1
X_13246_ _13250_/C _13245_/C _13245_/B vssd1 vssd1 vccd1 vccd1 _13247_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_1120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13177_ _13177_/A _13177_/B vssd1 vssd1 vccd1 vccd1 _13179_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11875__C _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__A1 _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12128_ _12127_/B _12128_/B vssd1 vssd1 vccd1 vccd1 _12130_/B sky130_fd_sc_hd__and2b_1
X_17985_ _17985_/A _18121_/B vssd1 vssd1 vccd1 vccd1 _17987_/A sky130_fd_sc_hd__or2_1
XANTENNA__20550__A _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15644__A _15645_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16936_ _16937_/A _16937_/B vssd1 vssd1 vccd1 vccd1 _16936_/Y sky130_fd_sc_hd__nand2b_1
X_12059_ _12109_/C _12269_/C vssd1 vssd1 vccd1 vccd1 _12104_/A sky130_fd_sc_hd__nand2_1
X_19724_ _19722_/X _19723_/Y _19291_/A _19291_/B vssd1 vssd1 vccd1 vccd1 _19847_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11313__B2 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16867_ _17144_/A _16968_/C _17013_/C _17129_/B vssd1 vssd1 vccd1 vccd1 _16867_/X
+ sky130_fd_sc_hd__a22o_1
X_19655_ _19497_/A _19496_/A _19496_/B _19492_/B _19492_/A vssd1 vssd1 vccd1 vccd1
+ _19656_/B sky130_fd_sc_hd__o32ai_4
XANTENNA__11864__A2 _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11383__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15818_ _15816_/B _15816_/C _15816_/A vssd1 vssd1 vccd1 vccd1 _15818_/Y sky130_fd_sc_hd__a21oi_2
X_18606_ _18606_/A _18606_/B _18606_/C vssd1 vssd1 vccd1 vccd1 _18608_/C sky130_fd_sc_hd__nand3_1
X_19586_ _19587_/A _19587_/B _20247_/D vssd1 vssd1 vccd1 vccd1 _19586_/X sky130_fd_sc_hd__and3_1
X_16798_ _16797_/B _16797_/C _16797_/A vssd1 vssd1 vccd1 vccd1 _16800_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_87_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11077__A0 _10919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18537_ _18537_/A _18839_/A vssd1 vssd1 vccd1 vccd1 _18537_/Y sky130_fd_sc_hd__xnor2_4
X_15749_ _15749_/A _15749_/B vssd1 vssd1 vccd1 vccd1 _15752_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_603 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18468_ _19535_/A _18624_/A _18466_/Y _18626_/A vssd1 vssd1 vccd1 vccd1 _18470_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_74_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17419_ _17417_/X _17419_/B vssd1 vssd1 vccd1 vccd1 _17420_/B sky130_fd_sc_hd__and2b_1
XANTENNA__13611__B _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18399_ _21791_/Q _19013_/C _19179_/C _18703_/A vssd1 vssd1 vccd1 vccd1 _18420_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_28_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_522 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20430_ _20433_/D vssd1 vssd1 vccd1 vccd1 _20430_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_71_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17505__A1_N _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15515__B1 _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20361_ _20214_/X _20217_/Y _20359_/Y _20360_/X vssd1 vssd1 vccd1 vccd1 _20363_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_130_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout115_A _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22100_ _22105_/CLK _22100_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[36] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20292_ _20292_/A _20292_/B vssd1 vssd1 vccd1 vccd1 _20294_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22031_ _22038_/CLK _22031_/D vssd1 vssd1 vccd1 vccd1 hold311/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11552__A1 _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18849__B _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19009__B2 _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout484_A _21748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11304__A1 _11303_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16369__B _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12897__B _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11068__A0 _10852_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18584__B _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21291__A _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21815_ _21817_/CLK _21815_/D vssd1 vssd1 vccd1 vccd1 _21815_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11607__A2 _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_1209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21746_ _22005_/CLK _21746_/D vssd1 vssd1 vccd1 vccd1 _21746_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_148_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14617__B _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout28_A fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21677_ _21682_/CLK _21677_/D vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_124_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11430_ hold228/A fanout28/X _11429_/X vssd1 vssd1 vccd1 vccd1 _11430_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_74_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20628_ _20628_/A _20628_/B _20627_/C _20627_/D vssd1 vssd1 vccd1 vccd1 _20628_/X
+ sky130_fd_sc_hd__or4bb_2
XFILLER_0_145_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12137__B _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11679__D _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_1085 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11240__A0 _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11361_ hold176/X fanout29/X _11360_/X vssd1 vssd1 vccd1 vccd1 _11361_/X sky130_fd_sc_hd__a21o_1
XANTENNA__11041__B _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20559_ _20559_/A _20559_/B vssd1 vssd1 vccd1 vccd1 _20567_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13100_ _13100_/A _13240_/A vssd1 vssd1 vccd1 vccd1 _13102_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_81_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14080_ _14078_/X _14080_/B vssd1 vssd1 vccd1 vccd1 _14081_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_120_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11292_ _12991_/D _11291_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21774_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_131_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13031_ _13031_/A _13031_/B vssd1 vssd1 vccd1 vccd1 _13067_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11543__A1 _11089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_2_clk_i_A _21822_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17770_ _17770_/A _17891_/A _17770_/C vssd1 vssd1 vccd1 vccd1 _17891_/B sky130_fd_sc_hd__nand3_2
X_14982_ _15218_/A _14982_/B _15075_/B vssd1 vssd1 vccd1 vccd1 _14984_/B sky130_fd_sc_hd__nand3_1
Xfanout170 _21828_/Q vssd1 vssd1 vccd1 vccd1 _19732_/A sky130_fd_sc_hd__buf_4
Xfanout181 _16868_/A vssd1 vssd1 vccd1 vccd1 _17144_/A sky130_fd_sc_hd__buf_4
XFILLER_0_89_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout192 _21823_/Q vssd1 vssd1 vccd1 vccd1 _17557_/B sky130_fd_sc_hd__clkbuf_4
X_16721_ _16721_/A _16721_/B _16721_/C vssd1 vssd1 vccd1 vccd1 _16723_/A sky130_fd_sc_hd__and3_1
X_13933_ _13933_/A _13933_/B _13933_/C vssd1 vssd1 vccd1 vccd1 _13936_/A sky130_fd_sc_hd__nand3_2
XANTENNA__20520__D _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19440_ _19441_/A _19441_/B _19441_/C vssd1 vssd1 vccd1 vccd1 _19440_/X sky130_fd_sc_hd__a21o_1
X_16652_ _16653_/A _16653_/B _16653_/C vssd1 vssd1 vccd1 vccd1 _16652_/X sky130_fd_sc_hd__and3_1
X_13864_ _21738_/Q _13864_/B _14354_/C _14663_/D vssd1 vssd1 vccd1 vccd1 _13867_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_18_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15603_ _15463_/X _15465_/X _15601_/Y _15602_/X vssd1 vssd1 vccd1 vccd1 _15605_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_97_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19371_ _19246_/A _19246_/B _19246_/C _19248_/X vssd1 vssd1 vccd1 vccd1 _19405_/A
+ sky130_fd_sc_hd__a31o_1
X_12815_ _12701_/A _12701_/C _12701_/B vssd1 vssd1 vccd1 vccd1 _12816_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_85_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16583_ _17199_/B _16582_/C _16582_/A vssd1 vssd1 vccd1 vccd1 _16583_/Y sky130_fd_sc_hd__a21oi_2
X_13795_ _13795_/A _13795_/B _13795_/C _13795_/D vssd1 vssd1 vccd1 vccd1 _13795_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_97_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18322_ _18322_/A _18322_/B vssd1 vssd1 vccd1 vccd1 _18324_/B sky130_fd_sc_hd__or2_1
X_15534_ _15534_/A _15714_/B vssd1 vssd1 vccd1 vccd1 _15545_/A sky130_fd_sc_hd__nand2_1
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12746_ _12652_/X _12655_/Y _12744_/Y _12745_/X vssd1 vssd1 vccd1 vccd1 _12837_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_139_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12973__D _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18253_ _18253_/A _18253_/B vssd1 vssd1 vccd1 vccd1 _18263_/A sky130_fd_sc_hd__or2_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15465_ _15323_/X _15325_/Y _15462_/Y _15464_/X vssd1 vssd1 vccd1 vccd1 _15465_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18850__A1_N _18851_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12677_ _12676_/B _12676_/C _12676_/A vssd1 vssd1 vccd1 vccd1 _12679_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_72_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17204_ _17504_/C _17636_/B _17201_/Y _17203_/B vssd1 vssd1 vccd1 vccd1 _17205_/B
+ sky130_fd_sc_hd__a22oi_1
X_14416_ _14416_/A _14416_/B vssd1 vssd1 vccd1 vccd1 _14419_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_127_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18184_ _18183_/B _18183_/C _18183_/A vssd1 vssd1 vccd1 vccd1 _18220_/B sky130_fd_sc_hd__a21oi_2
X_11628_ _12229_/A _12751_/B _12637_/B _12155_/B vssd1 vssd1 vccd1 vccd1 _11630_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15396_ _15541_/A vssd1 vssd1 vccd1 vccd1 _15398_/D sky130_fd_sc_hd__inv_2
XFILLER_0_128_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12047__B _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11231__B1 _11230_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17135_ _17134_/A _17134_/B _17134_/C vssd1 vssd1 vccd1 vccd1 _17135_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_128_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14347_ _14659_/A _14176_/C _15112_/D _15435_/A vssd1 vssd1 vccd1 vccd1 _14347_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11559_ _12094_/A _12877_/B _12751_/B _12094_/B vssd1 vssd1 vccd1 vccd1 _11560_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14543__A _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17557__C _17670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17066_ _17066_/A _17066_/B _17066_/C vssd1 vssd1 vccd1 vccd1 _17091_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14278_ _14277_/B _14277_/C _14277_/A vssd1 vssd1 vccd1 vccd1 _14279_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16017_ _15496_/B _15496_/C _15626_/A _16016_/X _15496_/A vssd1 vssd1 vccd1 vccd1
+ _16021_/B sky130_fd_sc_hd__a2111o_1
X_13229_ _13229_/A vssd1 vssd1 vccd1 vccd1 _13357_/A sky130_fd_sc_hd__inv_2
XANTENNA__17854__A _18851_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11534__A1 _11089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16473__A1 _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17968_ _17969_/A _18243_/A vssd1 vssd1 vccd1 vccd1 _17968_/Y sky130_fd_sc_hd__nor2_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15093__B _15093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19707_ _19706_/B _19903_/B _19706_/A vssd1 vssd1 vccd1 vccd1 _19708_/C sky130_fd_sc_hd__a21o_1
X_16919_ _17141_/A _16917_/C _16968_/C _17141_/B vssd1 vssd1 vccd1 vccd1 _16920_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17899_ _20583_/A _19892_/A _18319_/B _18622_/B vssd1 vssd1 vccd1 vccd1 _17901_/B
+ sky130_fd_sc_hd__nand4_1
X_19638_ hold137/X _19637_/X fanout4/A vssd1 vssd1 vccd1 vccd1 hold138/A sky130_fd_sc_hd__mux2_1
XFILLER_0_79_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13325__C _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14787__A1 _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19569_ _19569_/A _19569_/B vssd1 vssd1 vccd1 vccd1 _19578_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13044__D _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21600_ _21934_/CLK _21600_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[63] sky130_fd_sc_hd__dfrtp_4
XANTENNA__16636__C _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12262__A2 _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16528__A2 _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14539__A1 _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21531_ hold274/X sstream_i[108] _21536_/S vssd1 vssd1 vccd1 vccd1 _22058_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14539__B2 _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18851__C _18851_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21462_ hold182/X sstream_i[39] _21494_/S vssd1 vssd1 vccd1 vccd1 _21989_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19478__A1 _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20455__A _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15154__A2_N _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20413_ _20863_/C _21264_/A _20413_/C _20603_/A vssd1 vssd1 vccd1 vccd1 _20603_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13762__A2 _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21393_ _21420_/S _21393_/B vssd1 vssd1 vccd1 vccd1 _21393_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20344_ _20195_/X _20197_/Y _20341_/Y _20343_/X vssd1 vssd1 vccd1 vccd1 _20344_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_102_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11288__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20275_ _20275_/A _20275_/B vssd1 vssd1 vccd1 vccd1 _20277_/B sky130_fd_sc_hd__or2_1
XANTENNA__11525__A1 _11089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18579__B _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22014_ _22016_/CLK _22014_/D vssd1 vssd1 vccd1 vccd1 hold200/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__21286__A _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20796__B1 _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_2__f_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13711__A1_N _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold277_A hold277/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12420__B _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10930_ _10931_/B vssd1 vssd1 vccd1 vccd1 _10940_/A sky130_fd_sc_hd__inv_2
XANTENNA__13235__C _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10861_ mstream_o[44] _10860_/Y _10992_/S vssd1 vssd1 vccd1 vccd1 _21581_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_79_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ _12600_/A _12600_/B vssd1 vssd1 vccd1 vccd1 _21340_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_112_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ _13580_/A _13580_/B _13580_/C vssd1 vssd1 vccd1 vccd1 _13581_/B sky130_fd_sc_hd__and3_1
XFILLER_0_94_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10792_ sstream_i[114] vssd1 vssd1 vccd1 vccd1 _10792_/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_94_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12531_ _12530_/A _13012_/B _12530_/C _12530_/D vssd1 vssd1 vccd1 vccd1 _12532_/B
+ sky130_fd_sc_hd__a22o_1
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21729_ _22016_/CLK _21729_/D vssd1 vssd1 vccd1 vccd1 _21729_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15250_ _15108_/A _15250_/B vssd1 vssd1 vccd1 vccd1 _15252_/B sky130_fd_sc_hd__nand2b_2
XFILLER_0_152_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12462_ _12359_/A _12359_/C _12359_/B vssd1 vssd1 vccd1 vccd1 _12463_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_124_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11213__A0 _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14201_ _14201_/A _14201_/B _14201_/C vssd1 vssd1 vccd1 vccd1 _14203_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_34_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11413_ _11412_/X _20991_/C _11446_/S vssd1 vssd1 vccd1 vccd1 _21809_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_152_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15181_ _14954_/B _14956_/B _15179_/X _15180_/Y vssd1 vssd1 vccd1 vccd1 _15331_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12393_ _21725_/D hold132/X _11045_/X fanout6/X _12392_/Y vssd1 vssd1 vccd1 vccd1
+ _12393_/X sky130_fd_sc_hd__a221o_1
X_14132_ _14132_/A _14132_/B vssd1 vssd1 vccd1 vccd1 _14171_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_104_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11344_ _15698_/B _11343_/X _11348_/S vssd1 vssd1 vccd1 vccd1 _21787_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_50_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14082__B _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11198__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14063_ _13901_/A _13901_/C _13901_/B vssd1 vssd1 vccd1 vccd1 _14064_/C sky130_fd_sc_hd__a21bo_1
X_18940_ _18940_/A _19084_/A _18940_/C vssd1 vssd1 vccd1 vccd1 _19084_/B sky130_fd_sc_hd__nand3_1
X_11275_ fanout58/X v0z[12] fanout17/X _11274_/X vssd1 vssd1 vccd1 vccd1 _11275_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11516__A1 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20812__B _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13014_ _12444_/B _13152_/C _13152_/D _13864_/B vssd1 vssd1 vccd1 vccd1 _13014_/X
+ sky130_fd_sc_hd__a22o_1
X_18871_ _20032_/D _19487_/B _19053_/B _19199_/C vssd1 vssd1 vccd1 vccd1 _19028_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_24_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16455__A1 _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13707__A _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17822_ _17698_/A _17698_/C _17698_/B vssd1 vssd1 vccd1 vccd1 _17824_/B sky130_fd_sc_hd__o21ba_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
X_14965_ _14967_/A _14967_/B vssd1 vssd1 vccd1 vccd1 _14965_/X sky130_fd_sc_hd__or2_1
X_17753_ _17750_/X _17751_/Y _17651_/X _17654_/Y vssd1 vssd1 vccd1 vccd1 _17753_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__20003__A2 _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13916_ _13916_/A _13916_/B _14073_/B vssd1 vssd1 vccd1 vccd1 _13916_/X sky130_fd_sc_hd__and3_1
X_16704_ _16705_/A _16705_/B _16705_/C vssd1 vssd1 vccd1 vccd1 _16704_/X sky130_fd_sc_hd__and3_1
X_17684_ _17684_/A _17684_/B _17684_/C vssd1 vssd1 vccd1 vccd1 _17684_/Y sky130_fd_sc_hd__nand3_2
X_14896_ _14896_/A _14896_/B vssd1 vssd1 vccd1 vccd1 _14897_/B sky130_fd_sc_hd__xor2_2
Xclkbuf_leaf_22_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21942_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_1014 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16635_ _16634_/B _16634_/C _16634_/A vssd1 vssd1 vccd1 vccd1 _16635_/Y sky130_fd_sc_hd__a21oi_2
X_19423_ _19563_/B _19422_/C _19422_/A vssd1 vssd1 vccd1 vccd1 _19424_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_76_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13847_ _13685_/A _13686_/Y _13845_/Y _13846_/X vssd1 vssd1 vccd1 vccd1 _13847_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_18_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13572__A2_N _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13442__A _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16566_ _16566_/A _16566_/B _16566_/C vssd1 vssd1 vccd1 vccd1 _16651_/A sky130_fd_sc_hd__and3_1
X_19354_ _19354_/A _19354_/B _19504_/B vssd1 vssd1 vccd1 vccd1 _19356_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13778_ _14089_/A _14087_/A _14557_/D _15234_/C vssd1 vssd1 vccd1 vccd1 _13779_/C
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13441__A1 _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13441__B2 _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15517_ _15517_/A _15517_/B vssd1 vssd1 vccd1 vccd1 _15518_/B sky130_fd_sc_hd__xnor2_2
X_18305_ _18305_/A _18305_/B _18292_/Y vssd1 vssd1 vccd1 vccd1 _18305_/Y sky130_fd_sc_hd__nor3b_4
XFILLER_0_57_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_37_clk_i clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21845_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19285_ _19285_/A _19285_/B vssd1 vssd1 vccd1 vccd1 _19296_/A sky130_fd_sc_hd__xnor2_2
X_12729_ _12730_/A _12730_/B vssd1 vssd1 vccd1 vccd1 _12834_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_155_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16497_ _16781_/A _16781_/B vssd1 vssd1 vccd1 vccd1 _16503_/A sky130_fd_sc_hd__or2_1
XANTENNA__12058__A _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18236_ _18095_/B _18095_/Y _18386_/B _18235_/X vssd1 vssd1 vccd1 vccd1 _18389_/A
+ sky130_fd_sc_hd__a211o_2
X_15448_ _15449_/A _15448_/B vssd1 vssd1 vccd1 vccd1 _15448_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11204__A0 _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18167_ _19373_/B _18769_/B _18167_/C _18167_/D vssd1 vssd1 vccd1 vccd1 _18169_/A
+ sky130_fd_sc_hd__nand4_1
X_15379_ _15379_/A _15379_/B vssd1 vssd1 vccd1 vccd1 _15380_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_128_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__18132__A1 _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17118_ _17110_/B _17110_/C _17110_/A vssd1 vssd1 vccd1 vccd1 _17118_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18098_ _18095_/Y _18096_/X _17962_/B _17964_/A vssd1 vssd1 vccd1 vccd1 _18099_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_141_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15439__A_N _21735_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17049_ _17049_/A _17049_/B _17049_/C vssd1 vssd1 vccd1 vccd1 _17117_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_0_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20060_ _20167_/A _20059_/C _20059_/A vssd1 vssd1 vccd1 vccd1 _20060_/X sky130_fd_sc_hd__o21a_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16446__A1 _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17643__B1 _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16446__B2 _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14463__A_N _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout182_A _21825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_136_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20962_ _20790_/B _20830_/Y _20960_/X _20961_/Y vssd1 vssd1 vccd1 vccd1 _20964_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_36_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15551__B _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20893_ _20726_/A _20726_/B _20727_/Y vssd1 vssd1 vccd1 vccd1 _20895_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_36_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout447_A _21759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11443__A0 _11442_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17174__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21514_ hold238/X sstream_i[91] _21528_/S vssd1 vssd1 vccd1 vccd1 _22041_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_35_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15279__A _15279_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16813__D _17086_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21445_ hold297/X sstream_i[22] _21489_/S vssd1 vssd1 vccd1 vccd1 _21972_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19974__A _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20286__A1_N _21839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21376_ _14296_/Y _19169_/Y _21420_/S vssd1 vssd1 vccd1 vccd1 _21376_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_32_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20327_ _20328_/A _20327_/B vssd1 vssd1 vccd1 vccd1 _20327_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_43_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17925__C _19703_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout95_A fanout96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11060_ _11059_/Y hold66/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21659_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_101_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18426__A2 _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20258_ _20258_/A _20258_/B _20258_/C vssd1 vssd1 vccd1 vccd1 _20260_/C sky130_fd_sc_hd__nand3_1
XANTENNA__18102__B _21355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20189_ _20975_/D _20671_/B _19987_/X _19988_/X fanout96/X vssd1 vssd1 vccd1 vccd1
+ _20196_/A sky130_fd_sc_hd__a32oi_4
XANTENNA__16988__A2 _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_clk_i_A clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11692__D _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13120__B1 _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15660__A2 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14750_ _14750_/A _14750_/B vssd1 vssd1 vccd1 vccd1 _14751_/B sky130_fd_sc_hd__xnor2_4
XTAP_3844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11962_ _11969_/B _11960_/X _11954_/Y _11957_/Y vssd1 vssd1 vccd1 vccd1 _11964_/D
+ sky130_fd_sc_hd__o211a_1
XTAP_3855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13701_ _13697_/Y _13699_/X _13583_/X _13586_/Y vssd1 vssd1 vccd1 vccd1 _13702_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_3877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10913_ mstream_o[51] _10912_/X _10992_/S vssd1 vssd1 vccd1 vccd1 _21588_/D sky130_fd_sc_hd__mux2_1
XTAP_3888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14681_ _14521_/A _14521_/C _14521_/B vssd1 vssd1 vccd1 vccd1 _14682_/C sky130_fd_sc_hd__a21bo_1
X_11893_ _11830_/B _11830_/C _11830_/D _11833_/B vssd1 vssd1 vccd1 vccd1 _11893_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16420_ _16420_/A _16420_/B vssd1 vssd1 vccd1 vccd1 _16421_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13632_ _13632_/A _13632_/B _13632_/C vssd1 vssd1 vccd1 vccd1 _13635_/A sky130_fd_sc_hd__nand3_2
X_10844_ _11061_/A _11061_/B _10810_/A vssd1 vssd1 vccd1 vccd1 _11063_/A sky130_fd_sc_hd__o21a_2
XFILLER_0_6_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19868__B _19868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14077__B _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11434__A0 _11433_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18772__B _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16351_ _16368_/B _16351_/B vssd1 vssd1 vccd1 vccd1 _16354_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13563_ _13410_/A _13410_/B _13409_/B vssd1 vssd1 vccd1 vccd1 _13565_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__13974__A2 _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16573__A _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19587__C _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15302_ _15439_/D _15698_/B _15303_/C _15303_/D vssd1 vssd1 vccd1 vccd1 _15306_/A
+ sky130_fd_sc_hd__a22oi_1
X_19070_ _19379_/B _19240_/B _19070_/C _19235_/A vssd1 vssd1 vccd1 vccd1 _19235_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_54_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12514_ _12512_/X _12514_/B vssd1 vssd1 vccd1 vccd1 _12515_/B sky130_fd_sc_hd__and2b_1
X_16282_ _16173_/A _16284_/A _16027_/B vssd1 vssd1 vccd1 vccd1 _16283_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_125_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13494_ _13491_/X _13492_/Y _13343_/C _13342_/Y vssd1 vssd1 vccd1 vccd1 _13496_/D
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__21249__A1 _11550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13187__B1 _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18021_ _18020_/B _18020_/C _18020_/A vssd1 vssd1 vccd1 vccd1 _18021_/Y sky130_fd_sc_hd__a21oi_1
X_15233_ _15373_/B _16177_/B _16286_/B _15373_/A vssd1 vssd1 vccd1 vccd1 _15233_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_41_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12445_ _13017_/A _12771_/C _12897_/D _12444_/B vssd1 vssd1 vccd1 vccd1 _12446_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15164_ _14933_/X _14940_/B _14935_/B vssd1 vssd1 vccd1 vccd1 _15166_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_34_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12376_ _12375_/A _12375_/B _12375_/C _12375_/D vssd1 vssd1 vccd1 vccd1 _12376_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_61_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12325__B _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14115_ _13952_/C _13952_/Y _14113_/X _14114_/X vssd1 vssd1 vccd1 vccd1 _14117_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_50_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17873__B1 _20146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11327_ fanout58/X v0z[25] fanout18/X _11326_/X vssd1 vssd1 vccd1 vccd1 _11327_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15095_ _15373_/B _15368_/D _15234_/C _15373_/A vssd1 vssd1 vccd1 vccd1 _15098_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19972_ _19972_/A _20394_/B _19972_/C _21258_/B vssd1 vssd1 vccd1 vccd1 _20110_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__20542__B _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12044__C _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14046_ _14045_/B _14045_/C _14045_/A vssd1 vssd1 vccd1 vccd1 _14046_/Y sky130_fd_sc_hd__o21ai_1
X_18923_ _18758_/B _18758_/Y _19007_/A _18922_/Y vssd1 vssd1 vccd1 vccd1 _19007_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11258_ _11502_/A1 t1x[8] v2z[8] _11501_/B2 _11257_/X vssd1 vssd1 vccd1 vccd1 _11258_/X
+ sky130_fd_sc_hd__a221o_2
XANTENNA__16428__A1 _16173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14540__B _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13437__A _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18854_ _18854_/A _19017_/B _18855_/B vssd1 vssd1 vccd1 vccd1 _19024_/A sky130_fd_sc_hd__or3_1
X_11189_ _14384_/C _11188_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21746_/D sky130_fd_sc_hd__mux2_1
X_17805_ _17805_/A _17805_/B _17805_/C vssd1 vssd1 vccd1 vccd1 _17805_/Y sky130_fd_sc_hd__nand3_2
X_15997_ _15999_/C vssd1 vssd1 vccd1 vccd1 _16134_/B sky130_fd_sc_hd__inv_2
X_18785_ _19439_/A _19414_/C _18646_/X _18647_/X _19874_/B vssd1 vssd1 vccd1 vccd1
+ _18790_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_59_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14948_ _15838_/D _15717_/C _15976_/D _15702_/D vssd1 vssd1 vccd1 vccd1 _14951_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21373__B _21373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17736_ _17736_/A _17736_/B vssd1 vssd1 vccd1 vccd1 _17750_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14879_ _14699_/Y _14701_/X _14877_/X _14878_/Y vssd1 vssd1 vccd1 vccd1 _14881_/B
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__10796__A _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17667_ _17665_/Y _17666_/X _17915_/A _19439_/A vssd1 vssd1 vccd1 vccd1 _17669_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13172__A _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19406_ _19406_/A _19406_/B vssd1 vssd1 vccd1 vccd1 _19406_/X sky130_fd_sc_hd__and2_1
X_16618_ _16617_/B _16617_/C _16617_/A vssd1 vssd1 vccd1 vccd1 _16631_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_147_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17598_ hold215/X fanout3/X _17596_/Y _17597_/X vssd1 vssd1 vccd1 vccd1 _21890_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__11425__A0 _11424_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16549_ _16549_/A _17197_/A vssd1 vssd1 vccd1 vccd1 _16550_/B sky130_fd_sc_hd__nor2_1
X_19337_ _19185_/D _20178_/B _20721_/C _19337_/D vssd1 vssd1 vccd1 vccd1 _19340_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_45_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_1082 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19268_ _19268_/A _19406_/A _19268_/C vssd1 vssd1 vccd1 vccd1 _19406_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_61_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17729__D _19060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18219_ _18220_/A _18220_/B _18220_/C _18220_/D vssd1 vssd1 vccd1 vccd1 _18219_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_143_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19199_ _20178_/D _20032_/D _19199_/C _19199_/D vssd1 vssd1 vccd1 vccd1 _19348_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_115_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21230_ _21230_/A _21230_/B vssd1 vssd1 vccd1 vccd1 _21231_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_13_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14390__A2 _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold201 hold201/A vssd1 vssd1 vccd1 vccd1 hold201/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__19853__A1 _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20733__A _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold212 hold212/A vssd1 vssd1 vccd1 vccd1 hold212/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold223 hold223/A vssd1 vssd1 vccd1 vccd1 hold223/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold234 hold234/A vssd1 vssd1 vccd1 vccd1 hold234/X sky130_fd_sc_hd__dlygate4sd3_1
X_21161_ _21161_/A _21161_/B _21159_/Y vssd1 vssd1 vccd1 vccd1 _21162_/B sky130_fd_sc_hd__or3b_1
Xhold245 hold245/A vssd1 vssd1 vccd1 vccd1 hold245/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold256 hold256/A vssd1 vssd1 vccd1 vccd1 hold256/X sky130_fd_sc_hd__buf_4
Xhold267 hold267/A vssd1 vssd1 vccd1 vccd1 hold267/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 hold278/A vssd1 vssd1 vccd1 vccd1 hold278/X sky130_fd_sc_hd__dlygate4sd3_1
X_20112_ _20112_/A _20112_/B vssd1 vssd1 vccd1 vccd1 _20114_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold289 hold289/A vssd1 vssd1 vccd1 vccd1 hold289/X sky130_fd_sc_hd__dlygate4sd3_1
X_21092_ _21091_/A _21091_/B _21091_/C vssd1 vssd1 vccd1 vccd1 _21093_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_1_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15890__A2 _15888_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20043_ _20043_/A _20043_/B vssd1 vssd1 vccd1 vccd1 _20051_/A sky130_fd_sc_hd__nand2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17092__A1 _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18857__B _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17092__B2 _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout564_A _12621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21283__B _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11259__A3 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21994_ _22021_/CLK _21994_/D vssd1 vssd1 vccd1 vccd1 hold123/A sky130_fd_sc_hd__dfxtp_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_107 sstream_i[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_118 sstream_i[71] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20945_ _21054_/B vssd1 vssd1 vccd1 vccd1 _20946_/C sky130_fd_sc_hd__inv_2
XANTENNA_129 v1z[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18295__D _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19969__A _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14178__A _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18873__A _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20876_ _20873_/X _20874_/Y _20741_/Y _20743_/Y vssd1 vssd1 vccd1 vccd1 _20877_/C
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__19688__B _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_438 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11416__A0 _11415_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout10_A _11547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12426__A _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12230_ _12222_/A _12224_/B _12222_/B vssd1 vssd1 vccd1 vccd1 _12232_/B sky130_fd_sc_hd__o21ba_1
X_21428_ hold255/X sstream_i[5] _21442_/S vssd1 vssd1 vccd1 vccd1 _21955_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12145__B _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15159__D _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12161_ _12160_/A _12159_/Y _12115_/X _12133_/Y vssd1 vssd1 vccd1 vccd1 _12168_/A
+ sky130_fd_sc_hd__o211a_1
X_21359_ _21412_/A _13369_/B fanout40/X vssd1 vssd1 vccd1 vccd1 _21359_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_130_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11112_ _10934_/Y hold168/X _11112_/S vssd1 vssd1 vccd1 vccd1 _21706_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_124_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11984__B _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15456__B _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12092_ _12091_/B _12091_/C _12091_/A vssd1 vssd1 vccd1 vccd1 _12093_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__11476__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15920_ _15920_/A _16050_/B vssd1 vssd1 vccd1 vccd1 _15923_/A sky130_fd_sc_hd__or2_1
XFILLER_0_120_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11043_ _11045_/A _11043_/B vssd1 vssd1 vccd1 vccd1 _11043_/X sky130_fd_sc_hd__and2_2
XANTENNA__13892__A1 _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13892__B2 _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18767__B _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15851_ _15854_/D vssd1 vssd1 vccd1 vccd1 _15851_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17671__B _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16568__A _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14802_ _14802_/A _14802_/B vssd1 vssd1 vccd1 vccd1 _14804_/B sky130_fd_sc_hd__xnor2_1
X_15782_ _15907_/A _15782_/B _15782_/C vssd1 vssd1 vccd1 vccd1 _15784_/A sky130_fd_sc_hd__or3_1
X_18570_ _18565_/Y _18567_/X _18413_/Y _18416_/X vssd1 vssd1 vccd1 vccd1 _18572_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_3630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21167__B1 _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ _13860_/A _13573_/D _13128_/A _12993_/D vssd1 vssd1 vccd1 vccd1 _12995_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_3641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14733_ _14732_/B _14732_/C _14732_/A vssd1 vssd1 vccd1 vccd1 _14734_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_86_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17521_ _17520_/A _17300_/C _17520_/D _17520_/B vssd1 vssd1 vccd1 vccd1 _17522_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11945_ _11870_/Y _11942_/X _11941_/X _11927_/X vssd1 vssd1 vccd1 vccd1 _11964_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_2940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18583__A1 _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18583__B2 _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17452_ _17340_/A _17340_/C _17340_/B vssd1 vssd1 vccd1 vccd1 _17453_/C sky130_fd_sc_hd__a21bo_1
X_14664_ _15695_/A _15022_/B _14666_/C _14666_/D vssd1 vssd1 vccd1 vccd1 _14664_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_2973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11876_ _11879_/A vssd1 vssd1 vccd1 vccd1 _11876_/Y sky130_fd_sc_hd__inv_2
XTAP_2995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16403_ _16403_/A _16403_/B vssd1 vssd1 vccd1 vccd1 _16411_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_39_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11407__A0 _11406_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13615_ _13616_/B _13616_/A vssd1 vssd1 vccd1 vccd1 _13758_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_27_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11224__B _11555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17383_ _17294_/A _17294_/B _17292_/X vssd1 vssd1 vccd1 vccd1 _17409_/A sky130_fd_sc_hd__a21oi_1
X_10827_ hold212/A hold194/A vssd1 vssd1 vccd1 vccd1 _11045_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_131_1267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14595_ _14595_/A _14595_/B vssd1 vssd1 vccd1 vccd1 _14596_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_89_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16334_ _16335_/B _16335_/A vssd1 vssd1 vccd1 vccd1 _16388_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__16734__C _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19122_ _19123_/A _19123_/B vssd1 vssd1 vccd1 vccd1 _19126_/A sky130_fd_sc_hd__or2_1
X_13546_ _13545_/A _13545_/B _13669_/A _13545_/D vssd1 vssd1 vccd1 vccd1 _13546_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_54_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_471 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14535__B _15892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16897__A1 _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19053_ _20178_/D _19053_/B vssd1 vssd1 vccd1 vccd1 _19054_/B sky130_fd_sc_hd__nand2_1
X_16265_ _16414_/A _16266_/C _16414_/B _16391_/A vssd1 vssd1 vccd1 vccd1 _16265_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13477_ _13327_/A _13327_/C _13327_/B vssd1 vssd1 vccd1 vccd1 _13478_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__11878__C _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15216_ _15217_/A _16027_/B _15361_/A _15217_/D vssd1 vssd1 vccd1 vccd1 _15218_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18004_ _18004_/A _18004_/B vssd1 vssd1 vccd1 vccd1 _18005_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_51_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12428_ _12642_/A _14698_/A _13155_/D _12637_/A vssd1 vssd1 vccd1 vccd1 _12429_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16196_ _16196_/A _16196_/B _16399_/B _16409_/B vssd1 vssd1 vccd1 vccd1 _16309_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_23_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15147_ _15147_/A _15147_/B _15298_/B _15146_/D vssd1 vssd1 vccd1 vccd1 _15147_/X
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12359_ _12359_/A _12359_/B _12359_/C vssd1 vssd1 vccd1 vccd1 _12362_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_11_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15078_ _15217_/A _16380_/B _15361_/A _15217_/D vssd1 vssd1 vccd1 vccd1 _15080_/B
+ sky130_fd_sc_hd__a22o_1
X_19955_ _20088_/A _20247_/C _20087_/A _19955_/D vssd1 vssd1 vccd1 vccd1 _20087_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__21087__C _21853_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18958__A _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11386__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14029_ _14025_/X _14027_/Y _13863_/X _13866_/X vssd1 vssd1 vccd1 vccd1 _14030_/B
+ sky130_fd_sc_hd__a211o_1
X_18906_ _18906_/A _18906_/B vssd1 vssd1 vccd1 vccd1 _18914_/A sky130_fd_sc_hd__nand2_1
X_19886_ _19743_/X _19763_/X _19883_/Y _19885_/X vssd1 vssd1 vccd1 vccd1 _19923_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__21384__A _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18837_ _18837_/A _18837_/B vssd1 vssd1 vccd1 vccd1 _18841_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_101_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12221__D _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18768_ _19089_/B _18767_/X _18766_/X vssd1 vssd1 vccd1 vccd1 _18770_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_26_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17719_ _17962_/A _17719_/B vssd1 vssd1 vccd1 vccd1 _17819_/A sky130_fd_sc_hd__and2_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11646__B1 _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18699_ _18701_/A _18853_/B vssd1 vssd1 vccd1 vccd1 _18702_/A sky130_fd_sc_hd__or2_1
XFILLER_0_26_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20730_ _20730_/A _20730_/B vssd1 vssd1 vccd1 vccd1 _20738_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_133_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16925__B _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20661_ _20662_/B _20662_/A vssd1 vssd1 vccd1 vccd1 _20661_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_92_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18433__A2_N _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20592_ _20590_/D _21293_/B _21261_/B _20462_/D vssd1 vssd1 vccd1 vccd1 _20593_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_45_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__21330__B1 _11089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout312_A _21793_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16660__B _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21213_ _21286_/A _21311_/B vssd1 vssd1 vccd1 vccd1 _21214_/B sky130_fd_sc_hd__nand2_1
XANTENNA__21278__B _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21144_ hold146/X _21143_/X fanout1/X vssd1 vssd1 vccd1 vccd1 hold147/A sky130_fd_sc_hd__mux2_1
Xfanout500 _15717_/B vssd1 vssd1 vccd1 vccd1 _16196_/A sky130_fd_sc_hd__buf_4
XFILLER_0_6_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11296__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout511 _14195_/A vssd1 vssd1 vccd1 vccd1 _13155_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__20592__A2_N _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout522 _14813_/A vssd1 vssd1 vccd1 vccd1 _15838_/D sky130_fd_sc_hd__buf_4
Xfanout533 _21737_/Q vssd1 vssd1 vccd1 vccd1 _15435_/A sky130_fd_sc_hd__buf_4
X_21075_ _21075_/A _21228_/B _21075_/C vssd1 vssd1 vccd1 vccd1 _21077_/B sky130_fd_sc_hd__or3_1
XANTENNA__13874__A1 _21741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout544 _12750_/A vssd1 vssd1 vccd1 vccd1 _12637_/B sky130_fd_sc_hd__buf_4
XANTENNA__13874__B2 _13875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout555 _14774_/D vssd1 vssd1 vccd1 vccd1 _14306_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__20910__B _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17065__A1 _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout566 _12403_/B vssd1 vssd1 vccd1 vccd1 _12246_/C sky130_fd_sc_hd__buf_4
X_20026_ _20462_/D _20026_/B _20838_/C _20838_/D vssd1 vssd1 vccd1 vccd1 _20175_/A
+ sky130_fd_sc_hd__and4_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17065__B2 _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout577 _13525_/A vssd1 vssd1 vccd1 vccd1 _12302_/A sky130_fd_sc_hd__buf_4
Xfanout588 _11549_/A vssd1 vssd1 vccd1 vccd1 _11502_/A1 sky130_fd_sc_hd__buf_4
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout599 _16363_/A vssd1 vssd1 vccd1 vccd1 _21725_/D sky130_fd_sc_hd__buf_6
XANTENNA__13626__A1 _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13626__B2 _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout58_A fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21977_ _22021_/CLK _21977_/D vssd1 vssd1 vccd1 vccd1 hold220/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_95_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11730_ _12784_/A _13157_/A vssd1 vssd1 vccd1 vccd1 _11732_/B sky130_fd_sc_hd__and2_1
XFILLER_0_138_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20928_ _21048_/A vssd1 vssd1 vccd1 vccd1 _20930_/D sky130_fd_sc_hd__inv_2
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16835__B _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ _11659_/X _11661_/B vssd1 vssd1 vccd1 vccd1 _11662_/B sky130_fd_sc_hd__and2b_1
X_20859_ _21296_/A _21283_/B _21305_/B _20991_/C vssd1 vssd1 vccd1 vccd1 _20863_/D
+ sky130_fd_sc_hd__a22o_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13400_ _13400_/A _13400_/B vssd1 vssd1 vccd1 vccd1 _13501_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16554__C _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14380_ _14379_/B _14379_/C _14379_/A vssd1 vssd1 vccd1 vccd1 _14381_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18868__A2 _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11592_ _11593_/A _11593_/B vssd1 vssd1 vccd1 vccd1 _11592_/X sky130_fd_sc_hd__and2_1
XFILLER_0_91_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13331_ _13330_/A _13330_/B _13330_/C vssd1 vssd1 vccd1 vccd1 _13332_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_64_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19638__S fanout4/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_1015 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17540__A2 _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16050_ _16050_/A _16050_/B vssd1 vssd1 vccd1 vccd1 _16052_/B sky130_fd_sc_hd__or2_1
XFILLER_0_107_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13262_ _13121_/A _13121_/C _13121_/B vssd1 vssd1 vccd1 vccd1 _13263_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_121_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15001_ _15375_/A _15001_/B _15001_/C _15001_/D vssd1 vssd1 vccd1 vccd1 _15001_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_0_121_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12213_ _12183_/A _12183_/C _12183_/B vssd1 vssd1 vccd1 vccd1 _12219_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_122_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13193_ _13193_/A _13193_/B _13193_/C vssd1 vssd1 vccd1 vccd1 _13196_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_32_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12144_ _12144_/A _12144_/B vssd1 vssd1 vccd1 vccd1 _12146_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_130_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12117__A1 _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12117__B2 _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19740_ _19740_/A _19740_/B _19740_/C _19740_/D vssd1 vssd1 vccd1 vccd1 _19743_/B
+ sky130_fd_sc_hd__nand4_1
X_16952_ _16952_/A _16952_/B vssd1 vssd1 vccd1 vccd1 _16954_/B sky130_fd_sc_hd__or2_1
X_12075_ _12076_/A _12075_/B _12075_/C vssd1 vssd1 vccd1 vccd1 _12076_/B sky130_fd_sc_hd__nand3_1
XANTENNA__13865__A1 _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13418__C _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12668__A2 _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17056__A1 _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18497__B _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12322__C _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15903_ _16034_/A _15904_/B _15904_/C vssd1 vssd1 vccd1 vccd1 _15905_/A sky130_fd_sc_hd__o21ai_2
X_11026_ mstream_o[100] hold290/X _11027_/S vssd1 vssd1 vccd1 vccd1 _21637_/D sky130_fd_sc_hd__mux2_1
XANTENNA__21408__S _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19671_ _19660_/Y _19671_/B _19671_/C vssd1 vssd1 vccd1 vccd1 _19671_/X sky130_fd_sc_hd__and3b_1
X_16883_ _16989_/C _17145_/B vssd1 vssd1 vccd1 vccd1 _16935_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_155_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16803__B2 _16734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18622_ _19092_/A _18622_/B _18773_/B _19546_/D vssd1 vssd1 vccd1 vccd1 _18624_/D
+ sky130_fd_sc_hd__nand4_4
X_15834_ _15834_/A _15834_/B vssd1 vssd1 vccd1 vccd1 _15836_/B sky130_fd_sc_hd__or2_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18553_ _18849_/A _19199_/C _19199_/D _18849_/B vssd1 vssd1 vccd1 vccd1 _18553_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__11628__B1 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15765_ _15892_/B _16286_/B _16173_/B _15892_/A vssd1 vssd1 vccd1 vccd1 _15767_/A
+ sky130_fd_sc_hd__a22oi_1
XTAP_3460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12977_ _13381_/C _13997_/C _12976_/C _12976_/D vssd1 vssd1 vccd1 vccd1 _12978_/B
+ sky130_fd_sc_hd__a22oi_1
XTAP_3471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17504_ _17618_/A _17503_/Y _17504_/C _17741_/B vssd1 vssd1 vccd1 vccd1 _17618_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_59_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14716_ _14716_/A _16380_/B _14848_/B _14848_/C vssd1 vssd1 vccd1 vccd1 _14716_/Y
+ sky130_fd_sc_hd__nand4_2
X_11928_ _11928_/A _11928_/B _11928_/C vssd1 vssd1 vccd1 vccd1 _11941_/A sky130_fd_sc_hd__nand3_1
X_15696_ _15834_/A vssd1 vssd1 vccd1 vccd1 _15698_/D sky130_fd_sc_hd__inv_2
X_18484_ _18787_/A _19732_/B _18640_/B _19092_/C vssd1 vssd1 vccd1 vccd1 _18486_/D
+ sky130_fd_sc_hd__nand4_1
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12840__A2 _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14647_ _14647_/A _14647_/B vssd1 vssd1 vccd1 vccd1 _14649_/B sky130_fd_sc_hd__nor2_2
X_17435_ _19892_/A _19951_/A _19951_/B _17434_/B vssd1 vssd1 vccd1 vccd1 _17436_/B
+ sky130_fd_sc_hd__a22o_1
X_11859_ _12897_/C _12897_/D _12619_/A _13556_/A vssd1 vssd1 vccd1 vccd1 _11859_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_67_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20267__B _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_18 _11335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15790__A1 _15916_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14578_ _14579_/B _14579_/A vssd1 vssd1 vccd1 vccd1 _14578_/X sky130_fd_sc_hd__and2b_1
XANTENNA_29 _11343_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17366_ _17366_/A _17366_/B vssd1 vssd1 vccd1 vccd1 _17369_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19105_ _19105_/A _19105_/B vssd1 vssd1 vccd1 vccd1 _19139_/A sky130_fd_sc_hd__and2_1
X_16317_ _16206_/A _16321_/A _16205_/B _16202_/B _16202_/A vssd1 vssd1 vccd1 vccd1
+ _16319_/B sky130_fd_sc_hd__o32ai_4
X_13529_ _13975_/B _13682_/C _14155_/C _14155_/D vssd1 vssd1 vccd1 vccd1 _13678_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_83_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17857__A _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17297_ _17297_/A _17297_/B _17297_/C vssd1 vssd1 vccd1 vccd1 _17297_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_3_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16248_ _16248_/A _16248_/B vssd1 vssd1 vccd1 vccd1 _16250_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19036_ _19035_/B _19035_/C _19035_/A vssd1 vssd1 vccd1 vccd1 _19037_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_141_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16480__B _17141_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13553__B1 _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20418__A2 _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16179_ _16287_/A _16180_/B vssd1 vssd1 vccd1 vccd1 _16179_/X sky130_fd_sc_hd__or2_1
XFILLER_0_141_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15808__C _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14712__C _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15096__B _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12108__A1 _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12108__B2 _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21379__A0 _14449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19938_ _19936_/Y _19938_/B vssd1 vssd1 vccd1 vccd1 _19939_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_103_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19869_ _19869_/A _19869_/B vssd1 vssd1 vccd1 vccd1 _19877_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13625__A _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21900_ _21942_/CLK hold98/X vssd1 vssd1 vccd1 vccd1 hold97/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__19992__B1 _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16270__A2 _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21831_ _21837_/CLK _21831_/D vssd1 vssd1 vccd1 vccd1 _21831_/Q sky130_fd_sc_hd__dfxtp_2
XANTENNA_fanout262_A _21803_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21762_ _21963_/CLK _21762_/D vssd1 vssd1 vccd1 vccd1 _21762_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_37_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12292__B1 _11043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20458__A _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20713_ _20838_/B _21286_/B _21296_/B _20975_/D vssd1 vssd1 vccd1 vccd1 _20717_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_77_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14033__A1 _21742_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21693_ _22080_/CLK _21693_/D vssd1 vssd1 vccd1 vccd1 hold173/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14033__B2 _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout527_A _21738_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20644_ _20901_/A _20643_/Y _20902_/A vssd1 vssd1 vccd1 vccd1 _20645_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20575_ _20707_/B _20573_/X _20400_/X _20402_/X vssd1 vssd1 vccd1 vccd1 _20575_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_132_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_614 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12898__A2 _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18598__A _19531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11570__A2 _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21127_ _21238_/A _21125_/Y _21008_/A _21012_/B vssd1 vssd1 vccd1 vccd1 _21130_/B
+ sky130_fd_sc_hd__a211o_1
Xfanout330 _21787_/Q vssd1 vssd1 vccd1 vccd1 _16404_/B sky130_fd_sc_hd__clkbuf_8
Xfanout341 _21783_/Q vssd1 vssd1 vccd1 vccd1 _14635_/D sky130_fd_sc_hd__clkbuf_4
Xfanout352 _16414_/A vssd1 vssd1 vccd1 vccd1 _15112_/D sky130_fd_sc_hd__buf_4
Xfanout363 _21778_/Q vssd1 vssd1 vccd1 vccd1 _16273_/A sky130_fd_sc_hd__buf_4
X_21058_ _21169_/A _21171_/B _21169_/B vssd1 vssd1 vccd1 vccd1 _21059_/B sky130_fd_sc_hd__and3_1
Xfanout374 _21775_/Q vssd1 vssd1 vccd1 vccd1 _16286_/A sky130_fd_sc_hd__clkbuf_8
Xfanout385 _21773_/Q vssd1 vssd1 vccd1 vccd1 _16173_/A sky130_fd_sc_hd__buf_4
XANTENNA__18110__B _21791_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18786__A1 _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12900_ _14195_/A _12899_/B _13032_/A _12899_/D vssd1 vssd1 vccd1 vccd1 _12900_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18786__B2 _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout396 _21770_/Q vssd1 vssd1 vccd1 vccd1 _12319_/C sky130_fd_sc_hd__buf_4
X_20009_ _20009_/A _20154_/A _20009_/C vssd1 vssd1 vccd1 vccd1 _20154_/B sky130_fd_sc_hd__nand3_1
X_13880_ _13878_/X _13880_/B vssd1 vssd1 vccd1 vccd1 _13881_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_9_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12831_ _12947_/A _12820_/Y _12831_/C _12831_/D vssd1 vssd1 vccd1 vccd1 _12831_/X
+ sky130_fd_sc_hd__and4bb_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13254__B _14463_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22065__RESET_B fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15172__D _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15550_ _15553_/D vssd1 vssd1 vccd1 vccd1 _15550_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_55_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ _12762_/A _12762_/B vssd1 vssd1 vccd1 vccd1 _12764_/B sky130_fd_sc_hd__xor2_2
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14501_ _15435_/A _15788_/B vssd1 vssd1 vccd1 vccd1 _14502_/B sky130_fd_sc_hd__nand2_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11713_ _11711_/X _11713_/B vssd1 vssd1 vccd1 vccd1 _11714_/B sky130_fd_sc_hd__and2b_1
X_15481_ _15481_/A _15481_/B vssd1 vssd1 vccd1 vccd1 _15484_/A sky130_fd_sc_hd__and2_1
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ _12692_/A _12692_/B _12692_/C _12692_/D vssd1 vssd1 vccd1 vccd1 _12693_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_139_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14432_ _14268_/A _14268_/C _14268_/B vssd1 vssd1 vccd1 vccd1 _14434_/B sky130_fd_sc_hd__a21bo_2
X_17220_ _17297_/A _17219_/C _17219_/A vssd1 vssd1 vccd1 vccd1 _17256_/B sky130_fd_sc_hd__a21oi_2
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11644_ _11643_/A _11643_/B _11643_/C vssd1 vssd1 vccd1 vccd1 _11650_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17151_ _17148_/X _17149_/X _17150_/Y _17138_/X _17133_/B vssd1 vssd1 vccd1 vccd1
+ _17151_/X sky130_fd_sc_hd__o311a_1
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14363_ _14213_/A _14215_/B _14213_/B vssd1 vssd1 vccd1 vccd1 _14368_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__14516__D _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11575_ _12426_/B _12403_/A vssd1 vssd1 vccd1 vccd1 _11579_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13420__D _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16102_ _16102_/A _16102_/B vssd1 vssd1 vccd1 vccd1 _16110_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18710__A1 _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13314_ _13455_/B _13315_/C vssd1 vssd1 vccd1 vccd1 _13316_/B sky130_fd_sc_hd__nor2_1
XANTENNA__18710__B2 _19493_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14327__A2 _15174_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21199__A _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17082_ _17081_/B _17081_/C _17081_/A vssd1 vssd1 vccd1 vccd1 _17156_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_123_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14294_ _13518_/X _14294_/B _14294_/C _14294_/D vssd1 vssd1 vccd1 vccd1 _14295_/C
+ sky130_fd_sc_hd__nand4b_1
XFILLER_0_12_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14813__B _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16033_ _16034_/A _16034_/B _16150_/A vssd1 vssd1 vccd1 vccd1 _16035_/A sky130_fd_sc_hd__o21ai_2
X_13245_ _13250_/C _13245_/B _13245_/C vssd1 vssd1 vccd1 vccd1 _13400_/A sky130_fd_sc_hd__and3_1
XANTENNA__19892__A _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13176_ _13177_/A _13308_/B _13176_/C vssd1 vssd1 vccd1 vccd1 _13304_/A sky130_fd_sc_hd__or3_1
XFILLER_0_0_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11875__D _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11561__A2 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _12127_/A _12127_/B _12127_/C vssd1 vssd1 vccd1 vccd1 _12128_/B sky130_fd_sc_hd__or3_1
X_17984_ _17982_/A _17982_/B _17982_/C vssd1 vssd1 vccd1 vccd1 _18121_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__20550__B _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19723_ _19723_/A _19723_/B _19723_/C vssd1 vssd1 vccd1 vccd1 _19723_/Y sky130_fd_sc_hd__nand3_1
X_16935_ _16935_/A _16935_/B vssd1 vssd1 vccd1 vccd1 _16937_/B sky130_fd_sc_hd__xor2_2
X_12058_ _12229_/A _12155_/B _12246_/C _12246_/D vssd1 vssd1 vccd1 vccd1 _12058_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_74_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11009_ mstream_o[83] hold69/X _11012_/S vssd1 vssd1 vccd1 vccd1 _21620_/D sky130_fd_sc_hd__mux2_1
X_19654_ _19654_/A _19654_/B vssd1 vssd1 vccd1 vccd1 _19656_/A sky130_fd_sc_hd__xnor2_1
X_16866_ _16866_/A _16866_/B _16866_/C vssd1 vssd1 vccd1 vccd1 _16873_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_88_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18605_ _18606_/A _18606_/B _18606_/C vssd1 vssd1 vccd1 vccd1 _18608_/B sky130_fd_sc_hd__a21o_1
X_15817_ _15817_/A vssd1 vssd1 vccd1 vccd1 _15817_/Y sky130_fd_sc_hd__inv_2
X_19585_ _19585_/A _19585_/B vssd1 vssd1 vccd1 vccd1 _19613_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_137_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16797_ _16797_/A _16797_/B _16797_/C vssd1 vssd1 vccd1 vccd1 _16866_/A sky130_fd_sc_hd__nand3_1
XANTENNA__21381__B _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18536_ _18536_/A _18536_/B vssd1 vssd1 vccd1 vccd1 _18839_/A sky130_fd_sc_hd__nor2_2
X_15748_ _15745_/Y _15746_/X _15614_/Y _15616_/Y vssd1 vssd1 vccd1 vccd1 _15749_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__21533__A0 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18467_ _19092_/A _19092_/B _19089_/B _18773_/B vssd1 vssd1 vccd1 vccd1 _18626_/A
+ sky130_fd_sc_hd__and4_1
X_15679_ _15680_/A _15680_/B vssd1 vssd1 vccd1 vccd1 _15815_/B sky130_fd_sc_hd__nand2_1
XANTENNA_290 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13180__A _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_607 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17418_ _17417_/A _17417_/C _17417_/D _17525_/A vssd1 vssd1 vccd1 vccd1 _17419_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13611__C _14218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18398_ _18398_/A _18398_/B vssd1 vssd1 vccd1 vccd1 _18529_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17349_ _17348_/A _17348_/B _17348_/C vssd1 vssd1 vccd1 vccd1 _17351_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_43_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15515__A1 _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20360_ _20357_/Y _20358_/X _20207_/X _20209_/X vssd1 vssd1 vccd1 vccd1 _20360_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_130_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19019_ _19019_/A _19019_/B vssd1 vssd1 vccd1 vccd1 _19021_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_28_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20291_ _20292_/A _20292_/B vssd1 vssd1 vccd1 vccd1 _20440_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout108_A _19692_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22030_ _22038_/CLK _22030_/D vssd1 vssd1 vccd1 vccd1 hold285/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18849__C _21848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20721__A_N _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18768__A1 _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12897__C _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout644_A _21329_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21814_ _21816_/CLK _21814_/D vssd1 vssd1 vccd1 vccd1 hold332/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21524__A0 hold247/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21745_ _22005_/CLK _21745_/D vssd1 vssd1 vccd1 vccd1 _21745_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_93_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21676_ _21682_/CLK _21676_/D vssd1 vssd1 vccd1 vccd1 hold71/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_1176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20627_ _20628_/A _20628_/B _20627_/C _20627_/D vssd1 vssd1 vccd1 vccd1 _20627_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_970 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16832__C _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_1097 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ _21718_/D hold222/X _11126_/B hold209/X vssd1 vssd1 vccd1 vccd1 _11360_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20558_ _20558_/A _20558_/B vssd1 vssd1 vccd1 vccd1 _20569_/A sky130_fd_sc_hd__or2_1
XFILLER_0_62_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11291_ fanout58/X v0z[16] fanout17/X _11290_/X vssd1 vssd1 vccd1 vccd1 _11291_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20489_ _20342_/X _20344_/X _20487_/Y _20488_/X vssd1 vssd1 vccd1 vccd1 _20491_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_120_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13030_ _13029_/B _13029_/C _13029_/A vssd1 vssd1 vccd1 vccd1 _13031_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_131_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14981_ _21766_/Q _21755_/Q _14981_/C _15075_/A vssd1 vssd1 vccd1 vccd1 _15075_/B
+ sky130_fd_sc_hd__nand4_2
Xfanout160 _21829_/Q vssd1 vssd1 vccd1 vccd1 _16743_/B sky130_fd_sc_hd__clkbuf_4
Xfanout171 _16870_/A vssd1 vssd1 vccd1 vccd1 _17096_/A sky130_fd_sc_hd__buf_4
Xfanout182 _21825_/Q vssd1 vssd1 vccd1 vccd1 _16868_/A sky130_fd_sc_hd__clkbuf_2
X_16720_ _16686_/X _16687_/Y _16718_/A _16718_/Y vssd1 vssd1 vccd1 vccd1 _16721_/C
+ sky130_fd_sc_hd__o211ai_2
X_13932_ _13931_/A _13931_/B _13931_/C vssd1 vssd1 vccd1 vccd1 _13933_/C sky130_fd_sc_hd__a21o_1
Xfanout193 _21056_/B vssd1 vssd1 vccd1 vccd1 _20247_/D sky130_fd_sc_hd__buf_4
XFILLER_0_135_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17431__A1 _17417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13863_ _14027_/A _13864_/B _14354_/C _14663_/D vssd1 vssd1 vccd1 vccd1 _13863_/X
+ sky130_fd_sc_hd__and4_1
X_16651_ _16651_/A _16651_/B vssd1 vssd1 vccd1 vccd1 _16653_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_88_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15602_ _15599_/Y _15600_/X _15458_/Y _15460_/Y vssd1 vssd1 vccd1 vccd1 _15602_/X
+ sky130_fd_sc_hd__o211a_1
X_12814_ _12813_/B _12813_/C _12813_/A vssd1 vssd1 vccd1 vccd1 _12816_/B sky130_fd_sc_hd__o21ai_1
X_19370_ _19370_/A _19370_/B vssd1 vssd1 vccd1 vccd1 _19461_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13794_ _13795_/A _13795_/B _13795_/C _13795_/D vssd1 vssd1 vccd1 vccd1 _13794_/Y
+ sky130_fd_sc_hd__nor4_2
X_16582_ _16582_/A _17199_/B _16582_/C vssd1 vssd1 vccd1 vccd1 _17178_/A sky130_fd_sc_hd__and3_1
XFILLER_0_9_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18321_ _18321_/A _18321_/B vssd1 vssd1 vccd1 vccd1 _18324_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_139_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15533_ _15717_/B _15913_/B _15533_/C _15714_/A vssd1 vssd1 vccd1 vccd1 _15714_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_29_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ _12744_/B _12744_/C _12744_/A vssd1 vssd1 vccd1 vccd1 _12745_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_85_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15464_ _15464_/A _15464_/B _15464_/C vssd1 vssd1 vccd1 vccd1 _15464_/X sky130_fd_sc_hd__and3_1
X_18252_ _18143_/A _18142_/B _18142_/A vssd1 vssd1 vccd1 vccd1 _18265_/A sky130_fd_sc_hd__o21ba_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21716__SET_B _21329_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12676_ _12676_/A _12676_/B _12676_/C vssd1 vssd1 vccd1 vccd1 _12679_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_127_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14415_ _14848_/A _14557_/D vssd1 vssd1 vccd1 vccd1 _14416_/B sky130_fd_sc_hd__nand2_2
XANTENNA__21421__S _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17203_ _17281_/A _17203_/B _17504_/C _17636_/B vssd1 vssd1 vccd1 vccd1 _17281_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_5_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11627_ _11625_/X _11626_/Y _12223_/A _12751_/B vssd1 vssd1 vccd1 vccd1 _11787_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_155_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15395_ _15791_/A _16371_/A _16399_/A _16424_/A vssd1 vssd1 vccd1 vccd1 _15541_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_108_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18183_ _18183_/A _18183_/B _18183_/C vssd1 vssd1 vccd1 vccd1 _18183_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__15838__A_N _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14346_ _14201_/A _14201_/B _14201_/C _14203_/X vssd1 vssd1 vccd1 vccd1 _14379_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11231__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17200__A _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17134_ _17134_/A _17134_/B _17134_/C vssd1 vssd1 vccd1 vccd1 _17134_/Y sky130_fd_sc_hd__nand3_1
X_11558_ _12223_/A _12637_/B vssd1 vssd1 vccd1 vccd1 _11815_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14543__B _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17557__D _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17065_ _17146_/A _17063_/C _17086_/C _17146_/B vssd1 vssd1 vccd1 vccd1 _17066_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_69_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14277_ _14277_/A _14277_/B _14277_/C vssd1 vssd1 vccd1 vccd1 _14279_/A sky130_fd_sc_hd__and3_1
XFILLER_0_100_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19239__A2 _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11489_ _11498_/A1 t1y[13] t0x[13] _11501_/B2 vssd1 vssd1 vccd1 vccd1 _11489_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_110_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16016_ _16016_/A _16016_/B _16016_/C vssd1 vssd1 vccd1 vccd1 _16016_/X sky130_fd_sc_hd__or3_1
X_13228_ _12969_/A _12969_/B _13112_/B _13110_/Y vssd1 vssd1 vccd1 vccd1 _13229_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17854__B _17854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15655__A _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ _13020_/A _13020_/C _13020_/B vssd1 vssd1 vccd1 vccd1 _13160_/C sky130_fd_sc_hd__a21bo_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16473__A2 _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17967_ _17967_/A _17967_/B vssd1 vssd1 vccd1 vccd1 _18243_/A sky130_fd_sc_hd__xnor2_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19706_ _19706_/A _19706_/B _19903_/B vssd1 vssd1 vccd1 vccd1 _19708_/B sky130_fd_sc_hd__nand3_1
X_16918_ _17145_/A _17013_/C vssd1 vssd1 vccd1 vccd1 _16920_/B sky130_fd_sc_hd__and2_1
XANTENNA__11298__A1 _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17898_ _19823_/A _18624_/A vssd1 vssd1 vccd1 vccd1 _17901_/A sky130_fd_sc_hd__and2_1
X_19637_ hold169/A fanout7/X _21384_/B _11550_/A _19636_/Y vssd1 vssd1 vccd1 vccd1
+ _19637_/X sky130_fd_sc_hd__a221o_1
X_16849_ _16849_/A _16849_/B _16849_/C vssd1 vssd1 vccd1 vccd1 _16850_/B sky130_fd_sc_hd__or3_1
XANTENNA__13325__D _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16917__C _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12247__B1 _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19568_ _20103_/A _19906_/C vssd1 vssd1 vccd1 vccd1 _19569_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_149_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18519_ _18516_/X _18517_/Y _18368_/C _18367_/Y vssd1 vssd1 vccd1 vccd1 _18521_/D
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__16636__D _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19499_ _19499_/A _19499_/B vssd1 vssd1 vccd1 vccd1 _19501_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21530_ hold288/X sstream_i[107] _21536_/S vssd1 vssd1 vccd1 vccd1 _22057_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_91_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11470__A1 _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13747__B1 _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18851__D _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21461_ hold204/X sstream_i[38] _21481_/S vssd1 vssd1 vccd1 vccd1 _21988_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19478__A2 _19476_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout225_A _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20455__B _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_640 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20412_ _20863_/C _21264_/A _20413_/C _20603_/A vssd1 vssd1 vccd1 vccd1 _20414_/A
+ sky130_fd_sc_hd__a22o_1
X_21392_ _21390_/B _21391_/X _21390_/Y vssd1 vssd1 vccd1 vccd1 _21938_/D sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20343_ _20343_/A _20343_/B _20343_/C vssd1 vssd1 vccd1 vccd1 _20343_/X sky130_fd_sc_hd__and3_1
XFILLER_0_141_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_583 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20274_ _20274_/A _20421_/B vssd1 vssd1 vccd1 vccd1 _20277_/A sky130_fd_sc_hd__or2_1
XANTENNA_fanout594_A _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22013_ _22013_/CLK _22013_/D vssd1 vssd1 vccd1 vccd1 hold202/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_41_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18579__C _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20796__A1 _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20796__B2 _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15284__B _15284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14475__A1 _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14475__B2 _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11289__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17780__A _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12420__C _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13235__D _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17930__D _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_3_clk_i _21822_/CLK vssd1 vssd1 vccd1 vccd1 _22020_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_151_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10860_ _10866_/B _10860_/B vssd1 vssd1 vccd1 vccd1 _10860_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_6_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout40_A _21390_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ _11122_/A vssd1 vssd1 vccd1 vccd1 _10791_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_112_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12530_ _12530_/A _13012_/B _12530_/C _12530_/D vssd1 vssd1 vccd1 vccd1 _12532_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__15188__C1 _15050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11461__A1 _17666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21728_ _21974_/CLK _21728_/D vssd1 vssd1 vccd1 vccd1 _21728_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16924__B1 _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20646__A _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12461_ _12460_/B _12460_/C _12460_/A vssd1 vssd1 vccd1 vccd1 _12463_/B sky130_fd_sc_hd__a21o_1
X_21659_ _21934_/CLK _21659_/D vssd1 vssd1 vccd1 vccd1 hold66/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_clkbuf_leaf_24_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14200_ _14040_/A _14040_/C _14040_/B vssd1 vssd1 vccd1 vccd1 _14201_/C sky130_fd_sc_hd__a21bo_1
X_11412_ hold246/A fanout28/X _11411_/X vssd1 vssd1 vccd1 vccd1 _11412_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_151_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15180_ _15179_/B _15179_/C _15179_/A vssd1 vssd1 vccd1 vccd1 _15180_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__14950__A2 _15174_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12392_ fanout9/X _12392_/B vssd1 vssd1 vccd1 vccd1 _12392_/Y sky130_fd_sc_hd__nor2_1
X_14131_ _14131_/A _14131_/B vssd1 vssd1 vccd1 vccd1 _14173_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11479__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11343_ _21407_/S v0z[29] fanout20/X _11342_/X vssd1 vssd1 vccd1 vccd1 _11343_/X
+ sky130_fd_sc_hd__a31o_2
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_1272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14062_ _14062_/A _14062_/B _14062_/C vssd1 vssd1 vccd1 vccd1 _14064_/B sky130_fd_sc_hd__nand3_1
X_11274_ _11493_/A1 t1x[12] v2z[12] _11501_/B2 _11273_/X vssd1 vssd1 vccd1 vccd1 _11274_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_39_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13013_ _13013_/A _13864_/B _13152_/D vssd1 vssd1 vccd1 vccd1 _13013_/X sky130_fd_sc_hd__and3_1
XANTENNA__20812__C _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18870_ _20032_/D _19223_/B _19199_/C _19487_/B vssd1 vssd1 vccd1 vccd1 _18873_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16455__A2 _17063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17821_ _17821_/A _17821_/B vssd1 vssd1 vccd1 vccd1 _17824_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13707__B _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
X_17752_ _17651_/X _17654_/Y _17750_/X _17751_/Y vssd1 vssd1 vccd1 vccd1 _17852_/A
+ sky130_fd_sc_hd__a211o_2
X_14964_ _14964_/A _14964_/B vssd1 vssd1 vccd1 vccd1 _14967_/B sky130_fd_sc_hd__or2_1
X_16703_ _16703_/A _16703_/B vssd1 vssd1 vccd1 vccd1 _16705_/C sky130_fd_sc_hd__xor2_2
X_13915_ _14859_/A _14391_/B _13915_/C _14073_/A vssd1 vssd1 vccd1 vccd1 _14073_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_89_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17683_ _17684_/A _17684_/B _17684_/C vssd1 vssd1 vccd1 vccd1 _17683_/X sky130_fd_sc_hd__and3_1
X_14895_ _14896_/A _14896_/B vssd1 vssd1 vccd1 vccd1 _14895_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14819__A _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19422_ _19422_/A _19563_/B _19422_/C vssd1 vssd1 vccd1 vccd1 _19424_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_134_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16634_ _16634_/A _16634_/B _16634_/C vssd1 vssd1 vccd1 vccd1 _16634_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_57_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13846_ _13846_/A _13846_/B _13846_/C vssd1 vssd1 vccd1 vccd1 _13846_/X sky130_fd_sc_hd__and3_1
XFILLER_0_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13442__B _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19353_ _20032_/D _20193_/D _19353_/C _19504_/A vssd1 vssd1 vccd1 vccd1 _19504_/B
+ sky130_fd_sc_hd__nand4_2
X_13777_ _14087_/A _14557_/D _15234_/C _14089_/A vssd1 vssd1 vccd1 vccd1 _13779_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16565_ _16586_/B _16563_/C _16563_/A vssd1 vssd1 vccd1 vccd1 _16566_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_130_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13441__A2 _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10989_ mstream_o[63] _10988_/Y _11005_/S vssd1 vssd1 vccd1 vccd1 _21600_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18304_ _18304_/A _18304_/B _18304_/C vssd1 vssd1 vccd1 vccd1 _18305_/B sky130_fd_sc_hd__and3_1
X_15516_ _15763_/B _15516_/B vssd1 vssd1 vccd1 vccd1 _15517_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11452__A1 _17557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19284_ _19282_/X _19284_/B vssd1 vssd1 vccd1 vccd1 _19285_/B sky130_fd_sc_hd__and2b_1
X_12728_ _12728_/A _12728_/B vssd1 vssd1 vccd1 vccd1 _12730_/B sky130_fd_sc_hd__or2_2
X_16496_ _17739_/C _17387_/A vssd1 vssd1 vccd1 vccd1 _16781_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_128_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12058__B _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18235_ _18386_/A _18234_/C _18234_/A vssd1 vssd1 vccd1 vccd1 _18235_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_127_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15447_ _15449_/B vssd1 vssd1 vccd1 vccd1 _15448_/B sky130_fd_sc_hd__inv_2
X_12659_ _14024_/B _12899_/B vssd1 vssd1 vccd1 vccd1 _12663_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18166_ _18166_/A _19230_/A _18929_/B _18616_/D vssd1 vssd1 vccd1 vccd1 _18167_/D
+ sky130_fd_sc_hd__nand4_2
X_15378_ _15379_/A _15379_/B vssd1 vssd1 vccd1 vccd1 _15378_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_111_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11389__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17117_ _17117_/A _17117_/B _17117_/C vssd1 vssd1 vccd1 vccd1 _17117_/Y sky130_fd_sc_hd__nand3_1
X_14329_ _14329_/A _14329_/B _14474_/B vssd1 vssd1 vccd1 vccd1 _14331_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_40_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18097_ _17962_/B _17964_/A _18095_/Y _18096_/X vssd1 vssd1 vccd1 vccd1 _18241_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_29_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21387__A _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17048_ _17002_/Y _17009_/X _17040_/X _17114_/A vssd1 vssd1 vccd1 vccd1 _17049_/C
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_141_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17643__A1 _19823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16446__A2 _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17643__B2 _18030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18999_ _18999_/A _19160_/B _18999_/C vssd1 vssd1 vccd1 vccd1 _19000_/B sky130_fd_sc_hd__and3_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18696__A _19185_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15832__B _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20961_ _20960_/B _20960_/C _20960_/A vssd1 vssd1 vccd1 vccd1 _20961_/Y sky130_fd_sc_hd__o21ai_2
XANTENNA__14729__A _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout175_A _21827_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20892_ _20892_/A _20892_/B vssd1 vssd1 vccd1 vccd1 _20895_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13968__B1 _10867_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout342_A _16418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12249__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21513_ hold272/X sstream_i[90] _21528_/S vssd1 vssd1 vccd1 vccd1 _22040_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_119_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout607_A _21718_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21444_ hold302/X sstream_i[21] _21489_/S vssd1 vssd1 vccd1 vccd1 _21971_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_32_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19974__B _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21375_ hold191/X _21381_/B _21373_/Y _21374_/X vssd1 vssd1 vccd1 vccd1 _21932_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18296__A1_N _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20326_ _20328_/B vssd1 vssd1 vccd1 vccd1 _20327_/B sky130_fd_sc_hd__inv_2
XFILLER_0_141_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17925__D _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19990__A _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20257_ _20258_/A _20258_/B _20258_/C vssd1 vssd1 vccd1 vccd1 _20260_/B sky130_fd_sc_hd__a21o_1
X_20188_ _20188_/A _20188_/B vssd1 vssd1 vccd1 vccd1 _20198_/A sky130_fd_sc_hd__or2_1
XANTENNA__12459__B1 _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13120__A1 _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13120__B2 _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11961_ _11954_/Y _11957_/Y _11969_/B _11960_/X vssd1 vssd1 vccd1 vccd1 _11969_/C
+ sky130_fd_sc_hd__a211oi_2
XTAP_3834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_19 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10912_ _10917_/B _10912_/B vssd1 vssd1 vccd1 vccd1 _10912_/X sky130_fd_sc_hd__and2b_2
X_13700_ _13583_/X _13586_/Y _13697_/Y _13699_/X vssd1 vssd1 vccd1 vccd1 _13819_/A
+ sky130_fd_sc_hd__a211oi_2
XTAP_3878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14680_ _14679_/B _14679_/C _14679_/A vssd1 vssd1 vccd1 vccd1 _14682_/B sky130_fd_sc_hd__a21o_1
X_11892_ _11872_/Y _11873_/X _11899_/B _11892_/D vssd1 vssd1 vccd1 vccd1 _11892_/X
+ sky130_fd_sc_hd__and4bb_2
XFILLER_0_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13631_ _13630_/A _13630_/B _13630_/C vssd1 vssd1 vccd1 vccd1 _13632_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_79_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10843_ _10843_/A _10843_/B _10843_/C vssd1 vssd1 vccd1 vccd1 _11061_/B sky130_fd_sc_hd__and3_2
XFILLER_0_6_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16350_ _16349_/A _16349_/B _16349_/C vssd1 vssd1 vccd1 vccd1 _16351_/B sky130_fd_sc_hd__o21ai_1
X_13562_ _13562_/A _13714_/B vssd1 vssd1 vccd1 vccd1 _13565_/A sky130_fd_sc_hd__or2_1
XANTENNA__11434__A1 _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19230__A _19230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16573__B _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15301_ _15437_/A vssd1 vssd1 vccd1 vccd1 _15303_/D sky130_fd_sc_hd__inv_2
XFILLER_0_82_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11985__A2 _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12513_ _12512_/A _12858_/C _12991_/D _12214_/C vssd1 vssd1 vccd1 vccd1 _12514_/B
+ sky130_fd_sc_hd__a22o_1
X_16281_ _16176_/A _16178_/B _16176_/B vssd1 vssd1 vccd1 vccd1 _16383_/S sky130_fd_sc_hd__o21ba_1
XFILLER_0_136_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13493_ _13343_/C _13342_/Y _13491_/X _13492_/Y vssd1 vssd1 vccd1 vccd1 _13496_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13187__A1 _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18020_ _18020_/A _18020_/B _18020_/C vssd1 vssd1 vccd1 vccd1 _18020_/X sky130_fd_sc_hd__and3_1
XFILLER_0_30_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15232_ _15232_/A _15407_/B vssd1 vssd1 vccd1 vccd1 _15242_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_136_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13187__B2 _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12444_ _13017_/A _12444_/B _12771_/C _12897_/D vssd1 vssd1 vccd1 vccd1 _12444_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11198__A0 _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15163_ _15163_/A _15163_/B vssd1 vssd1 vccd1 vccd1 _15166_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_50_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12375_ _12375_/A _12375_/B _12375_/C _12375_/D vssd1 vssd1 vccd1 vccd1 _12375_/X
+ sky130_fd_sc_hd__or4_4
X_14114_ _14113_/A _14113_/B _14111_/Y _14112_/X vssd1 vssd1 vccd1 vccd1 _14114_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_105_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17873__A1 _18008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11326_ _11544_/A1 t1x[25] v2z[25] _11543_/B2 _11325_/X vssd1 vssd1 vccd1 vccd1 _11326_/X
+ sky130_fd_sc_hd__a221o_2
X_15094_ _15094_/A _15094_/B vssd1 vssd1 vccd1 vccd1 _15101_/A sky130_fd_sc_hd__xor2_1
X_19971_ _20394_/B _19972_/C _21258_/B _19972_/A vssd1 vssd1 vccd1 vccd1 _19974_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17873__B2 _18010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14045_ _14045_/A _14045_/B _14045_/C vssd1 vssd1 vccd1 vccd1 _14174_/B sky130_fd_sc_hd__or3_1
X_18922_ _19049_/B _18920_/Y _18780_/X _18817_/A vssd1 vssd1 vccd1 vccd1 _18922_/Y
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__12044__D _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20542__C _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11257_ _11325_/A1 t2y[8] t0y[8] _11498_/A1 vssd1 vssd1 vccd1 vccd1 _11257_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_24_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16428__A2 _16284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13437__B _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18853_ _18853_/A _18853_/B vssd1 vssd1 vccd1 vccd1 _18855_/B sky130_fd_sc_hd__nor2_1
X_11188_ hold166/X fanout22/X _11187_/X vssd1 vssd1 vccd1 vccd1 _11188_/X sky130_fd_sc_hd__a21o_1
X_17804_ _17805_/A _17805_/B _17805_/C vssd1 vssd1 vccd1 vccd1 _17804_/X sky130_fd_sc_hd__and3_1
XFILLER_0_59_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18784_ _18784_/A _18784_/B vssd1 vssd1 vccd1 vccd1 _18793_/A sky130_fd_sc_hd__nand2_1
X_15996_ _15996_/A _16134_/A _15996_/C vssd1 vssd1 vccd1 vccd1 _15999_/C sky130_fd_sc_hd__and3_1
XFILLER_0_89_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17735_ _17736_/A _17736_/B vssd1 vssd1 vccd1 vccd1 _17847_/B sky130_fd_sc_hd__or2_1
X_14947_ _15838_/D _15788_/B _14810_/X _14811_/X _15653_/C vssd1 vssd1 vccd1 vccd1
+ _14952_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_89_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17666_ _17666_/A _19587_/B _17915_/D _17924_/B vssd1 vssd1 vccd1 vccd1 _17666_/X
+ sky130_fd_sc_hd__and4_1
X_14878_ _21769_/Q _16266_/C _14878_/C _14878_/D vssd1 vssd1 vccd1 vccd1 _14878_/Y
+ sky130_fd_sc_hd__nand4_4
XFILLER_0_106_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19405_ _19405_/A _19405_/B vssd1 vssd1 vccd1 vccd1 _19457_/A sky130_fd_sc_hd__xor2_2
XANTENNA__18963__B _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13172__B _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16617_ _16617_/A _16617_/B _16617_/C vssd1 vssd1 vccd1 vccd1 _16631_/A sky130_fd_sc_hd__nand3_2
X_13829_ _13985_/A _16406_/B vssd1 vssd1 vccd1 vccd1 _13831_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17597_ hold60/X fanout7/X _17595_/Y _11550_/A _11553_/Y vssd1 vssd1 vccd1 vccd1
+ _17597_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_15_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20976__A1_N _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11425__A1 _21040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19336_ _19336_/A _19336_/B vssd1 vssd1 vccd1 vccd1 _19341_/A sky130_fd_sc_hd__xnor2_2
X_16548_ _16548_/A _16548_/B vssd1 vssd1 vccd1 vccd1 _17197_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_57_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16364__A1 _10984_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19267_ _19266_/A _19266_/B _19266_/C vssd1 vssd1 vccd1 vccd1 _19268_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_143_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16479_ _17041_/A _16899_/B _17019_/C _17123_/C vssd1 vssd1 vccd1 vccd1 _16479_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_116_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16364__B2 _12291_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18218_ _18214_/X _18216_/Y _18077_/B _18077_/Y vssd1 vssd1 vccd1 vccd1 _18220_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_26_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19198_ _20178_/D _19030_/C _19199_/D _20032_/D vssd1 vssd1 vccd1 vccd1 _19201_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11189__A0 _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18149_ _19644_/A _19240_/B _18293_/A _18147_/Y vssd1 vssd1 vccd1 vccd1 _18150_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_142_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold202 hold202/A vssd1 vssd1 vccd1 vccd1 hold202/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19853__A2 _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold213 hold213/A vssd1 vssd1 vccd1 vccd1 hold213/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20733__B _20991_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14127__B1 _10874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold224 hold224/A vssd1 vssd1 vccd1 vccd1 hold224/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 hold235/A vssd1 vssd1 vccd1 vccd1 hold235/X sky130_fd_sc_hd__dlygate4sd3_1
X_21160_ _21161_/A _21161_/B _21159_/Y vssd1 vssd1 vccd1 vccd1 _21162_/A sky130_fd_sc_hd__o21bai_1
Xhold246 hold246/A vssd1 vssd1 vccd1 vccd1 hold246/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold257 hold257/A vssd1 vssd1 vccd1 vccd1 hold257/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 hold268/A vssd1 vssd1 vccd1 vccd1 hold268/X sky130_fd_sc_hd__dlygate4sd3_1
X_20111_ _20112_/A _20112_/B vssd1 vssd1 vccd1 vccd1 _20258_/A sky130_fd_sc_hd__nand2_1
Xhold279 hold279/A vssd1 vssd1 vccd1 vccd1 hold279/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21091_ _21091_/A _21091_/B _21091_/C vssd1 vssd1 vccd1 vccd1 _21093_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_141_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20042_ _19902_/A _19901_/B _19899_/X vssd1 vssd1 vccd1 vccd1 _20053_/A sky130_fd_sc_hd__a21o_1
XANTENNA__20462__A_N _18008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15627__B1 _10946_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16939__A _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17092__A2 _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18857__C _19181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11113__A0 _10941_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21993_ _22020_/CLK _21993_/D vssd1 vssd1 vccd1 vccd1 hold211/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__14459__A _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16667__A1_N _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout557_A _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_108 sstream_i[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20944_ _21171_/A _21256_/B _20944_/C _20944_/D vssd1 vssd1 vccd1 vccd1 _21054_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA_119 v0z[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20923__A1 _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19969__B _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14178__B _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18873__B _21847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20875_ _20741_/Y _20743_/Y _20873_/X _20874_/Y vssd1 vssd1 vccd1 vccd1 _20877_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11416__A1 _17670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20192__A2_N _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20687__B1 _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20924__A _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12426__B _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21427_ hold249/X sstream_i[4] _21442_/S vssd1 vssd1 vccd1 vccd1 _21954_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_60_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_21_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21945_/CLK sky130_fd_sc_hd__clkbuf_16
X_12160_ _12160_/A _12160_/B _12160_/C vssd1 vssd1 vccd1 vccd1 _12160_/X sky130_fd_sc_hd__or3_1
XFILLER_0_102_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21358_ _21420_/S _21358_/B vssd1 vssd1 vccd1 vccd1 _21358_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11111_ _10926_/X hold26/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21705_/D sky130_fd_sc_hd__mux2_1
X_20309_ _20721_/D _20590_/D _21286_/B _21296_/B vssd1 vssd1 vccd1 vccd1 _20460_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_102_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12091_ _12091_/A _12091_/B _12091_/C vssd1 vssd1 vccd1 vccd1 _12141_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_60_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21289_ _21293_/A _21291_/B _21193_/A _21191_/B vssd1 vssd1 vccd1 vccd1 _21290_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11042_ hold212/A hold194/A vssd1 vssd1 vccd1 vccd1 _11043_/B sky130_fd_sc_hd__or2_1
XFILLER_0_21_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13892__A2 _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_36_clk_i clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21853_/CLK sky130_fd_sc_hd__clkbuf_16
X_15850_ _16196_/B _16396_/B _16418_/B _16196_/A vssd1 vssd1 vccd1 vccd1 _15854_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18280__A1 _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18767__C _19087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17671__C _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16568__B _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18173__A1_N _19379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14801_ _14802_/B _14802_/A vssd1 vssd1 vccd1 vccd1 _14925_/A sky130_fd_sc_hd__and2b_1
XANTENNA__11104__A0 _10874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15781_ _15781_/A _15907_/B vssd1 vssd1 vccd1 vccd1 _15782_/C sky130_fd_sc_hd__nor2_1
XTAP_3620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21167__A1 _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12993_ _13860_/A _13573_/D _13128_/A _12993_/D vssd1 vssd1 vccd1 vccd1 _13128_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_3642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17520_ _17520_/A _17520_/B _20774_/A _17520_/D vssd1 vssd1 vccd1 vccd1 _17522_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_19_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_3653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14732_ _14732_/A _14732_/B _14732_/C vssd1 vssd1 vccd1 vccd1 _14734_/A sky130_fd_sc_hd__nand3_1
XTAP_3664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11944_ _11927_/X _11941_/X _11942_/X _11870_/Y vssd1 vssd1 vccd1 vccd1 _11944_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_59_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17451_ _17450_/B _17450_/C _17450_/A vssd1 vssd1 vccd1 vccd1 _17453_/B sky130_fd_sc_hd__a21o_1
XANTENNA__15397__A2 _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14663_ _16084_/A _16203_/D _14817_/C _14663_/D vssd1 vssd1 vccd1 vccd1 _14666_/D
+ sky130_fd_sc_hd__nand4_1
X_11875_ _12020_/A _12326_/D _12511_/A _12402_/A vssd1 vssd1 vccd1 vccd1 _11879_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16402_ _16406_/A _16404_/B _16308_/A _16306_/B vssd1 vssd1 vccd1 vccd1 _16403_/B
+ sky130_fd_sc_hd__a31o_1
XTAP_2996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13614_ _13614_/A _13614_/B vssd1 vssd1 vccd1 vccd1 _13616_/B sky130_fd_sc_hd__or2_1
XFILLER_0_55_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11407__A1 _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10826_ hold206/A hold223/A vssd1 vssd1 vccd1 vccd1 _10830_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17382_ _17382_/A _17382_/B vssd1 vssd1 vccd1 vccd1 _17475_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_39_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14594_ _14595_/A _14595_/B vssd1 vssd1 vccd1 vccd1 _14594_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19121_ _18964_/A _18964_/B _18964_/C vssd1 vssd1 vccd1 vccd1 _19129_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_54_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16333_ _16333_/A _16333_/B vssd1 vssd1 vccd1 vccd1 _16335_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13545_ _13545_/A _13545_/B _13669_/A _13545_/D vssd1 vssd1 vccd1 vccd1 _13669_/B
+ sky130_fd_sc_hd__nor4_2
XANTENNA__16734__D _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19895__A _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14535__C _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19052_ _19221_/C _19051_/X _19050_/X vssd1 vssd1 vccd1 vccd1 _19054_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_152_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16264_ _16032_/B _16150_/B _16032_/A vssd1 vssd1 vccd1 vccd1 _16372_/A sky130_fd_sc_hd__a21boi_4
X_13476_ _13475_/B _13475_/C _13475_/A vssd1 vssd1 vccd1 vccd1 _13478_/B sky130_fd_sc_hd__a21o_1
XANTENNA__16897__A2 _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15579__A_N _15439_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11878__D _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18003_ _18002_/A _18002_/B _18002_/C vssd1 vssd1 vccd1 vccd1 _18004_/B sky130_fd_sc_hd__a21oi_1
X_15215_ _15361_/A _15215_/B vssd1 vssd1 vccd1 vccd1 _15221_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12427_ _12642_/A _12637_/A _13155_/C _13155_/D vssd1 vssd1 vccd1 vccd1 _12427_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16195_ _16196_/B _16399_/B _16409_/B _16196_/A vssd1 vssd1 vccd1 vccd1 _16199_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15146_ _15147_/A _15147_/B _15298_/B _15146_/D vssd1 vssd1 vccd1 vccd1 _15146_/X
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_10_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12358_ _13173_/C _12357_/C _13034_/D _12458_/A vssd1 vssd1 vccd1 vccd1 _12359_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19119__B _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11309_ _11349_/A1 t2y[21] t0y[21] _21723_/D vssd1 vssd1 vccd1 vccd1 _11309_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15077_ _15076_/A _15076_/B _16173_/B vssd1 vssd1 vccd1 vccd1 _15217_/D sky130_fd_sc_hd__o21a_1
X_19954_ _20088_/A _20247_/C _20087_/A _19955_/D vssd1 vssd1 vccd1 vccd1 _19956_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12289_ _12289_/A _12289_/B vssd1 vssd1 vccd1 vccd1 _17173_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__21087__D _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14028_ _13863_/X _13866_/X _14025_/X _14027_/Y vssd1 vssd1 vccd1 vccd1 _14028_/X
+ sky130_fd_sc_hd__o211a_1
X_18905_ _18905_/A _18905_/B vssd1 vssd1 vccd1 vccd1 _18919_/A sky130_fd_sc_hd__xnor2_1
X_19885_ _19885_/A _19885_/B _19885_/C _19885_/D vssd1 vssd1 vccd1 vccd1 _19885_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__11343__B1 _11342_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18836_ _18837_/A _18837_/B vssd1 vssd1 vccd1 vccd1 _18836_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21384__B _21384_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18767_ _19535_/A _18767_/B _19087_/B vssd1 vssd1 vccd1 vccd1 _18767_/X sky130_fd_sc_hd__and3_1
X_15979_ _15979_/A _16101_/B vssd1 vssd1 vccd1 vccd1 _15981_/B sky130_fd_sc_hd__or2_1
X_17718_ _17718_/A _17718_/B _17718_/C vssd1 vssd1 vccd1 vccd1 _17719_/B sky130_fd_sc_hd__or3_1
XFILLER_0_37_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11646__A1 _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19220__B1 _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18698_ _18853_/A _19181_/B _18857_/B _18698_/D vssd1 vssd1 vccd1 vccd1 _18853_/B
+ sky130_fd_sc_hd__and4b_1
XANTENNA__11646__B2 _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17649_ _17650_/A _17650_/B vssd1 vssd1 vccd1 vccd1 _17649_/X sky130_fd_sc_hd__and2_1
XFILLER_0_37_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16925__C _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20660_ _20913_/A _20660_/B vssd1 vssd1 vccd1 vccd1 _20662_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19319_ _19320_/A _19320_/B _19320_/C vssd1 vssd1 vccd1 vccd1 _19319_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21330__A1 _21349_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20591_ _20593_/A vssd1 vssd1 vccd1 vccd1 _20728_/A sky130_fd_sc_hd__inv_2
XFILLER_0_156_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout138_A _18929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_971 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_678 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout305_A _21794_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21212_ _21212_/A _21212_/B vssd1 vssd1 vccd1 vccd1 _21214_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_13_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11582__B1 _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21143_ hold189/A fanout8/X _21415_/B _11550_/A _21142_/Y vssd1 vssd1 vccd1 vccd1
+ _21143_/X sky130_fd_sc_hd__a221o_1
XANTENNA__15276__C _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout501 _16406_/A vssd1 vssd1 vccd1 vccd1 _15717_/B sky130_fd_sc_hd__buf_2
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout512 _21741_/Q vssd1 vssd1 vccd1 vccd1 _14195_/A sky130_fd_sc_hd__clkbuf_8
Xfanout523 _13877_/A vssd1 vssd1 vccd1 vccd1 _14813_/A sky130_fd_sc_hd__buf_4
X_21074_ _21228_/B _21075_/C _21075_/A vssd1 vssd1 vccd1 vccd1 _21077_/A sky130_fd_sc_hd__o21ai_1
Xfanout534 _21737_/Q vssd1 vssd1 vccd1 vccd1 _15579_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__21397__A1 _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13874__A2 _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout545 _21734_/Q vssd1 vssd1 vccd1 vccd1 _12750_/A sky130_fd_sc_hd__clkbuf_8
Xfanout556 _21732_/Q vssd1 vssd1 vccd1 vccd1 _14774_/D sky130_fd_sc_hd__buf_4
XANTENNA__17065__A2 _17063_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20025_ _20462_/D _20838_/C _20838_/D _20026_/B vssd1 vssd1 vccd1 vccd1 _20025_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout567 _12403_/B vssd1 vssd1 vccd1 vccd1 _12511_/A sky130_fd_sc_hd__buf_4
Xfanout578 _13525_/A vssd1 vssd1 vccd1 vccd1 _13983_/B sky130_fd_sc_hd__buf_4
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout589 _11549_/A vssd1 vssd1 vccd1 vccd1 _11493_/A1 sky130_fd_sc_hd__buf_2
XANTENNA__21725__D _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13626__A2 _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13093__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11606__A _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21976_ _22013_/CLK _21976_/D vssd1 vssd1 vccd1 vccd1 hold119/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16025__B1 _10965_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20927_ _21267_/A _21841_/Q _21816_/Q _21278_/B vssd1 vssd1 vccd1 vccd1 _21048_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_90_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16576__A1 _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ _12402_/A _12858_/C _12991_/D _13525_/A vssd1 vssd1 vccd1 vccd1 _11661_/B
+ sky130_fd_sc_hd__a22o_1
X_20858_ _20858_/A _20858_/B vssd1 vssd1 vccd1 vccd1 _20866_/A sky130_fd_sc_hd__nand2_1
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19650__A_N _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12062__A1 _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16554__D _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11591_ _11591_/A _11591_/B vssd1 vssd1 vccd1 vccd1 _11593_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_135_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20789_ _20788_/A _20788_/B _20788_/C vssd1 vssd1 vccd1 vccd1 _20790_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_148_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18868__A3 _19030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13330_ _13330_/A _13330_/B _13330_/C vssd1 vssd1 vccd1 vccd1 _13332_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_135_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15000__A1 _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13261_ _13554_/B _14018_/C _13411_/A _13260_/D vssd1 vssd1 vccd1 vccd1 _13263_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18555__A2_N _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19278__B1 _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14652__A _14652_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17666__C _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15000_ _15375_/A _15370_/B _15001_/C _15001_/D vssd1 vssd1 vccd1 vccd1 _15000_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12212_ _12193_/A _12193_/C _12193_/B vssd1 vssd1 vccd1 vccd1 _12228_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_60_771 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13192_ _13191_/A _13191_/B _13191_/C vssd1 vssd1 vccd1 vccd1 _13193_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_121_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12143_ _12267_/A _12242_/B _12214_/C _12246_/C vssd1 vssd1 vccd1 vccd1 _12144_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_20_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12117__A2 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16951_ _16951_/A _16997_/A vssd1 vssd1 vccd1 vccd1 _16952_/B sky130_fd_sc_hd__nor2_1
X_12074_ _12011_/Y _12067_/X _12065_/Y _12066_/A vssd1 vssd1 vccd1 vccd1 _12075_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA__21388__A1 _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13865__A2 _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13418__D _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15902_ _15902_/A _15902_/B vssd1 vssd1 vccd1 vccd1 _15904_/C sky130_fd_sc_hd__and2_1
X_11025_ mstream_o[99] hold256/X _11027_/S vssd1 vssd1 vccd1 vccd1 hold257/A sky130_fd_sc_hd__mux2_1
XANTENNA__17056__A2 _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12322__D _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19670_ _19669_/B _19669_/C _19669_/A vssd1 vssd1 vccd1 vccd1 _19671_/C sky130_fd_sc_hd__a21o_1
X_16882_ _17029_/A _17029_/B _17019_/C vssd1 vssd1 vccd1 vccd1 _16882_/X sky130_fd_sc_hd__and3_1
X_18621_ _18622_/B _18773_/B _19546_/D _19092_/A vssd1 vssd1 vccd1 vccd1 _18624_/C
+ sky130_fd_sc_hd__a22o_1
X_15833_ _15833_/A _15959_/B vssd1 vssd1 vccd1 vccd1 _15835_/B sky130_fd_sc_hd__or2_1
XANTENNA__16803__A2 _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18552_ _18552_/A _18552_/B vssd1 vssd1 vccd1 vccd1 _18561_/A sky130_fd_sc_hd__or2_1
XANTENNA__11628__A1 _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15764_ _15764_/A _15764_/B vssd1 vssd1 vccd1 vccd1 _15778_/A sky130_fd_sc_hd__nand2_1
XTAP_3450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11628__B2 _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12976_ _13525_/A _13997_/C _12976_/C _12976_/D vssd1 vssd1 vccd1 vccd1 _13102_/B
+ sky130_fd_sc_hd__and4_1
XTAP_3472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17503_ _17619_/B _21056_/A _21169_/A _17621_/C vssd1 vssd1 vccd1 vccd1 _17503_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_3483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14715_ _14716_/A _16380_/B _14848_/B _14848_/C vssd1 vssd1 vccd1 vccd1 _14715_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18483_ _18787_/B _18640_/B _19092_/C _18787_/A vssd1 vssd1 vccd1 vccd1 _18486_/C
+ sky130_fd_sc_hd__a22o_1
X_11927_ _11928_/A _11928_/B _11928_/C vssd1 vssd1 vccd1 vccd1 _11927_/X sky130_fd_sc_hd__and3_1
X_15695_ _15695_/A _15961_/D _16084_/C _16084_/D vssd1 vssd1 vccd1 vccd1 _15834_/A
+ sky130_fd_sc_hd__and4_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17764__B1 _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17434_ _19892_/A _17434_/B _19951_/A _19951_/B vssd1 vssd1 vccd1 vccd1 _17434_/X
+ sky130_fd_sc_hd__and4_1
X_14646_ _14800_/B _14646_/B vssd1 vssd1 vccd1 vccd1 _14649_/A sky130_fd_sc_hd__nand2b_2
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _11857_/A _11857_/C _11857_/B vssd1 vssd1 vccd1 vccd1 _11870_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_28_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19505__A1 _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19505__B2 fanout96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_19 _11335_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10809_ hold219/A hold58/A vssd1 vssd1 vccd1 vccd1 _10810_/B sky130_fd_sc_hd__or2_1
X_17365_ _17365_/A _17365_/B vssd1 vssd1 vccd1 vccd1 _17366_/B sky130_fd_sc_hd__xnor2_4
X_14577_ _14423_/A _14423_/B _14421_/Y vssd1 vssd1 vccd1 vccd1 _14579_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11789_ _11788_/B _11788_/C _11788_/A vssd1 vssd1 vccd1 vccd1 _11791_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_82_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19104_ _19103_/B _19103_/C _19103_/A vssd1 vssd1 vccd1 vccd1 _19105_/B sky130_fd_sc_hd__a21o_1
X_16316_ _16316_/A _16316_/B vssd1 vssd1 vccd1 vccd1 _16319_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13528_ _13975_/B _14155_/C _14155_/D _13682_/C vssd1 vssd1 vccd1 vccd1 _13528_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17857__B _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17296_ _17296_/A vssd1 vssd1 vccd1 vccd1 _17382_/A sky130_fd_sc_hd__inv_2
XFILLER_0_125_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19035_ _19035_/A _19035_/B _19035_/C vssd1 vssd1 vccd1 vccd1 _19037_/B sky130_fd_sc_hd__nand3_2
X_16247_ _16352_/B _16245_/X _16132_/A _16133_/Y vssd1 vssd1 vccd1 vccd1 _16248_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_140_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13459_ _15076_/A _15076_/B _14212_/D _14384_/D vssd1 vssd1 vccd1 vccd1 _13461_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_70_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13553__A1 _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13553__B2 _13554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16178_ _16178_/A _16178_/B vssd1 vssd1 vccd1 vccd1 _16180_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15129_ _15931_/B _16326_/A _16418_/A _15931_/A vssd1 vssd1 vccd1 vccd1 _15129_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_142_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12108__A2 _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19937_ _19937_/A _19937_/B vssd1 vssd1 vccd1 vccd1 _19938_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11316__A0 _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21379__A1 _19322_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16489__A _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18244__B2 _17969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19868_ _20103_/A _19868_/B vssd1 vssd1 vccd1 vccd1 _19869_/B sky130_fd_sc_hd__and2_1
XFILLER_0_128_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19992__A1 _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13625__B _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18819_ _18669_/C _18668_/Y _18817_/X _18818_/X vssd1 vssd1 vccd1 vccd1 _18822_/C
+ sky130_fd_sc_hd__o211a_2
XANTENNA__19992__B2 _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19799_ _19679_/A _19679_/B _19677_/Y vssd1 vssd1 vccd1 vccd1 _19843_/A sky130_fd_sc_hd__o21ba_1
X_21830_ _21837_/CLK _21830_/D vssd1 vssd1 vccd1 vccd1 _21830_/Q sky130_fd_sc_hd__dfxtp_4
X_21761_ _21974_/CLK _21761_/D vssd1 vssd1 vccd1 vccd1 _21761_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__12292__A1 _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16558__A1 _16870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12292__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout255_A _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20712_ _20712_/A _20712_/B _20712_/C vssd1 vssd1 vccd1 vccd1 _20755_/B sky130_fd_sc_hd__or3_2
XFILLER_0_148_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21692_ _22080_/CLK _21692_/D vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__15230__A1 _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14033__A2 _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_1251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20643_ _20643_/A _20643_/B vssd1 vssd1 vccd1 vccd1 _20643_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_117_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout422_A _12771_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20574_ _20400_/X _20402_/X _20707_/B _20573_/X vssd1 vssd1 vccd1 vccd1 _20574_/X
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_2_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18483__A1 _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18483__B2 _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18598__B _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__C _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21126_ _21008_/A _21012_/B _21238_/A _21125_/Y vssd1 vssd1 vccd1 vccd1 _21238_/B
+ sky130_fd_sc_hd__o211ai_2
Xfanout320 _21791_/Q vssd1 vssd1 vccd1 vccd1 _17493_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__11307__B1 _11306_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout331 _16084_/D vssd1 vssd1 vccd1 vccd1 _15954_/D sky130_fd_sc_hd__buf_4
Xfanout342 _16418_/B vssd1 vssd1 vccd1 vccd1 _15976_/D sky130_fd_sc_hd__buf_4
Xfanout353 _16414_/A vssd1 vssd1 vccd1 vccd1 _15911_/C sky130_fd_sc_hd__buf_4
X_21057_ _21169_/A _21171_/B _21169_/B vssd1 vssd1 vccd1 vccd1 _21059_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__12720__A _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout70_A _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout364 _21778_/Q vssd1 vssd1 vccd1 vccd1 _14018_/C sky130_fd_sc_hd__clkbuf_8
XANTENNA__15049__A1 _15046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout375 _14828_/B vssd1 vssd1 vccd1 vccd1 _12991_/D sky130_fd_sc_hd__buf_4
XANTENNA__18110__C _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout386 _15768_/A vssd1 vssd1 vccd1 vccd1 _13012_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__18786__A2 _21040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20008_ _20007_/B _20143_/B _20007_/A vssd1 vssd1 vccd1 vccd1 _20009_/C sky130_fd_sc_hd__o21ai_1
Xfanout397 _14993_/A vssd1 vssd1 vccd1 vccd1 _14384_/A sky130_fd_sc_hd__buf_4
X_12830_ hold227/X _12829_/X fanout4/A vssd1 vssd1 vccd1 vccd1 _21859_/D sky130_fd_sc_hd__mux2_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13254__C _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20649__A _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ _12762_/A _12762_/B vssd1 vssd1 vccd1 vccd1 _12761_/X sky130_fd_sc_hd__and2_1
XFILLER_0_9_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21959_ _21963_/CLK _21959_/D vssd1 vssd1 vccd1 vccd1 hold314/A sky130_fd_sc_hd__dfxtp_1
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14500_ _13858_/C _14499_/X _14498_/X vssd1 vssd1 vccd1 vccd1 _14502_/A sky130_fd_sc_hd__a21bo_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _12443_/A _12897_/C _12897_/D _12642_/A vssd1 vssd1 vccd1 vccd1 _11713_/B
+ sky130_fd_sc_hd__a22o_1
X_15480_ _15477_/Y _15478_/X _15338_/B _15340_/A vssd1 vssd1 vccd1 vccd1 _15481_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_1086 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ _12692_/A _12692_/B _12692_/C _12692_/D vssd1 vssd1 vccd1 vccd1 _12692_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_37_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14431_ _14431_/A _14431_/B vssd1 vssd1 vccd1 vccd1 _14434_/A sky130_fd_sc_hd__xnor2_4
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _11643_/A _11643_/B _11643_/C vssd1 vssd1 vccd1 vccd1 _11650_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17150_ _17150_/A _17150_/B vssd1 vssd1 vccd1 vccd1 _17150_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_52_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14362_ _14362_/A _14362_/B vssd1 vssd1 vccd1 vccd1 _14370_/A sky130_fd_sc_hd__nand2_1
X_11574_ _11821_/A _11821_/B vssd1 vssd1 vccd1 vccd1 _11610_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16101_ _16101_/A _16101_/B vssd1 vssd1 vccd1 vccd1 _16112_/A sky130_fd_sc_hd__or2_1
XANTENNA__18710__A2 _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13313_ _15217_/A _13034_/D _13310_/Y _13455_/A vssd1 vssd1 vccd1 vccd1 _13315_/C
+ sky130_fd_sc_hd__o2bb2a_1
X_14293_ _14293_/A _14294_/B _14294_/C vssd1 vssd1 vccd1 vccd1 _14295_/B sky130_fd_sc_hd__nand3_1
X_17081_ _17081_/A _17081_/B _17081_/C vssd1 vssd1 vccd1 vccd1 _17156_/A sky130_fd_sc_hd__or3_1
XFILLER_0_134_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16032_ _16032_/A _16032_/B vssd1 vssd1 vccd1 vccd1 _16150_/A sky130_fd_sc_hd__and2_1
XFILLER_0_122_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13244_ _13244_/A _13244_/B vssd1 vssd1 vccd1 vccd1 _13245_/C sky130_fd_sc_hd__or2_1
XANTENNA__19892__B _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18789__A _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13175_ _13308_/B _13176_/C vssd1 vssd1 vccd1 vccd1 _13177_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_27_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21419__S _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ _12076_/B _12084_/X _12124_/A _12123_/Y vssd1 vssd1 vccd1 vccd1 _12127_/C
+ sky130_fd_sc_hd__a211oi_1
X_17983_ _18127_/C vssd1 vssd1 vccd1 vccd1 _17985_/A sky130_fd_sc_hd__inv_2
XANTENNA__13838__A2 _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19722_ _19723_/A _20247_/D _19723_/B _19723_/C vssd1 vssd1 vccd1 vccd1 _19722_/X
+ sky130_fd_sc_hd__a22o_1
X_16934_ _16926_/A _16928_/B _16926_/B vssd1 vssd1 vccd1 vccd1 _16937_/A sky130_fd_sc_hd__o21ba_1
X_12057_ _12057_/A _12057_/B vssd1 vssd1 vccd1 vccd1 _12063_/A sky130_fd_sc_hd__xor2_1
X_11008_ mstream_o[82] hold70/X _11012_/S vssd1 vssd1 vccd1 vccd1 _21619_/D sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_19_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19653_ _19653_/A _19653_/B vssd1 vssd1 vccd1 vccd1 _19654_/B sky130_fd_sc_hd__nor2_1
X_16865_ _16797_/A _16797_/C _16797_/B vssd1 vssd1 vccd1 vccd1 _16866_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_74_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18604_ _18606_/A _18606_/B _18606_/C vssd1 vssd1 vccd1 vccd1 _18604_/Y sky130_fd_sc_hd__a21oi_2
X_15816_ _15816_/A _15816_/B _15816_/C vssd1 vssd1 vccd1 vccd1 _15817_/A sky130_fd_sc_hd__and3_2
X_19584_ _19583_/B _19583_/C _19583_/A vssd1 vssd1 vccd1 vccd1 _19585_/B sky130_fd_sc_hd__a21oi_1
X_16796_ _17141_/A _17223_/A _16860_/C _17141_/B vssd1 vssd1 vccd1 vccd1 _16797_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_99_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18535_ _18687_/A _18534_/C _18534_/A vssd1 vssd1 vccd1 vccd1 _18536_/B sky130_fd_sc_hd__a21oi_1
X_15747_ _15614_/Y _15616_/Y _15745_/Y _15746_/X vssd1 vssd1 vccd1 vccd1 _15749_/A
+ sky130_fd_sc_hd__o211ai_4
XTAP_3280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12959_ _12831_/X _12949_/X _12956_/X _12958_/Y _12951_/B vssd1 vssd1 vccd1 vccd1
+ _12959_/X sky130_fd_sc_hd__a221o_1
XANTENNA__14557__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14776__A2_N _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13461__A _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18466_ _19092_/B _19089_/B _18773_/B _18319_/B vssd1 vssd1 vccd1 vccd1 _18466_/Y
+ sky130_fd_sc_hd__a22oi_1
X_15678_ _15678_/A _15678_/B vssd1 vssd1 vccd1 vccd1 _15680_/B sky130_fd_sc_hd__xnor2_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_280 hold283/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_291 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13180__B _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17417_ _17417_/A _17525_/A _17417_/C _17417_/D vssd1 vssd1 vccd1 vccd1 _17417_/X
+ sky130_fd_sc_hd__and4_1
X_14629_ _14629_/A _14629_/B vssd1 vssd1 vccd1 vccd1 _14630_/B sky130_fd_sc_hd__and2_1
X_18397_ _17841_/Y _18394_/Y _18396_/Y vssd1 vssd1 vccd1 vccd1 _18537_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__13611__D _14873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13774__A1 _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17348_ _17348_/A _17348_/B _17348_/C vssd1 vssd1 vccd1 vccd1 _17351_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_71_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_546 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15515__A2 _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17279_ _17279_/A _17488_/A vssd1 vssd1 vccd1 vccd1 _17294_/A sky130_fd_sc_hd__and2_1
XFILLER_0_31_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19018_ _19019_/A _19019_/B vssd1 vssd1 vccd1 vccd1 _19190_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_67_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20290_ _20290_/A _20290_/B vssd1 vssd1 vccd1 vccd1 _20292_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18849__D _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12897__D _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout372_A _21775_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17976__B1 _21847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_1184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_1168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21813_ _21816_/CLK _21813_/D vssd1 vssd1 vccd1 vccd1 hold323/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout637_A _11089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_936 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21744_ _22005_/CLK _21744_/D vssd1 vssd1 vccd1 vccd1 _21744_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_149_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17778__A _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21675_ _21939_/CLK _21675_/D vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13765__A1 _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20626_ _20623_/X _20624_/Y _20491_/B _20492_/Y vssd1 vssd1 vccd1 vccd1 _20627_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_149_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19993__A _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13923__A2_N _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16832__D _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20557_ _20742_/B _20557_/B vssd1 vssd1 vccd1 vccd1 _20572_/A sky130_fd_sc_hd__and2_1
XFILLER_0_149_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17900__B1 _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14714__B1 _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11290_ _11493_/A1 t1x[16] v2z[16] _11507_/B2 _11289_/X vssd1 vssd1 vccd1 vccd1 _11290_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20488_ _20485_/Y _20486_/X _20337_/Y _20339_/Y vssd1 vssd1 vccd1 vccd1 _20488_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14930__A _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21109_ _21110_/A _21110_/B _21110_/C vssd1 vssd1 vccd1 vccd1 _21109_/Y sky130_fd_sc_hd__a21oi_2
X_14980_ _14859_/A _21755_/Q _14981_/C _15075_/A vssd1 vssd1 vccd1 vccd1 _14982_/B
+ sky130_fd_sc_hd__a22o_1
X_22089_ _22096_/CLK _22089_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[25] sky130_fd_sc_hd__dfrtp_4
Xfanout150 _17417_/C vssd1 vssd1 vccd1 vccd1 _17041_/A sky130_fd_sc_hd__buf_4
XFILLER_0_22_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout161 _17324_/D vssd1 vssd1 vccd1 vccd1 _19951_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA_clkbuf_leaf_20_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout172 _21827_/Q vssd1 vssd1 vccd1 vccd1 _16870_/A sky130_fd_sc_hd__buf_2
X_13931_ _13931_/A _13931_/B _13931_/C vssd1 vssd1 vccd1 vccd1 _13933_/B sky130_fd_sc_hd__nand3_1
Xfanout183 _17666_/A vssd1 vssd1 vccd1 vccd1 _19587_/A sky130_fd_sc_hd__buf_4
Xfanout194 hold327/X vssd1 vssd1 vccd1 vccd1 _21056_/B sky130_fd_sc_hd__buf_4
XFILLER_0_156_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16650_ _16566_/A _16566_/C _16566_/B vssd1 vssd1 vccd1 vccd1 _16651_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__17431__A2 _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13862_ _14027_/A _14354_/C _14663_/D _13864_/B vssd1 vssd1 vccd1 vccd1 _13867_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15601_ _15458_/Y _15460_/Y _15599_/Y _15600_/X vssd1 vssd1 vccd1 vccd1 _15601_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_97_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12813_ _12813_/A _12813_/B _12813_/C vssd1 vssd1 vccd1 vccd1 _12816_/A sky130_fd_sc_hd__or3_1
X_16581_ _17199_/A _16580_/C _16580_/A vssd1 vssd1 vccd1 vccd1 _16582_/C sky130_fd_sc_hd__a21o_1
X_13793_ _13789_/X _13791_/Y _13638_/B _13638_/Y vssd1 vssd1 vccd1 vccd1 _13795_/D
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_85_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18320_ _18320_/A _18320_/B vssd1 vssd1 vccd1 vccd1 _18321_/B sky130_fd_sc_hd__nand2_1
X_15532_ _15717_/B _15913_/B _15533_/C _15714_/A vssd1 vssd1 vccd1 vccd1 _15534_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_273 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12744_ _12744_/A _12744_/B _12744_/C vssd1 vssd1 vccd1 vccd1 _12744_/Y sky130_fd_sc_hd__nor3_4
XANTENNA__13712__C _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18392__B1 _18390_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18251_ _18117_/A _18116_/B _18114_/Y vssd1 vssd1 vccd1 vccd1 _18267_/A sky130_fd_sc_hd__a21o_1
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12008__A1 _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15463_ _15464_/A _15464_/B _15464_/C vssd1 vssd1 vccd1 vccd1 _15463_/X sky130_fd_sc_hd__a21o_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16942__A1 _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16592__A _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12675_ _12785_/B _14384_/C _14384_/D _14248_/A vssd1 vssd1 vccd1 vccd1 _12676_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_139_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17202_ _17619_/B _17300_/C _17520_/D _17621_/C vssd1 vssd1 vccd1 vccd1 _17203_/B
+ sky130_fd_sc_hd__a22o_1
X_14414_ _14250_/B _14242_/X _14413_/X vssd1 vssd1 vccd1 vccd1 _14416_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18182_ _18183_/A _18183_/B _18183_/C vssd1 vssd1 vccd1 vccd1 _18220_/A sky130_fd_sc_hd__and3_1
X_11626_ _12094_/A _12443_/A _12642_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _11626_/Y
+ sky130_fd_sc_hd__a22oi_1
X_15394_ _16371_/A _16399_/A _16424_/A _15791_/A vssd1 vssd1 vccd1 vccd1 _15398_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17133_ _17133_/A _17133_/B vssd1 vssd1 vccd1 vccd1 _17134_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_53_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14345_ _14345_/A _14345_/B vssd1 vssd1 vccd1 vccd1 _14435_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__17200__B _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11557_ _12094_/A _12094_/B _12877_/B _12751_/B vssd1 vssd1 vccd1 vccd1 _11557_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_53_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15001__A _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17064_ _17145_/A _17123_/C vssd1 vssd1 vccd1 vccd1 _17066_/B sky130_fd_sc_hd__and2_1
XFILLER_0_40_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14276_ _14273_/X _14274_/Y _14111_/Y _14113_/X vssd1 vssd1 vccd1 vccd1 _14277_/C
+ sky130_fd_sc_hd__o211ai_4
X_11488_ _11487_/X _18767_/B _11521_/S vssd1 vssd1 vccd1 vccd1 _21834_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_150_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16015_ _16015_/A _16015_/B vssd1 vssd1 vccd1 vccd1 _16021_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13227_ hold219/X _13226_/X fanout3/X vssd1 vssd1 vccd1 vccd1 _21862_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_27_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17854__C _19051_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ _13157_/A _13157_/B _13298_/A _13157_/D vssd1 vssd1 vccd1 vccd1 _13160_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ _12110_/A _12108_/Y _12109_/C _12269_/D vssd1 vssd1 vccd1 vccd1 _12153_/A
+ sky130_fd_sc_hd__and4bb_1
X_17966_ _17966_/A _17966_/B vssd1 vssd1 vccd1 vccd1 _17967_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13089_ _13091_/A _13091_/B vssd1 vssd1 vccd1 vccd1 _13089_/X sky130_fd_sc_hd__and2b_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16917_ _17141_/A _17141_/B _16917_/C _16968_/C vssd1 vssd1 vccd1 vccd1 _16920_/A
+ sky130_fd_sc_hd__nand4_2
X_19705_ _20148_/C _19705_/B _19705_/C _19903_/A vssd1 vssd1 vccd1 vccd1 _19903_/B
+ sky130_fd_sc_hd__nand4_2
X_17897_ _17897_/A _17897_/B vssd1 vssd1 vccd1 vccd1 _17906_/A sky130_fd_sc_hd__xor2_1
X_19636_ _19636_/A _19636_/B vssd1 vssd1 vccd1 vccd1 _19636_/Y sky130_fd_sc_hd__nor2_1
X_16848_ _16849_/B _16849_/C _16849_/A vssd1 vssd1 vccd1 vccd1 _16855_/A sky130_fd_sc_hd__o21ai_2
X_19567_ _19868_/B _19566_/X _19565_/X vssd1 vssd1 vccd1 vccd1 _19569_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_125_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16779_ _16756_/Y _16776_/X _16777_/X _16712_/Y vssd1 vssd1 vccd1 vccd1 _16785_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_88_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_87_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18518_ _18368_/C _18367_/Y _18516_/X _18517_/Y vssd1 vssd1 vccd1 vccd1 _18521_/C
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_73_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19498_ _19341_/A _19340_/A _19340_/B _19336_/B _19336_/A vssd1 vssd1 vccd1 vccd1
+ _19499_/B sky130_fd_sc_hd__o32ai_4
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18449_ _18606_/A _18449_/B vssd1 vssd1 vccd1 vccd1 _18451_/B sky130_fd_sc_hd__and2_1
XFILLER_0_111_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20190__B1 _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13747__A1 _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13747__B2 _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21460_ hold139/X sstream_i[37] _21494_/S vssd1 vssd1 vccd1 vccd1 _21987_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_145_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20411_ _21291_/A _21296_/A _21278_/A _21301_/A vssd1 vssd1 vccd1 vccd1 _20603_/A
+ sky130_fd_sc_hd__nand4_2
X_21391_ _15070_/B _19944_/Y _21420_/S vssd1 vssd1 vccd1 vccd1 _21391_/X sky130_fd_sc_hd__mux2_1
XANTENNA_fanout120_A _20562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20342_ _20343_/A _20343_/B _20343_/C vssd1 vssd1 vccd1 vccd1 _20342_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_141_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20273_ _20273_/A _20419_/A _20273_/C _20273_/D vssd1 vssd1 vccd1 vccd1 _20421_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_80_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22012_ _22013_/CLK _22012_/D vssd1 vssd1 vccd1 vccd1 hold201/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__18579__D _18894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20796__A2 _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout587_A _11549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14475__A2 _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17780__B _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12420__D _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19053__A _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16396__B _16396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16621__B1 _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13435__B1 _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19988__A _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18892__A _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10790_ mstream_i vssd1 vssd1 vccd1 vccd1 _10790_/Y sky130_fd_sc_hd__inv_2
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout33_A _21490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20927__A _21267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15188__B1 _15046_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21727_ _22016_/CLK _21727_/D vssd1 vssd1 vccd1 vccd1 _21727_/Q sky130_fd_sc_hd__dfxtp_2
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16924__A1 _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16924__B2 _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21658_ _21934_/CLK _21658_/D vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__dfxtp_1
X_12460_ _12460_/A _12460_/B _12460_/C vssd1 vssd1 vccd1 vccd1 _12463_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_124_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11411_ _11447_/A1 hold301/A fanout47/X hold142/A vssd1 vssd1 vccd1 vccd1 _11411_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12391_ _12391_/A _12497_/A vssd1 vssd1 vccd1 vccd1 _12392_/B sky130_fd_sc_hd__xnor2_4
X_20609_ _20609_/A _20729_/B vssd1 vssd1 vccd1 vccd1 _20611_/B sky130_fd_sc_hd__or2_1
XFILLER_0_151_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21589_ _21888_/CLK _21589_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[52] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14130_ _14015_/A _14015_/C _14015_/B vssd1 vssd1 vccd1 vccd1 _14277_/A sky130_fd_sc_hd__a21bo_1
X_11342_ _11544_/A1 t1x[29] v2z[29] _11543_/B2 _11341_/X vssd1 vssd1 vccd1 vccd1 _11342_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_105_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14061_ _14062_/B _14062_/C _14062_/A vssd1 vssd1 vccd1 vccd1 _14064_/A sky130_fd_sc_hd__a21o_1
X_11273_ _11325_/A1 t2y[12] t0y[12] _11498_/A1 vssd1 vssd1 vccd1 vccd1 _11273_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_120_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13012_ _13867_/A _13012_/B vssd1 vssd1 vccd1 vccd1 _13016_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_982 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17820_ _17819_/B _17819_/C _17819_/A vssd1 vssd1 vccd1 vccd1 _17821_/B sky130_fd_sc_hd__a21o_1
XANTENNA__17971__A _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17751_ _17750_/B _17750_/C _17750_/A vssd1 vssd1 vccd1 vccd1 _17751_/Y sky130_fd_sc_hd__a21oi_2
X_14963_ _14959_/X _14960_/Y _14795_/X _14797_/Y vssd1 vssd1 vccd1 vccd1 _14964_/B
+ sky130_fd_sc_hd__a211oi_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16587__A _21825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16702_ _16701_/A _16701_/C _16701_/B vssd1 vssd1 vccd1 vccd1 _16705_/B sky130_fd_sc_hd__a21o_1
X_13914_ _14859_/A _14391_/B _13915_/C _14073_/A vssd1 vssd1 vccd1 vccd1 _13916_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17682_ _17681_/A _17681_/B _17681_/C vssd1 vssd1 vccd1 vccd1 _17684_/C sky130_fd_sc_hd__a21o_1
X_14894_ _14743_/A _14743_/B _14741_/X vssd1 vssd1 vccd1 vccd1 _14896_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__16612__B1 _17334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19421_ _19563_/A _19420_/C _19420_/A vssd1 vssd1 vccd1 vccd1 _19422_/C sky130_fd_sc_hd__a21o_1
X_16633_ _16634_/A _16634_/B _16634_/C vssd1 vssd1 vccd1 vccd1 _16633_/X sky130_fd_sc_hd__and3_1
X_13845_ _13846_/A _13846_/B _13846_/C vssd1 vssd1 vccd1 vccd1 _13845_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_0_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19352_ _20032_/D _20193_/D _19353_/C _19504_/A vssd1 vssd1 vccd1 vccd1 _19354_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16564_ _16564_/A _16564_/B vssd1 vssd1 vccd1 vccd1 _16566_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13776_ _14572_/A _15098_/B vssd1 vssd1 vccd1 vccd1 _13779_/A sky130_fd_sc_hd__and2_1
XANTENNA__13442__C _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10988_ _10988_/A _10988_/B vssd1 vssd1 vccd1 vccd1 _10988_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_58_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18303_ _18304_/A _18304_/B _18304_/C vssd1 vssd1 vccd1 vccd1 _18305_/A sky130_fd_sc_hd__a21oi_4
X_15515_ _15514_/A _15514_/B _16173_/B vssd1 vssd1 vccd1 vccd1 _15516_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_139_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19283_ _19282_/B _19427_/B _19282_/A vssd1 vssd1 vccd1 vccd1 _19284_/B sky130_fd_sc_hd__a21o_1
X_12727_ _12851_/B _12727_/B vssd1 vssd1 vccd1 vccd1 _12730_/A sky130_fd_sc_hd__or2_2
X_16495_ _16495_/A _16495_/B vssd1 vssd1 vccd1 vccd1 _16781_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_139_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18234_ _18234_/A _18386_/A _18234_/C vssd1 vssd1 vccd1 vccd1 _18386_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_26_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12058__C _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15446_ _15446_/A _15446_/B vssd1 vssd1 vccd1 vccd1 _15449_/B sky130_fd_sc_hd__xnor2_2
X_12658_ _12563_/A _12562_/B _12562_/A vssd1 vssd1 vccd1 vccd1 _12665_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_154_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18165_ _19892_/A _18929_/B _18616_/D _19230_/A vssd1 vssd1 vccd1 vccd1 _18167_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11609_ _11887_/A _11887_/B vssd1 vssd1 vccd1 vccd1 _11609_/X sky130_fd_sc_hd__and2_1
X_15377_ _15377_/A _15377_/B vssd1 vssd1 vccd1 vccd1 _15379_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_5_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19865__B1 _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12589_ _12479_/C _12479_/Y _12587_/X _12588_/X vssd1 vssd1 vccd1 vccd1 _12589_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17116_ _17111_/X _17159_/A _17158_/A vssd1 vssd1 vccd1 vccd1 _17117_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_25_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14328_ _14936_/D _15174_/D _14328_/C _14474_/A vssd1 vssd1 vccd1 vccd1 _14474_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18096_ _18095_/B _18095_/C _18095_/A vssd1 vssd1 vccd1 vccd1 _18096_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_25_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14154__A1 _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14154__B2 _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17047_ _17040_/X _17114_/A _17002_/Y _17009_/X vssd1 vssd1 vccd1 vccd1 _17049_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_25_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14259_ _14258_/A _14258_/B _14258_/C vssd1 vssd1 vccd1 vccd1 _14260_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13186__A _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17643__A2 _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18998_ _19160_/B _18999_/C _18999_/A vssd1 vssd1 vccd1 vccd1 _19000_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__15654__A1 _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18696__B _19008_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17949_ _17948_/B _17948_/C _17948_/A vssd1 vssd1 vccd1 vccd1 _17949_/Y sky130_fd_sc_hd__o21ai_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20960_ _20960_/A _20960_/B _20960_/C vssd1 vssd1 vccd1 vccd1 _20960_/X sky130_fd_sc_hd__or3_2
XFILLER_0_139_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19619_ _19620_/A _19620_/B vssd1 vssd1 vccd1 vccd1 _19619_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_71_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13417__B1 _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20891_ _20888_/Y _20889_/X _20757_/X _20759_/Y vssd1 vssd1 vccd1 vccd1 _20892_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__15551__D _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout168_A _19732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13968__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19601__A _19732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13968__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12249__B _21727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12640__A1 _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout335_A _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21512_ hold228/X sstream_i[89] _21528_/S vssd1 vssd1 vccd1 vccd1 _22039_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_35_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21443_ hold267/X sstream_i[20] _21490_/S vssd1 vssd1 vccd1 vccd1 _21970_/D sky130_fd_sc_hd__mux2_1
XANTENNA_fanout502_A _21744_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21374_ _21420_/S _14126_/X _21403_/S vssd1 vssd1 vccd1 vccd1 _21374_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20325_ _20325_/A _20325_/B vssd1 vssd1 vccd1 vccd1 _20328_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15893__A1 _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20256_ _20256_/A _20256_/B vssd1 vssd1 vccd1 vccd1 _20258_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19990__B _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17791__A _21824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20187_ _20000_/A _20000_/B _19999_/A vssd1 vssd1 vccd1 vccd1 _20200_/A sky130_fd_sc_hd__o21a_1
XTAP_3802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13120__A2 _21776_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11960_ _11960_/A _11960_/B _11960_/C vssd1 vssd1 vccd1 vccd1 _11960_/X sky130_fd_sc_hd__and3_1
XTAP_3835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18595__B1 _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10911_ _10911_/A _10911_/B _10911_/C vssd1 vssd1 vccd1 vccd1 _10912_/B sky130_fd_sc_hd__or3_1
XTAP_3868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11891_ _11899_/A _11889_/Y _11880_/X _11886_/X vssd1 vssd1 vccd1 vccd1 _11892_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_6_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13630_ _13630_/A _13630_/B _13630_/C vssd1 vssd1 vccd1 vccd1 _13632_/B sky130_fd_sc_hd__nand3_1
X_10842_ _10817_/Y _10835_/Y _10837_/X _11059_/B _11057_/A vssd1 vssd1 vccd1 vccd1
+ _10843_/C sky130_fd_sc_hd__a311o_1
XFILLER_0_128_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13561_ _13558_/Y _13714_/A _21734_/Q _16273_/A vssd1 vssd1 vccd1 vccd1 _13714_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_6_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18772__D _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19230__B _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_928 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15300_ _15702_/D _15435_/A _15829_/C _15954_/D vssd1 vssd1 vccd1 vccd1 _15437_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_82_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12512_ _12512_/A _12621_/C _12858_/C _12991_/D vssd1 vssd1 vccd1 vccd1 _12512_/X
+ sky130_fd_sc_hd__and4_1
X_16280_ _16181_/A _16181_/B _16179_/X vssd1 vssd1 vccd1 vccd1 _16291_/A sky130_fd_sc_hd__a21bo_1
XANTENNA__20990__A2_N _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13492_ _13491_/A _13491_/B _13491_/C _13491_/D vssd1 vssd1 vccd1 vccd1 _13492_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_109_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15231_ _16027_/A _16266_/C _15231_/C _15407_/A vssd1 vssd1 vccd1 vccd1 _15407_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13187__A2 _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17966__A _17966_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12443_ _12443_/A _12899_/B vssd1 vssd1 vccd1 vccd1 _12447_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_87_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16870__A _16870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20457__A1 _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15162_ _15162_/A _15162_/B vssd1 vssd1 vccd1 vccd1 _15163_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_90_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12374_ _12369_/X _12371_/Y _11753_/B _11753_/Y vssd1 vssd1 vccd1 vccd1 _12375_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14113_ _14113_/A _14113_/B _14111_/Y _14112_/X vssd1 vssd1 vccd1 vccd1 _14113_/X
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_132_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11325_ _11325_/A1 t2y[25] t0y[25] _11089_/B vssd1 vssd1 vccd1 vccd1 _11325_/X sky130_fd_sc_hd__a22o_1
X_15093_ _16027_/A _15093_/B vssd1 vssd1 vccd1 vccd1 _15094_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17873__A2 _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19970_ _19970_/A _19970_/B vssd1 vssd1 vccd1 vccd1 _19977_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_132_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14044_ _14043_/A _14043_/B _14043_/C vssd1 vssd1 vccd1 vccd1 _14045_/C sky130_fd_sc_hd__a21oi_1
X_11256_ _12155_/B _11255_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21765_/D sky130_fd_sc_hd__mux2_1
X_18921_ _18780_/X _18817_/A _19049_/B _18920_/Y vssd1 vssd1 vccd1 vccd1 _19007_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__20542__D _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14540__D _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18852_ _18854_/A _19017_/B vssd1 vssd1 vccd1 vccd1 _18855_/A sky130_fd_sc_hd__nor2_1
X_11187_ hold267/X fanout51/X fanout47/X hold235/A vssd1 vssd1 vccd1 vccd1 _11187_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17803_ _17802_/A _17802_/B _17802_/C vssd1 vssd1 vccd1 vccd1 _17805_/C sky130_fd_sc_hd__a21o_1
XANTENNA__15933__B _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18783_ _18780_/X _18781_/Y _18627_/Y _18629_/X vssd1 vssd1 vccd1 vccd1 _18817_/B
+ sky130_fd_sc_hd__o211a_1
X_15995_ _15992_/A _15993_/Y _15819_/Y _15823_/B vssd1 vssd1 vccd1 vccd1 _15996_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_89_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17734_ _17734_/A _17734_/B vssd1 vssd1 vccd1 vccd1 _17736_/B sky130_fd_sc_hd__xor2_2
X_14946_ _14946_/A _14946_/B vssd1 vssd1 vccd1 vccd1 _14954_/A sky130_fd_sc_hd__nand2_1
XANTENNA__17206__A _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17665_ _19587_/B _17915_/D _17924_/B _19587_/A vssd1 vssd1 vccd1 vccd1 _17665_/Y
+ sky130_fd_sc_hd__a22oi_1
X_14877_ _21769_/Q _16266_/C _14878_/C _14878_/D vssd1 vssd1 vccd1 vccd1 _14877_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16061__A1 _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16616_ _16615_/A _16615_/B _16615_/C vssd1 vssd1 vccd1 vccd1 _16617_/C sky130_fd_sc_hd__a21o_1
XANTENNA__18963__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19404_ _19404_/A _19404_/B vssd1 vssd1 vccd1 vccd1 _19405_/B sky130_fd_sc_hd__nor2_1
X_13828_ _13828_/A _13828_/B vssd1 vssd1 vccd1 vccd1 _13831_/A sky130_fd_sc_hd__xor2_1
XANTENNA__13172__C _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17596_ _21142_/A _21343_/B vssd1 vssd1 vccd1 vccd1 _17596_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_85_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16547_ _16547_/A _16547_/B vssd1 vssd1 vccd1 vccd1 _16548_/B sky130_fd_sc_hd__and2_1
X_19335_ _19013_/C _19179_/X _19182_/A _19182_/B vssd1 vssd1 vccd1 vccd1 _19336_/B
+ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13759_ _13599_/Y _13601_/X _13757_/X _13758_/Y vssd1 vssd1 vccd1 vccd1 _13795_/A
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__20145__B1 _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14565__A _14712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19266_ _19266_/A _19266_/B _19266_/C vssd1 vssd1 vccd1 vccd1 _19406_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_127_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16478_ _16478_/A _16478_/B vssd1 vssd1 vccd1 vccd1 _16485_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16364__A2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16696__A2_N _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18217_ _18077_/B _18077_/Y _18214_/X _18216_/Y vssd1 vssd1 vccd1 vccd1 _18220_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_54_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15429_ _15426_/Y _15427_/X _15251_/Y _15291_/Y vssd1 vssd1 vccd1 vccd1 _15475_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_116_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19197_ _20178_/D _19053_/B _19050_/X _19051_/X _18894_/B vssd1 vssd1 vccd1 vccd1
+ _19202_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_66_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18148_ _18293_/A _18147_/Y _19644_/A _19240_/B vssd1 vssd1 vccd1 vccd1 _18293_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_25_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold203 hold203/A vssd1 vssd1 vccd1 vccd1 hold203/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14127__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold214 hold214/A vssd1 vssd1 vccd1 vccd1 hold214/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14127__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20733__C _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_clk_i _21822_/CLK vssd1 vssd1 vccd1 vccd1 _22016_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18079_ _17943_/B _17943_/Y _18076_/X _18078_/Y vssd1 vssd1 vccd1 vccd1 _18082_/B
+ sky130_fd_sc_hd__a211oi_4
Xhold225 hold225/A vssd1 vssd1 vccd1 vccd1 hold225/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 hold236/A vssd1 vssd1 vccd1 vccd1 hold236/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold247 hold247/A vssd1 vssd1 vccd1 vccd1 hold247/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__B1 _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold258 hold258/A vssd1 vssd1 vccd1 vccd1 hold258/X sky130_fd_sc_hd__buf_4
X_20110_ _20110_/A _20110_/B vssd1 vssd1 vccd1 vccd1 _20112_/B sky130_fd_sc_hd__nand2_1
Xhold269 hold269/A vssd1 vssd1 vccd1 vccd1 hold269/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21090_ _21090_/A _21090_/B vssd1 vssd1 vccd1 vccd1 _21091_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__19066__A1 _19087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14623__A1_N _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19066__B2 _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20041_ _20041_/A _20041_/B vssd1 vssd1 vccd1 vccd1 _20059_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_141_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15627__A1 _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15627__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16939__B _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18857__D _19185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout285_A _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21992_ _22020_/CLK _21992_/D vssd1 vssd1 vccd1 vccd1 hold210/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__14459__B _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_109 sstream_i[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20943_ _21171_/A _21256_/B _20944_/C _20944_/D vssd1 vssd1 vccd1 vccd1 _20946_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12861__A1 _13554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20923__A2 _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19331__A _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20874_ _20870_/Y _20872_/X _20737_/Y _20739_/Y vssd1 vssd1 vccd1 vccd1 _20874_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_72_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20687__A1 _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20687__B2 _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14366__A1 _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20924__B _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21426_ hold230/X sstream_i[3] _21489_/S vssd1 vssd1 vccd1 vccd1 _21953_/D sky130_fd_sc_hd__mux2_1
XANTENNA__17304__A1 _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10927__A1 _10926_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21357_ hold63/X _21381_/B _21356_/X vssd1 vssd1 vccd1 vccd1 _21926_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_20_817 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11110_ _10919_/X hold64/X _11121_/S vssd1 vssd1 vccd1 vccd1 _21704_/D sky130_fd_sc_hd__mux2_1
X_20308_ _20721_/D _21286_/B _21296_/B _20590_/D vssd1 vssd1 vccd1 vccd1 _20312_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12090_ _12261_/A _12639_/A _12530_/A _12269_/B vssd1 vssd1 vccd1 vccd1 _12091_/C
+ sky130_fd_sc_hd__a22o_1
X_21288_ _21264_/A _21283_/A _21150_/X _21151_/X _21046_/B vssd1 vssd1 vccd1 vccd1
+ _21290_/A sky130_fd_sc_hd__a32o_1
X_11041_ _11041_/A _21725_/D vssd1 vssd1 vccd1 vccd1 _11084_/S sky130_fd_sc_hd__nand2_2
XFILLER_0_120_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20239_ _20239_/A _20239_/B vssd1 vssd1 vccd1 vccd1 _20260_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__18280__A2 _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17671__D _18789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14800_ _14800_/A _14800_/B vssd1 vssd1 vccd1 vccd1 _14802_/B sky130_fd_sc_hd__nor2_1
XANTENNA__13554__A _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15780_ _16036_/A _15780_/B vssd1 vssd1 vccd1 vccd1 _15907_/B sky130_fd_sc_hd__nor2_1
XTAP_3610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12992_ _21735_/Q _13269_/C _13269_/D _13858_/B vssd1 vssd1 vccd1 vccd1 _12993_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21167__A2 _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12301__B1 _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14731_ _14730_/B _14854_/B _14730_/A vssd1 vssd1 vccd1 vccd1 _14732_/C sky130_fd_sc_hd__a21o_1
XTAP_3654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11943_ _11927_/X _11941_/X _11942_/X _11870_/Y vssd1 vssd1 vccd1 vccd1 _11964_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_3665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17450_ _17450_/A _17450_/B _17450_/C vssd1 vssd1 vccd1 vccd1 _17453_/A sky130_fd_sc_hd__nand3_1
XTAP_3698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14662_ _16374_/A _16203_/D _14817_/C _14817_/D vssd1 vssd1 vccd1 vccd1 _14662_/X
+ sky130_fd_sc_hd__and4_1
XTAP_2953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14054__B1 _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11874_ _11874_/A _11874_/B vssd1 vssd1 vccd1 vccd1 _11881_/A sky130_fd_sc_hd__xnor2_1
XTAP_2975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_16401_ _16377_/A _16268_/B _16265_/X _16266_/X _16414_/B vssd1 vssd1 vccd1 vccd1
+ _16403_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_131_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21623__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13613_ _15217_/A _14212_/D _13613_/C _13613_/D vssd1 vssd1 vccd1 vccd1 _13614_/B
+ sky130_fd_sc_hd__and4_1
XTAP_2997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17381_ _17381_/A _17381_/B _17381_/C vssd1 vssd1 vccd1 vccd1 _17483_/C sky130_fd_sc_hd__or3_1
XANTENNA__20127__B1 _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10825_ hold113/A hold134/A vssd1 vssd1 vccd1 vccd1 _11047_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_156_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14593_ _14439_/A _14439_/B _14437_/X vssd1 vssd1 vccd1 vccd1 _14595_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_82_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19120_ _19120_/A _19120_/B vssd1 vssd1 vccd1 vccd1 _19130_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_67_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16332_ _16330_/Y _16332_/B vssd1 vssd1 vccd1 vccd1 _16333_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_109_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13544_ _13540_/Y _13542_/X _13387_/X _13389_/Y vssd1 vssd1 vccd1 vccd1 _13545_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_94_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19895__B _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19051_ _19051_/A _20026_/B _19051_/C vssd1 vssd1 vccd1 vccd1 _19051_/X sky130_fd_sc_hd__and3_1
X_16263_ _16183_/A _16183_/B _16184_/X vssd1 vssd1 vccd1 vccd1 _16297_/A sky130_fd_sc_hd__o21ba_1
X_13475_ _13475_/A _13475_/B _13475_/C vssd1 vssd1 vccd1 vccd1 _13478_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_129_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18002_ _18002_/A _18002_/B _18002_/C vssd1 vssd1 vccd1 vccd1 _18004_/A sky130_fd_sc_hd__and3_1
XFILLER_0_153_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15214_ _15167_/A _15167_/B _15165_/Y vssd1 vssd1 vccd1 vccd1 _15351_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_35_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12426_ _12750_/A _12426_/B vssd1 vssd1 vccd1 vccd1 _12430_/A sky130_fd_sc_hd__nand2_1
X_16194_ _16193_/A _16193_/B _16193_/C vssd1 vssd1 vccd1 vccd1 _16240_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_51_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15145_ _15298_/A _15143_/X _15041_/Y _15043_/X vssd1 vssd1 vccd1 vccd1 _15146_/D
+ sky130_fd_sc_hd__a211o_1
X_12357_ _12458_/A _13173_/C _12357_/C _13034_/D vssd1 vssd1 vccd1 vccd1 _12359_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11308_ _14018_/C _11307_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21778_/D sky130_fd_sc_hd__mux2_1
X_15076_ _15076_/A _15076_/B _16173_/B vssd1 vssd1 vccd1 vccd1 _15361_/A sky130_fd_sc_hd__nand3_4
X_19953_ _20087_/A _19955_/D vssd1 vssd1 vccd1 vccd1 _20089_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12288_ _12294_/B _12288_/B _12288_/C vssd1 vssd1 vccd1 vccd1 _12289_/B sky130_fd_sc_hd__and3_2
XFILLER_0_120_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14027_ _14027_/A _14817_/D _14027_/C _14027_/D vssd1 vssd1 vccd1 vccd1 _14027_/Y
+ sky130_fd_sc_hd__nand4_1
X_18904_ _18902_/X _18904_/B vssd1 vssd1 vccd1 vccd1 _18905_/B sky130_fd_sc_hd__and2b_1
X_11239_ fanout59/X v0z[3] fanout19/X _11238_/X vssd1 vssd1 vccd1 vccd1 _11239_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__18958__C _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19884_ _19885_/A _19885_/B _19885_/C _19885_/D vssd1 vssd1 vccd1 vccd1 _19884_/Y
+ sky130_fd_sc_hd__nor4_1
XANTENNA__11343__A1 _21407_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18835_ _18837_/A _18837_/B vssd1 vssd1 vccd1 vccd1 _18835_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__16282__A1 _16173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15978_ _16101_/A _15978_/B _16196_/A _15978_/D vssd1 vssd1 vccd1 vccd1 _16101_/B
+ sky130_fd_sc_hd__and4b_1
X_18766_ _19535_/A _19087_/B _19089_/B _18767_/B vssd1 vssd1 vccd1 vccd1 _18766_/X
+ sky130_fd_sc_hd__a22o_1
X_14929_ _15159_/D _15698_/B _14930_/C _14930_/D vssd1 vssd1 vccd1 vccd1 _14934_/A
+ sky130_fd_sc_hd__a22o_1
X_17717_ _17718_/A _17718_/B _17718_/C vssd1 vssd1 vccd1 vccd1 _17962_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__19220__A1 _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19220__B2 _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11646__A2 _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18697_ _18857_/B _19181_/B _18695_/Y _18853_/A vssd1 vssd1 vccd1 vccd1 _18701_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17648_ _17648_/A _17648_/B vssd1 vssd1 vccd1 vccd1 _17650_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_33_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16925__D _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17579_ _17602_/B _17580_/B _17580_/C _17580_/D vssd1 vssd1 vccd1 vccd1 _17579_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__21315__C1 _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19318_ _19318_/A _19318_/B vssd1 vssd1 vccd1 vccd1 _19320_/C sky130_fd_sc_hd__xor2_1
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20590_ _20462_/D _21293_/B _20721_/C _20590_/D vssd1 vssd1 vccd1 vccd1 _20593_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_46_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18731__B1 _18894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21330__A2 _11549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19249_ _19248_/B _19248_/C _19248_/A vssd1 vssd1 vccd1 vccd1 _19249_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_983 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12246__C _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19287__A1 _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15838__B _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21211_ _21311_/A _21305_/A _21283_/B _21305_/B vssd1 vssd1 vccd1 vccd1 _21212_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout200_A _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11582__A1 _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21142_ _21142_/A _21142_/B vssd1 vssd1 vccd1 vccd1 _21142_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__11582__B2 _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout502 _21744_/Q vssd1 vssd1 vccd1 vccd1 _16406_/A sky130_fd_sc_hd__clkbuf_4
Xfanout513 _21741_/Q vssd1 vssd1 vccd1 vccd1 _16092_/D sky130_fd_sc_hd__buf_4
X_21073_ _21228_/A _21071_/X _20952_/B _20953_/Y vssd1 vssd1 vccd1 vccd1 _21075_/C
+ sky130_fd_sc_hd__o211a_1
Xfanout524 _21739_/Q vssd1 vssd1 vccd1 vccd1 _13877_/A sky130_fd_sc_hd__buf_4
XFILLER_0_67_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21397__A2 _15356_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout535 _12642_/A vssd1 vssd1 vccd1 vccd1 _12877_/B sky130_fd_sc_hd__buf_4
Xfanout546 _21734_/Q vssd1 vssd1 vccd1 vccd1 _13858_/B sky130_fd_sc_hd__clkbuf_8
X_20024_ _20024_/A _20024_/B vssd1 vssd1 vccd1 vccd1 _20066_/A sky130_fd_sc_hd__nand2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout557 _13556_/A vssd1 vssd1 vccd1 vccd1 _12512_/A sky130_fd_sc_hd__buf_4
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout568 _14312_/D vssd1 vssd1 vccd1 vccd1 _13682_/C sky130_fd_sc_hd__buf_4
Xfanout579 _13525_/A vssd1 vssd1 vccd1 vccd1 _13381_/C sky130_fd_sc_hd__buf_2
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11098__A0 _11061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13093__B _21352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11606__B _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21975_ _22016_/CLK _21975_/D vssd1 vssd1 vccd1 vccd1 hold293/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__16025__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16025__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20926_ _21258_/A _21046_/B _21278_/B _21267_/A vssd1 vssd1 vccd1 vccd1 _20930_/C
+ sky130_fd_sc_hd__a22o_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_1208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16576__A2 _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20857_ _20857_/A _20857_/B vssd1 vssd1 vccd1 vccd1 _20868_/A sky130_fd_sc_hd__or2_1
XFILLER_0_7_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12062__A2 _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11590_ _13012_/B _12302_/A _11589_/C _11589_/D vssd1 vssd1 vccd1 vccd1 _11591_/B
+ sky130_fd_sc_hd__a22oi_1
X_20788_ _20788_/A _20788_/B _20788_/C vssd1 vssd1 vccd1 vccd1 _20790_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_135_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18868__A4 _21847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_148_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15000__A2 _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13260_ _13554_/B _14018_/C _13411_/A _13260_/D vssd1 vssd1 vccd1 vccd1 _13411_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__19278__A1 _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19278__B2 _19430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17666__D _17924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12211_ _12203_/A _12203_/C _12203_/B vssd1 vssd1 vccd1 vccd1 _12211_/Y sky130_fd_sc_hd__o21ai_2
X_21409_ _21412_/A _21409_/B vssd1 vssd1 vccd1 vccd1 _21409_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13191_ _13191_/A _13191_/B _13191_/C vssd1 vssd1 vccd1 vccd1 _13193_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_20_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15839__B2 _14659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12142_ _12267_/A _12214_/C _12246_/C _12242_/B vssd1 vssd1 vccd1 vccd1 _12144_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_124_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16950_ _16943_/A _16943_/B _16936_/Y vssd1 vssd1 vccd1 vccd1 _16954_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_21_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12073_ _12073_/A _12080_/A vssd1 vssd1 vccd1 vccd1 _12075_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11325__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21388__A2 _14918_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11325__B2 _11089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15901_ _16031_/A _15901_/B vssd1 vssd1 vccd1 vccd1 _15902_/B sky130_fd_sc_hd__or2_1
X_11024_ mstream_o[98] hold239/X _11027_/S vssd1 vssd1 vccd1 vccd1 hold240/A sky130_fd_sc_hd__mux2_1
X_16881_ _16881_/A _16881_/B vssd1 vssd1 vccd1 vccd1 _16888_/A sky130_fd_sc_hd__xor2_1
X_15832_ _15961_/D _16404_/B _15832_/C _15832_/D vssd1 vssd1 vccd1 vccd1 _15959_/B
+ sky130_fd_sc_hd__and4_1
X_18620_ _18620_/A _18620_/B vssd1 vssd1 vccd1 vccd1 _18630_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_21_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15763_ _15763_/A _15763_/B vssd1 vssd1 vccd1 vccd1 _15764_/B sky130_fd_sc_hd__nand2_1
XTAP_3440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18551_ _18707_/A _18551_/B vssd1 vssd1 vccd1 vccd1 _18572_/A sky130_fd_sc_hd__or2_1
XFILLER_0_99_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12975_ _13682_/C _14176_/C _13402_/D _13822_/B vssd1 vssd1 vccd1 vccd1 _12976_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11628__A2 _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14714_ _14713_/A _14713_/B _16173_/B vssd1 vssd1 vccd1 vccd1 _14848_/C sky130_fd_sc_hd__o21a_2
X_17502_ _17619_/B _17621_/C _21056_/A _21169_/A vssd1 vssd1 vccd1 vccd1 _17618_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18482_ _19723_/A _19092_/C _18347_/B _18345_/X vssd1 vssd1 vccd1 vccd1 _18489_/A
+ sky130_fd_sc_hd__a31o_1
X_11926_ _11854_/A _11854_/B _11854_/C vssd1 vssd1 vccd1 vccd1 _11928_/C sky130_fd_sc_hd__a21o_1
X_15694_ _15695_/A _16084_/C _16084_/D _15961_/D vssd1 vssd1 vccd1 vccd1 _15698_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17764__A1 _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17764__B2 _19823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17433_ _17433_/A _19432_/A vssd1 vssd1 vccd1 vccd1 _17437_/A sky130_fd_sc_hd__nand2_1
X_14645_ _14800_/A _14643_/Y _14482_/B _14484_/B vssd1 vssd1 vccd1 vccd1 _14646_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _11857_/A _11857_/B _11857_/C vssd1 vssd1 vccd1 vccd1 _11870_/A sky130_fd_sc_hd__nand3_4
XFILLER_0_74_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19505__A2 _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10808_ hold219/A hold58/A vssd1 vssd1 vccd1 vccd1 _10810_/A sky130_fd_sc_hd__nand2_1
X_17364_ _17365_/A _17365_/B vssd1 vssd1 vccd1 vccd1 _17364_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_131_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14576_ _14576_/A _14576_/B vssd1 vssd1 vccd1 vccd1 _14579_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_83_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11788_ _11788_/A _11788_/B _11788_/C vssd1 vssd1 vccd1 vccd1 _11819_/A sky130_fd_sc_hd__nand3_2
X_16315_ _16315_/A _16400_/A vssd1 vssd1 vccd1 vccd1 _16316_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_103_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19103_ _19103_/A _19103_/B _19103_/C vssd1 vssd1 vccd1 vccd1 _19105_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_43_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13527_ _13527_/A _13527_/B vssd1 vssd1 vccd1 vccd1 _13536_/A sky130_fd_sc_hd__or2_1
XFILLER_0_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17295_ _17297_/A _17297_/B _17297_/C vssd1 vssd1 vccd1 vccd1 _17296_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_153_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_15_clk_i_A _21806_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20564__B _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19034_ _19031_/Y _19032_/X _18894_/D _18895_/B vssd1 vssd1 vccd1 vccd1 _19035_/C
+ sky130_fd_sc_hd__o211ai_2
X_16246_ _16132_/A _16133_/Y _16352_/B _16245_/X vssd1 vssd1 vccd1 vccd1 _16248_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_153_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15658__B _15916_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13458_ _15076_/A _15076_/B _14212_/D _14218_/B vssd1 vssd1 vccd1 vccd1 _13608_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_88_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13459__A _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13553__A2 _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12409_ _12410_/A _12410_/B vssd1 vssd1 vccd1 vccd1 _12521_/B sky130_fd_sc_hd__nand2_1
X_16177_ _16286_/A _16177_/B vssd1 vssd1 vccd1 vccd1 _16178_/B sky130_fd_sc_hd__nand2_1
X_13389_ _13390_/A _13390_/B vssd1 vssd1 vccd1 vccd1 _13389_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_88_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15128_ _14994_/A _14996_/B _14994_/B vssd1 vssd1 vccd1 vccd1 _15133_/A sky130_fd_sc_hd__a21boi_1
XANTENNA__15096__D _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15059_ _15059_/A _15059_/B vssd1 vssd1 vccd1 vccd1 _15060_/B sky130_fd_sc_hd__xnor2_1
X_19936_ _19937_/A _19937_/B vssd1 vssd1 vccd1 vccd1 _19936_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__18050__A _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11316__A1 _11315_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16489__B _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12513__B1 _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19867_ _19867_/A _19867_/B vssd1 vssd1 vccd1 vccd1 _19869_/A sky130_fd_sc_hd__nand2_1
X_18818_ _18817_/A _18817_/B _18815_/X _18816_/Y vssd1 vssd1 vccd1 vccd1 _18818_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__19992__A2 _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13625__C _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19798_ _19798_/A _19798_/B vssd1 vssd1 vccd1 vccd1 _19934_/A sky130_fd_sc_hd__or2_1
X_18749_ _19686_/A _19686_/B _19068_/C _20146_/B vssd1 vssd1 vccd1 vccd1 _18906_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_144_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14314__A2_N _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21760_ _21963_/CLK _21760_/D vssd1 vssd1 vccd1 vccd1 _21760_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_20_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21939_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__16558__A2 _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20711_ _20712_/A _20712_/B _20712_/C vssd1 vssd1 vccd1 vccd1 _20755_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_93_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21691_ _22080_/CLK _21691_/D vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15230__A2 _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout248_A _19379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_382 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20642_ _20513_/A _20509_/Y _20511_/B vssd1 vssd1 vccd1 vccd1 _20902_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11252__A0 _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_35_clk_i clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _22069_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_34_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20573_ _20707_/A _20572_/C _20572_/A vssd1 vssd1 vccd1 vccd1 _20573_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_128_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout415_A _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20193__C _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13369__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_1046 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18483__A2 _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21125_ _21232_/B _21123_/X _20964_/A _21014_/A vssd1 vssd1 vccd1 vccd1 _21125_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__19056__A _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12423__D _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout310 _21793_/Q vssd1 vssd1 vccd1 vccd1 _17490_/A sky130_fd_sc_hd__clkbuf_8
Xfanout321 _21791_/Q vssd1 vssd1 vccd1 vccd1 _18857_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__16399__B _16399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout332 _16409_/B vssd1 vssd1 vccd1 vccd1 _16084_/D sky130_fd_sc_hd__buf_4
Xfanout343 _21783_/Q vssd1 vssd1 vccd1 vccd1 _16418_/B sky130_fd_sc_hd__clkbuf_4
X_21056_ _21056_/A _21056_/B vssd1 vssd1 vccd1 vccd1 _21169_/B sky130_fd_sc_hd__and2_1
Xfanout354 _13402_/D vssd1 vssd1 vccd1 vccd1 _16414_/A sky130_fd_sc_hd__clkbuf_8
Xfanout365 _21777_/Q vssd1 vssd1 vccd1 vccd1 _13258_/D sky130_fd_sc_hd__buf_4
XANTENNA__12720__B _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout376 _14828_/B vssd1 vssd1 vccd1 vccd1 _13269_/D sky130_fd_sc_hd__clkbuf_4
X_20007_ _20007_/A _20007_/B _20143_/B vssd1 vssd1 vccd1 vccd1 _20154_/A sky130_fd_sc_hd__or3_1
Xfanout387 _15768_/A vssd1 vssd1 vccd1 vccd1 _14537_/A sky130_fd_sc_hd__buf_4
XANTENNA__18110__D _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11617__A _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout398 _14993_/A vssd1 vssd1 vccd1 vccd1 _15892_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout63_A _19185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14928__A _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12760_ _12642_/A _13157_/B _12645_/B _12643_/X vssd1 vssd1 vccd1 vccd1 _12762_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_139_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21958_ _21963_/CLK _21958_/D vssd1 vssd1 vccd1 vccd1 hold248/A sky130_fd_sc_hd__dfxtp_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11711_ _12443_/A _12897_/C _12897_/D _12642_/A vssd1 vssd1 vccd1 vccd1 _11711_/X
+ sky130_fd_sc_hd__and4_1
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20909_ hold145/X _20908_/X fanout2/X vssd1 vssd1 vccd1 vccd1 _21913_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12691_ _12692_/A _12692_/B _12692_/C _12692_/D vssd1 vssd1 vccd1 vccd1 _12691_/Y
+ sky130_fd_sc_hd__nor4_2
X_21889_ _21923_/CLK hold91/X vssd1 vssd1 vccd1 vccd1 hold90/A sky130_fd_sc_hd__dfxtp_1
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14430_ _14430_/A _14430_/B vssd1 vssd1 vccd1 vccd1 _14431_/B sky130_fd_sc_hd__xnor2_4
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11642_ _12426_/B _12403_/A _11576_/X _11577_/X _12619_/A vssd1 vssd1 vccd1 vccd1
+ _11643_/C sky130_fd_sc_hd__a32o_1
XANTENNA__14980__A1 _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14361_ _14361_/A _14361_/B vssd1 vssd1 vccd1 vccd1 _14375_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__15759__A fanout9/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11243__B1 _11242_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11573_ _11573_/A _11573_/B vssd1 vssd1 vccd1 vccd1 _11821_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18135__A _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16100_ _16100_/A _16100_/B vssd1 vssd1 vccd1 vccd1 _16119_/A sky130_fd_sc_hd__xnor2_2
X_13312_ _13310_/Y _13455_/A _15217_/A _14365_/D vssd1 vssd1 vccd1 vccd1 _13455_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_134_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17080_ _17038_/X _17060_/Y _17078_/A _17077_/Y vssd1 vssd1 vccd1 vccd1 _17081_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_52_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14292_ _14285_/B _14123_/C _14290_/X _14294_/C _13966_/A vssd1 vssd1 vccd1 vccd1
+ _14295_/A sky130_fd_sc_hd__a32oi_2
XFILLER_0_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_722 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21199__C _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22074__RESET_B fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16031_ _16031_/A _16031_/B vssd1 vssd1 vccd1 vccd1 _16032_/B sky130_fd_sc_hd__or2_1
X_13243_ _13243_/A _13243_/B vssd1 vssd1 vccd1 vccd1 _13245_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_66_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18789__B _18789_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13174_ _13173_/C _15217_/A _13171_/Y _13308_/A vssd1 vssd1 vccd1 vccd1 _13176_/C
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_62_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12125_ _12124_/A _12123_/Y _12076_/B _12084_/X vssd1 vssd1 vccd1 vccd1 _12127_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12911__A _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17982_ _17982_/A _17982_/B _17982_/C vssd1 vssd1 vccd1 vccd1 _18127_/C sky130_fd_sc_hd__nand3_2
X_19721_ _19721_/A _19721_/B vssd1 vssd1 vccd1 vccd1 _19769_/A sky130_fd_sc_hd__nor2_2
X_16933_ _16933_/A _16933_/B _16933_/C vssd1 vssd1 vccd1 vccd1 _16946_/A sky130_fd_sc_hd__and3_2
X_12056_ _12057_/A _12057_/B vssd1 vssd1 vccd1 vccd1 _12056_/X sky130_fd_sc_hd__and2_1
X_11007_ mstream_o[81] hold48/X _11012_/S vssd1 vssd1 vccd1 vccd1 _21618_/D sky130_fd_sc_hd__mux2_1
X_19652_ _19650_/D _20178_/B _21261_/B _19493_/D vssd1 vssd1 vccd1 vccd1 _19653_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_16864_ _16863_/B _16863_/C _16863_/A vssd1 vssd1 vccd1 vccd1 _16866_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_137_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18603_ _18603_/A _18603_/B vssd1 vssd1 vccd1 vccd1 _18606_/C sky130_fd_sc_hd__xnor2_2
X_15815_ _15815_/A _15815_/B _15815_/C vssd1 vssd1 vccd1 vccd1 _15816_/C sky130_fd_sc_hd__nand3_1
X_16795_ _17145_/A _16917_/C vssd1 vssd1 vccd1 vccd1 _16797_/B sky130_fd_sc_hd__and2_1
X_19583_ _19583_/A _19583_/B _19583_/C vssd1 vssd1 vccd1 vccd1 _19585_/A sky130_fd_sc_hd__and3_1
XANTENNA__19187__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13742__A _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14936__A_N _14774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15746_ _15743_/Y _15744_/X _15607_/X _15612_/C vssd1 vssd1 vccd1 vccd1 _15746_/X
+ sky130_fd_sc_hd__a211o_1
X_18534_ _18534_/A _18687_/A _18534_/C vssd1 vssd1 vccd1 vccd1 _18534_/Y sky130_fd_sc_hd__nand3_1
XTAP_3270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12958_ _12957_/B _12708_/X _12825_/X vssd1 vssd1 vccd1 vccd1 _12958_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_73_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14557__B _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13461__B _14212_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11909_ _11907_/A _11909_/B vssd1 vssd1 vccd1 vccd1 _12035_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_75_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15677_ _15678_/B _15678_/A vssd1 vssd1 vccd1 vccd1 _15815_/A sky130_fd_sc_hd__nand2b_1
X_18465_ _18465_/A _18465_/B vssd1 vssd1 vccd1 vccd1 _18475_/A sky130_fd_sc_hd__nand2_1
XANTENNA_270 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12889_ _12889_/A _13010_/A _12889_/C vssd1 vssd1 vccd1 vccd1 _13010_/B sky130_fd_sc_hd__nand3_2
XANTENNA_281 hold283/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_292 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14628_ _14629_/A _14629_/B vssd1 vssd1 vccd1 vccd1 _14630_/A sky130_fd_sc_hd__nor2_1
X_17416_ _17520_/A _20249_/A vssd1 vssd1 vccd1 vccd1 _17420_/A sky130_fd_sc_hd__nand2_1
X_18396_ _18100_/B _18394_/A _18242_/Y _18394_/C _18395_/X vssd1 vssd1 vccd1 vccd1
+ _18396_/Y sky130_fd_sc_hd__o41ai_4
XFILLER_0_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17347_ _17245_/A _17245_/C _17245_/B vssd1 vssd1 vccd1 vccd1 _17348_/C sky130_fd_sc_hd__a21bo_1
X_14559_ _14859_/A _15001_/B _14559_/C _14724_/A vssd1 vssd1 vccd1 vccd1 _14724_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_126_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17278_ _17278_/A vssd1 vssd1 vccd1 vccd1 _17488_/A sky130_fd_sc_hd__inv_2
XFILLER_0_125_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16229_ _16225_/Y _16226_/X _16109_/Y _16111_/Y vssd1 vssd1 vccd1 vccd1 _16229_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_113_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19017_ _19017_/A _19017_/B vssd1 vssd1 vccd1 vccd1 _19019_/B sky130_fd_sc_hd__or2_1
XFILLER_0_140_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11537__A1 _11089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11201__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19662__A1 _19531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19662__B2 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20272__A2 _20419_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19919_ _19759_/Y _19763_/C _19917_/X _19918_/Y vssd1 vssd1 vccd1 vccd1 _19919_/X
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17976__A1 _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17976__B2 _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19178__B1 _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout365_A _21777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17124__A _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21812_ _21816_/CLK _21812_/D vssd1 vssd1 vccd1 vccd1 hold328/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21743_ _22021_/CLK _21743_/D vssd1 vssd1 vccd1 vccd1 _21743_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_148_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12268__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout532_A _21737_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21674_ _21939_/CLK _21674_/D vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__17778__B _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_549 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21288__A1 _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13765__A2 _14218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21288__B2 _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20625_ _20491_/B _20492_/Y _20623_/X _20624_/Y vssd1 vssd1 vccd1 vccd1 _20627_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_47_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_950 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19350__B1 _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19993__B _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20556_ _20556_/A _20556_/B vssd1 vssd1 vccd1 vccd1 _20557_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17900__A1 _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17900__B2 _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14714__A1 _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11528__A1 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20487_ _20337_/Y _20339_/Y _20485_/Y _20486_/X vssd1 vssd1 vccd1 vccd1 _20487_/Y
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_120_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14930__B _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16467__A1 _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21108_ _21222_/B _21108_/B vssd1 vssd1 vccd1 vccd1 _21110_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_121_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout140 _21834_/Q vssd1 vssd1 vccd1 vccd1 _18929_/B sky130_fd_sc_hd__buf_4
X_22088_ _22096_/CLK _22088_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[24] sky130_fd_sc_hd__dfrtp_4
Xfanout151 _21831_/Q vssd1 vssd1 vccd1 vccd1 _17417_/C sky130_fd_sc_hd__buf_2
Xfanout162 _17324_/D vssd1 vssd1 vccd1 vccd1 _18787_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13930_ _13779_/A _13779_/B _13779_/C vssd1 vssd1 vccd1 vccd1 _13931_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_156_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21039_ _21040_/A _21264_/A _21040_/C _21040_/D vssd1 vssd1 vccd1 vccd1 _21041_/A
+ sky130_fd_sc_hd__a22oi_1
Xfanout173 _19723_/A vssd1 vssd1 vccd1 vccd1 _19439_/A sky130_fd_sc_hd__buf_4
Xfanout184 _17666_/A vssd1 vssd1 vccd1 vccd1 _19438_/A sky130_fd_sc_hd__buf_4
Xfanout195 _21171_/B vssd1 vssd1 vccd1 vccd1 _20247_/C sky130_fd_sc_hd__buf_4
X_13861_ _13861_/A _13861_/B vssd1 vssd1 vccd1 vccd1 _13871_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_92_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15600_ _15600_/A _15600_/B _15600_/C vssd1 vssd1 vccd1 vccd1 _15600_/X sky130_fd_sc_hd__and3_1
X_12812_ _12813_/A _12813_/B _12813_/C vssd1 vssd1 vccd1 vccd1 _12812_/Y sky130_fd_sc_hd__nor3_2
X_16580_ _16580_/A _17199_/A _16580_/C vssd1 vssd1 vccd1 vccd1 _17199_/B sky130_fd_sc_hd__nand3_1
X_13792_ _13638_/B _13638_/Y _13789_/X _13791_/Y vssd1 vssd1 vccd1 vccd1 _13795_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_97_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15531_ _16404_/A _16305_/B _15911_/A _15911_/C vssd1 vssd1 vccd1 vccd1 _15714_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__17969__A _17969_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12743_ _12743_/A _12743_/B _12743_/C vssd1 vssd1 vccd1 vccd1 _12744_/C sky130_fd_sc_hd__and3_1
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13712__D _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18392__B2 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18250_ _18250_/A _18250_/B vssd1 vssd1 vccd1 vccd1 _18275_/A sky130_fd_sc_hd__nand2_1
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15462_ _15464_/A _15464_/B _15464_/C vssd1 vssd1 vccd1 vccd1 _15462_/Y sky130_fd_sc_hd__a21oi_1
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12008__A2 _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12674_ _14248_/A _12785_/B _14384_/C _14384_/D vssd1 vssd1 vccd1 vccd1 _12676_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11216__A0 _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16942__A2 _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17201_ _17281_/A vssd1 vssd1 vccd1 vccd1 _17201_/Y sky130_fd_sc_hd__inv_2
XANTENNA__16592__B _16813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14413_ _14713_/B _15234_/C _14250_/B _14713_/A vssd1 vssd1 vccd1 vccd1 _14413_/X
+ sky130_fd_sc_hd__a22o_1
X_18181_ _18181_/A _18181_/B _18181_/C vssd1 vssd1 vccd1 vccd1 _18183_/C sky130_fd_sc_hd__nand3_2
X_11625_ _12094_/A _12094_/B _12443_/A _12877_/B vssd1 vssd1 vccd1 vccd1 _11625_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_53_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15393_ _15393_/A _15588_/B vssd1 vssd1 vccd1 vccd1 _15404_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_93_992 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17132_ _17133_/A _17132_/B _17132_/C vssd1 vssd1 vccd1 vccd1 _17133_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_53_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14344_ _14345_/A _14345_/B vssd1 vssd1 vccd1 vccd1 _14453_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_108_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11556_ _12094_/A _12242_/B _12751_/B vssd1 vssd1 vccd1 vccd1 _11556_/X sky130_fd_sc_hd__and3_1
XFILLER_0_80_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11231__A3 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17200__C _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17063_ _17146_/A _17146_/B _17063_/C _17086_/C vssd1 vssd1 vccd1 vccd1 _17066_/A
+ sky130_fd_sc_hd__nand4_2
X_14275_ _14111_/Y _14113_/X _14273_/X _14274_/Y vssd1 vssd1 vccd1 vccd1 _14277_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_64_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11487_ _11493_/A1 t2x[12] v1z[12] fanout20/X _11486_/X vssd1 vssd1 vccd1 vccd1 _11487_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__11519__A1 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16014_ _16014_/A _16014_/B vssd1 vssd1 vccd1 vccd1 _16015_/B sky130_fd_sc_hd__nand2_1
X_13226_ _21725_/D hold63/X _11061_/X fanout6/X _13225_/Y vssd1 vssd1 vccd1 vccd1
+ _13226_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_110_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17854__D _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13157_ _13157_/A _13157_/B _13298_/A _13157_/D vssd1 vssd1 vccd1 vccd1 _13298_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12671__A2_N _12781_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ _12229_/A _12246_/D _12269_/C _12155_/B vssd1 vssd1 vccd1 vccd1 _12108_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17965_ _17966_/B _17966_/A vssd1 vssd1 vccd1 vccd1 _18100_/A sky130_fd_sc_hd__nand2b_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ _13088_/A _13088_/B vssd1 vssd1 vccd1 vccd1 _13091_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_100_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19704_ _20148_/C _19705_/B _19705_/C _19903_/A vssd1 vssd1 vccd1 vccd1 _19706_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16916_ _16916_/A _16916_/B vssd1 vssd1 vccd1 vccd1 _16916_/Y sky130_fd_sc_hd__nand2_1
X_12039_ _12458_/A _12637_/B _12639_/A _12357_/C vssd1 vssd1 vccd1 vccd1 _12040_/C
+ sky130_fd_sc_hd__a22o_1
X_17896_ _18767_/B _17894_/X _17895_/X vssd1 vssd1 vccd1 vccd1 _17897_/B sky130_fd_sc_hd__a21bo_1
X_19635_ _19635_/A _19787_/B vssd1 vssd1 vccd1 vccd1 _21384_/B sky130_fd_sc_hd__xnor2_2
X_16847_ _16776_/X _16845_/Y _16844_/X _16826_/Y vssd1 vssd1 vccd1 vccd1 _16851_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_26_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13472__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12247__A2 _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19566_ _20101_/A _20101_/B _19906_/D vssd1 vssd1 vccd1 vccd1 _19566_/X sky130_fd_sc_hd__and3_1
X_16778_ _16756_/Y _16776_/X _16777_/X _16712_/Y vssd1 vssd1 vccd1 vccd1 _16778_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_125_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18517_ _18516_/A _18516_/B _18516_/C _18516_/D vssd1 vssd1 vccd1 vccd1 _18517_/Y
+ sky130_fd_sc_hd__o22ai_2
X_15729_ _15725_/Y _15727_/X _15595_/Y _15597_/Y vssd1 vssd1 vccd1 vccd1 _15729_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_87_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19497_ _19497_/A _19497_/B vssd1 vssd1 vccd1 vccd1 _19499_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18448_ _18445_/X _18594_/B _18314_/D _18316_/A vssd1 vssd1 vccd1 vccd1 _18449_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__20190__A1 _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20190__B2 _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11207__A0 _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13747__A2 _14212_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18379_ _18398_/B _18378_/B _18377_/C _18377_/D vssd1 vssd1 vccd1 vccd1 _18379_/Y
+ sky130_fd_sc_hd__a2bb2oi_2
XFILLER_0_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20410_ _21296_/A _21278_/A _21301_/A _21291_/A vssd1 vssd1 vccd1 vccd1 _20413_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16146__B1 _10972_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21390_ hold87/X _21390_/B vssd1 vssd1 vccd1 vccd1 _21390_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_16_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_344 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20341_ _20343_/A _20343_/B _20343_/C vssd1 vssd1 vccd1 vccd1 _20341_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout113_A _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20272_ _20273_/A _20419_/A _20273_/C _20273_/D vssd1 vssd1 vccd1 vccd1 _20274_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_80_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22011_ _22013_/CLK _22011_/D vssd1 vssd1 vccd1 vccd1 hold180/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__12551__A _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout482_A _21748_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19053__B _19053_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16621__A1 _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16621__B2 _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13435__A1 _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19988__B _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13435__B2 _13875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11446__A0 _11445_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18892__B _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20927__B _21841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21726_ _22016_/CLK _21726_/D vssd1 vssd1 vccd1 vccd1 _21726_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16924__A2 _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout26_A _11348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14417__S _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21657_ _21934_/CLK _21657_/D vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_81_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19323__B1 _14449_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11630__A _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11410_ _11409_/X _21293_/A _11446_/S vssd1 vssd1 vccd1 vccd1 _21808_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_34_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20608_ _20729_/A _21311_/B _21087_/D _20608_/D vssd1 vssd1 vccd1 vccd1 _20729_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_90_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12390_ _12496_/B _12390_/B vssd1 vssd1 vccd1 vccd1 _12497_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_62_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21588_ _21888_/CLK _21588_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[51] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11341_ _11349_/A1 t2y[29] t0y[29] _21723_/D vssd1 vssd1 vccd1 vccd1 _11341_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_50_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19509__A _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20539_ _20539_/A _20539_/B vssd1 vssd1 vccd1 vccd1 _20712_/A sky130_fd_sc_hd__and2_1
XFILLER_0_127_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14060_ _14859_/A _15373_/A _14873_/B _14217_/D vssd1 vssd1 vccd1 vccd1 _14062_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_132_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11272_ _12426_/B _11271_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21769_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_120_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13011_ _12904_/A _12903_/B _12901_/X vssd1 vssd1 vccd1 vccd1 _13027_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_30_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17029__A _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17971__B _21352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14962_ _14964_/A vssd1 vssd1 vccd1 vccd1 _14962_/Y sky130_fd_sc_hd__inv_2
X_17750_ _17750_/A _17750_/B _17750_/C vssd1 vssd1 vccd1 vccd1 _17750_/X sky130_fd_sc_hd__and3_2
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__16587__B _16734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16701_ _16701_/A _16701_/B _16701_/C vssd1 vssd1 vccd1 vccd1 _16705_/A sky130_fd_sc_hd__nand3_2
X_13913_ _14557_/A _14557_/B _13913_/C _14077_/B vssd1 vssd1 vccd1 vccd1 _14073_/A
+ sky130_fd_sc_hd__nand4_1
X_14893_ _14893_/A _14893_/B vssd1 vssd1 vccd1 vccd1 _14896_/A sky130_fd_sc_hd__xnor2_2
X_17681_ _17681_/A _17681_/B _17681_/C vssd1 vssd1 vccd1 vccd1 _17684_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_57_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16612__A1 _21822_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19420_ _19420_/A _19563_/A _19420_/C vssd1 vssd1 vccd1 vccd1 _19563_/B sky130_fd_sc_hd__nand3_1
X_13844_ _13844_/A _13844_/B vssd1 vssd1 vccd1 vccd1 _13846_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__16612__B2 _21823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16632_ _16631_/A _16631_/B _16631_/C vssd1 vssd1 vccd1 vccd1 _16634_/C sky130_fd_sc_hd__a21o_1
XANTENNA__14623__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11437__A0 _11436_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19351_ _20026_/B _20178_/D _20733_/C _20606_/D vssd1 vssd1 vccd1 vccd1 _19504_/A
+ sky130_fd_sc_hd__nand4_2
X_13775_ _13775_/A _13775_/B vssd1 vssd1 vccd1 vccd1 _13784_/A sky130_fd_sc_hd__xor2_1
X_16563_ _16563_/A _16586_/B _16563_/C vssd1 vssd1 vccd1 vccd1 _16566_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_58_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13442__D _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987_ hold232/A hold121/A vssd1 vssd1 vccd1 vccd1 _10988_/B sky130_fd_sc_hd__xnor2_2
X_18302_ _18302_/A _18302_/B vssd1 vssd1 vccd1 vccd1 _18304_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_1255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15514_ _15514_/A _15514_/B _16173_/B vssd1 vssd1 vccd1 vccd1 _15763_/B sky130_fd_sc_hd__and3_1
XFILLER_0_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12726_ _13822_/B _14018_/C _12725_/C _12725_/D vssd1 vssd1 vccd1 vccd1 _12727_/B
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_128_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16494_ _16484_/X _16492_/X _16493_/Y _16715_/A vssd1 vssd1 vccd1 vccd1 _16715_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19282_ _19282_/A _19282_/B _19427_/B vssd1 vssd1 vccd1 vccd1 _19282_/X sky130_fd_sc_hd__and3_1
XFILLER_0_73_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20172__A1 _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15445_ _15446_/A _15446_/B vssd1 vssd1 vccd1 vccd1 _15445_/Y sky130_fd_sc_hd__nand2_1
X_18233_ _18229_/X _18231_/Y _18091_/B _18091_/Y vssd1 vssd1 vccd1 vccd1 _18234_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12058__D _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12657_ _13013_/A _12899_/B _12553_/B _12551_/X vssd1 vssd1 vccd1 vccd1 _12667_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_155_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_154_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11608_ _11612_/B _11608_/B vssd1 vssd1 vccd1 vccd1 _11887_/B sky130_fd_sc_hd__nor2_1
X_15376_ _15376_/A _15376_/B vssd1 vssd1 vccd1 vccd1 _15379_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_128_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18164_ _18164_/A _18164_/B vssd1 vssd1 vccd1 vccd1 _18183_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19865__A1 _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ _12604_/B _12587_/B _12585_/Y _12586_/X vssd1 vssd1 vccd1 vccd1 _12588_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19865__B2 _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14327_ _14936_/D _15174_/D _14328_/C _14474_/A vssd1 vssd1 vccd1 vccd1 _14329_/B
+ sky130_fd_sc_hd__a22o_1
X_17115_ _17114_/A _17114_/B _17114_/C vssd1 vssd1 vccd1 vccd1 _17158_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_68_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18095_ _18095_/A _18095_/B _18095_/C vssd1 vssd1 vccd1 vccd1 _18095_/Y sky130_fd_sc_hd__nand3_4
X_11539_ _11538_/X _19181_/B _11545_/S vssd1 vssd1 vccd1 vccd1 _21851_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17046_ _17046_/A _17046_/B _17046_/C vssd1 vssd1 vccd1 vccd1 _17114_/A sky130_fd_sc_hd__or3_2
X_14258_ _14258_/A _14258_/B _14258_/C vssd1 vssd1 vccd1 vccd1 _14260_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_123_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14154__A2 _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13467__A _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13209_ _13230_/B _13209_/B _13209_/C _13209_/D vssd1 vssd1 vccd1 vccd1 _13209_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14189_ _14189_/A _14189_/B vssd1 vssd1 vccd1 vccd1 _14203_/A sky130_fd_sc_hd__xnor2_2
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13186__B _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18997_ _19160_/B _18999_/C vssd1 vssd1 vccd1 vccd1 _18997_/Y sky130_fd_sc_hd__nand2_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13114__B1 _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18696__C _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17948_ _17948_/A _17948_/B _17948_/C vssd1 vssd1 vccd1 vccd1 _17948_/X sky130_fd_sc_hd__or3_1
XFILLER_0_31_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17879_ _17878_/B _17878_/C _17878_/A vssd1 vssd1 vccd1 vccd1 _17881_/B sky130_fd_sc_hd__a21o_1
XANTENNA__11140__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19618_ _19457_/A _19457_/B _19455_/Y vssd1 vssd1 vccd1 vccd1 _19620_/B sky130_fd_sc_hd__a21boi_2
XANTENNA__13417__A1 _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20890_ _20757_/X _20759_/Y _20888_/Y _20889_/X vssd1 vssd1 vccd1 vccd1 _20892_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__14614__B1 _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13417__B2 _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11428__A0 _11427_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_926 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19549_ _19549_/A _19549_/B _19700_/B vssd1 vssd1 vccd1 vccd1 _19551_/B sky130_fd_sc_hd__nand3_1
XANTENNA__19601__B _19732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__22106__RESET_B _11089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12640__A2 _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21511_ hold271/X sstream_i[88] _21528_/S vssd1 vssd1 vccd1 vccd1 _22038_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_91_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21442_ hold301/X sstream_i[19] _21442_/S vssd1 vssd1 vccd1 vccd1 _21969_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_44_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21373_ _21420_/S _21373_/B vssd1 vssd1 vccd1 vccd1 _21373_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_82_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20324_ _20325_/A _20325_/B vssd1 vssd1 vccd1 vccd1 _20324_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_114_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15893__A2 _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20255_ _20255_/A _20255_/B vssd1 vssd1 vccd1 vccd1 _20256_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_110_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17791__B _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20186_ _20186_/A _20186_/B vssd1 vssd1 vccd1 vccd1 _20202_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12459__A2 _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold275_A hold275/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13824__B _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20926__B1 _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18595__A1 _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11131__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10910_ _10911_/A _10911_/B _10911_/C vssd1 vssd1 vccd1 vccd1 _10917_/B sky130_fd_sc_hd__o21a_1
XANTENNA__18595__B2 _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11890_ _11880_/X _11886_/X _11899_/A _11889_/Y vssd1 vssd1 vccd1 vccd1 _11899_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_54_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11419__A0 _11418_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10841_ _10843_/A _10841_/B vssd1 vssd1 vccd1 vccd1 _11059_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_6_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13560_ _13858_/B _16273_/A _13558_/Y _13714_/A vssd1 vssd1 vccd1 vccd1 _13562_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_137_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_1083 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12511_ _12511_/A _13573_/D vssd1 vssd1 vccd1 vccd1 _12515_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_137_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21709_ _22096_/CLK _21709_/D vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dfxtp_1
X_13491_ _13491_/A _13491_/B _13491_/C _13491_/D vssd1 vssd1 vccd1 vccd1 _13491_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_81_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15230_ _16027_/A _14234_/C _15231_/C _15407_/A vssd1 vssd1 vccd1 vccd1 _15232_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12442_ _12355_/A _12354_/A _12354_/B vssd1 vssd1 vccd1 vccd1 _12449_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16870__B _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15161_ _21734_/Q _15838_/B _16374_/B _21733_/Q vssd1 vssd1 vccd1 vccd1 _15162_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_90_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12373_ _12375_/C vssd1 vssd1 vccd1 vccd1 _12373_/Y sky130_fd_sc_hd__inv_2
X_14112_ _14109_/X _14110_/X _13948_/C _13947_/Y vssd1 vssd1 vccd1 vccd1 _14112_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_50_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11324_ _14477_/C _11323_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21782_/D sky130_fd_sc_hd__mux2_1
X_15092_ _15001_/B _15091_/X _15090_/X vssd1 vssd1 vccd1 vccd1 _15094_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14043_ _14043_/A _14043_/B _14043_/C vssd1 vssd1 vccd1 vccd1 _14045_/B sky130_fd_sc_hd__and3_1
X_18920_ _18919_/B _18919_/C _18919_/A vssd1 vssd1 vccd1 vccd1 _18920_/Y sky130_fd_sc_hd__o21ai_1
X_11255_ fanout59/X v0z[7] fanout19/X _11254_/X vssd1 vssd1 vccd1 vccd1 _11255_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_1190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1092 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18851_ _18848_/Y _19017_/A _18851_/C _19179_/C vssd1 vssd1 vccd1 vccd1 _19017_/B
+ sky130_fd_sc_hd__and4bb_1
X_11186_ _14386_/B _11185_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21745_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11370__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17802_ _17802_/A _17802_/B _17802_/C vssd1 vssd1 vccd1 vccd1 _17805_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_98_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18782_ _18627_/Y _18629_/X _18780_/X _18781_/Y vssd1 vssd1 vccd1 vccd1 _18817_/A
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__15933__C _15933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15994_ _15819_/Y _15823_/B _15992_/A _15993_/Y vssd1 vssd1 vccd1 vccd1 _16134_/A
+ sky130_fd_sc_hd__o211ai_4
X_17733_ _17734_/A _17734_/B vssd1 vssd1 vccd1 vccd1 _17847_/A sky130_fd_sc_hd__nand2b_1
X_14945_ _14824_/A _14823_/B _14821_/X vssd1 vssd1 vccd1 vccd1 _14956_/A sky130_fd_sc_hd__a21o_1
XANTENNA__17206__B _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17664_ _17664_/A _17664_/B vssd1 vssd1 vccd1 vccd1 _17684_/A sky130_fd_sc_hd__xnor2_2
X_14876_ _15514_/A _15514_/B _16414_/B _16391_/B vssd1 vssd1 vccd1 vccd1 _14878_/D
+ sky130_fd_sc_hd__nand4_4
XANTENNA__16061__A2 _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21443__S _21490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19403_ _19400_/X _19401_/Y _19271_/Y _19275_/A vssd1 vssd1 vccd1 vccd1 _19404_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16615_ _16615_/A _16615_/B _16615_/C vssd1 vssd1 vccd1 vccd1 _16617_/B sky130_fd_sc_hd__nand3_2
X_13827_ _13827_/A _13979_/B _13828_/B vssd1 vssd1 vccd1 vccd1 _13992_/A sky130_fd_sc_hd__or3b_2
XANTENNA__13172__D _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17595_ _17595_/A _17595_/B vssd1 vssd1 vccd1 vccd1 _17595_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__13750__A _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19334_ _19334_/A _19334_/B vssd1 vssd1 vccd1 vccd1 _19336_/A sky130_fd_sc_hd__xnor2_2
X_13758_ _13758_/A _13758_/B _13758_/C vssd1 vssd1 vccd1 vccd1 _13758_/Y sky130_fd_sc_hd__nor3_2
X_16546_ _16546_/A vssd1 vssd1 vccd1 vccd1 _16548_/A sky130_fd_sc_hd__inv_2
XANTENNA__20145__A1 _20562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20145__B2 _19906_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14565__B _14712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_586 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_2_1__f_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12709_ _12600_/A _12600_/B _12708_/X vssd1 vssd1 vccd1 vccd1 _12710_/B sky130_fd_sc_hd__a21boi_4
XFILLER_0_73_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19265_ _19095_/A _19095_/C _19095_/B vssd1 vssd1 vccd1 vccd1 _19266_/C sky130_fd_sc_hd__a21bo_1
X_13689_ _13689_/A vssd1 vssd1 vccd1 vccd1 _13689_/Y sky130_fd_sc_hd__inv_2
X_16477_ _16493_/A _16493_/B _16493_/C vssd1 vssd1 vccd1 vccd1 _16715_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_31_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18216_ _18215_/B _18215_/C _18215_/A vssd1 vssd1 vccd1 vccd1 _18216_/Y sky130_fd_sc_hd__a21oi_2
X_15428_ _15251_/Y _15291_/Y _15426_/Y _15427_/X vssd1 vssd1 vccd1 vccd1 _15475_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19196_ _20032_/D _19810_/D _19199_/C _21847_/Q _19032_/X vssd1 vssd1 vccd1 vccd1
+ _19204_/A sky130_fd_sc_hd__a41o_1
XFILLER_0_54_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20583__A _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15359_ hold109/X _15358_/X fanout4/X vssd1 vssd1 vccd1 vccd1 hold110/A sky130_fd_sc_hd__mux2_1
X_18147_ _19051_/A _19068_/C _19238_/C _20317_/D vssd1 vssd1 vccd1 vccd1 _18147_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_26_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold204 hold204/A vssd1 vssd1 vccd1 vccd1 hold204/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold215 hold215/A vssd1 vssd1 vccd1 vccd1 hold215/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__20733__D _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold226 hold226/A vssd1 vssd1 vccd1 vccd1 hold226/X sky130_fd_sc_hd__dlygate4sd3_1
X_18078_ _18077_/B _18077_/C _18077_/A vssd1 vssd1 vccd1 vccd1 _18078_/Y sky130_fd_sc_hd__a21oi_2
Xhold237 hold237/A vssd1 vssd1 vccd1 vccd1 hold237/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold248 hold248/A vssd1 vssd1 vccd1 vccd1 hold248/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold259 hold259/A vssd1 vssd1 vccd1 vccd1 hold259/X sky130_fd_sc_hd__dlygate4sd3_1
X_17029_ _17029_/A _17029_/B _17146_/C _17146_/D vssd1 vssd1 vccd1 vccd1 _17030_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_40_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1110 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19066__A2 _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20040_ _20041_/A _20041_/B vssd1 vssd1 vccd1 vccd1 _20222_/B sky130_fd_sc_hd__nor2_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11361__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13925__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout180_A _21826_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21991_ _22020_/CLK _21991_/D vssd1 vssd1 vccd1 vccd1 hold199/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout278_A _21799_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20942_ _21054_/A vssd1 vssd1 vccd1 vccd1 _20944_/D sky130_fd_sc_hd__inv_2
XANTENNA__16588__B1 _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12861__A2 _12402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20873_ _20737_/Y _20739_/Y _20870_/Y _20872_/X vssd1 vssd1 vccd1 vccd1 _20873_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__19331__B _19650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout445_A _12785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20687__A2 _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14366__A2 _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15563__A1 _15381_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17786__B _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21425_ hold222/X sstream_i[2] _21442_/S vssd1 vssd1 vccd1 vccd1 _21952_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19059__A _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17304__A2 _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21356_ _21720_/D _18101_/X _21403_/S _21355_/Y vssd1 vssd1 vccd1 vccd1 _21356_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13326__B1 _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20307_ _20307_/A _20307_/B vssd1 vssd1 vccd1 vccd1 _20352_/A sky130_fd_sc_hd__nand2_1
X_21287_ _21287_/A _21287_/B vssd1 vssd1 vccd1 vccd1 _21299_/A sky130_fd_sc_hd__xor2_1
XANTENNA_fanout93_A _19051_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11040_ mstream_o[115] sstream_i[115] _21721_/D vssd1 vssd1 vccd1 vccd1 _21651_/D
+ sky130_fd_sc_hd__mux2_1
X_20238_ _20239_/B vssd1 vssd1 vccd1 vccd1 _20238_/Y sky130_fd_sc_hd__inv_2
XANTENNA__17307__A _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20169_ _20590_/D _20838_/C _20838_/D _20462_/D vssd1 vssd1 vccd1 vccd1 _20173_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13554__B _13554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12991_ _13858_/A _13858_/B _13269_/C _12991_/D vssd1 vssd1 vccd1 vccd1 _13128_/A
+ sky130_fd_sc_hd__nand4_2
XTAP_3611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12301__A1 _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12301__B2 _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14730_ _14730_/A _14730_/B _14854_/B vssd1 vssd1 vccd1 vccd1 _14732_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_118_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11942_ _11870_/A _11870_/B _11870_/C vssd1 vssd1 vccd1 vccd1 _11942_/X sky130_fd_sc_hd__a21o_1
XTAP_3644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14661_ _16374_/A _14817_/C _14817_/D _16203_/D vssd1 vssd1 vccd1 vccd1 _14666_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_2943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11873_ _11822_/X _11871_/Y _11870_/Y _11870_/A vssd1 vssd1 vccd1 vccd1 _11873_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14666__A _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14054__A1 _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14054__B2 _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16400_ _16400_/A _16400_/B vssd1 vssd1 vccd1 vccd1 _16412_/A sky130_fd_sc_hd__xor2_1
XTAP_2976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13612_ _15217_/A _14212_/D _13613_/C _13613_/D vssd1 vssd1 vccd1 vccd1 _13614_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10824_ hold113/A hold134/A vssd1 vssd1 vccd1 vccd1 _11047_/A sky130_fd_sc_hd__and2_1
XTAP_2998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14592_ _14592_/A _14592_/B vssd1 vssd1 vccd1 vccd1 _14595_/A sky130_fd_sc_hd__xnor2_2
X_17380_ _17381_/C _17380_/B vssd1 vssd1 vccd1 vccd1 _17483_/B sky130_fd_sc_hd__or2_1
XANTENNA__20127__A1 _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20127__B2 _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16331_ _16331_/A _16331_/B vssd1 vssd1 vccd1 vccd1 _16332_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_95_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13543_ _13387_/X _13389_/Y _13540_/Y _13542_/X vssd1 vssd1 vccd1 vccd1 _13669_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_82_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17977__A _21791_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_428 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12186__A _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19895__C _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16262_ _15907_/A _16151_/B _16261_/X vssd1 vssd1 vccd1 vccd1 _16298_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_82_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19050_ _19051_/A _19051_/C _19221_/C _20026_/B vssd1 vssd1 vccd1 vccd1 _19050_/X
+ sky130_fd_sc_hd__a22o_1
X_13474_ _14087_/A _15370_/B _15098_/B _14089_/A vssd1 vssd1 vccd1 vccd1 _13475_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15213_ _15201_/A _15201_/B _15200_/A vssd1 vssd1 vccd1 vccd1 _15354_/A sky130_fd_sc_hd__a21o_2
X_18001_ _18849_/B _19060_/B _17863_/B _17861_/X vssd1 vssd1 vccd1 vccd1 _18002_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_51_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12425_ _12510_/B _12425_/B vssd1 vssd1 vccd1 vccd1 _12435_/A sky130_fd_sc_hd__nor2_1
X_16193_ _16193_/A _16193_/B _16193_/C vssd1 vssd1 vccd1 vccd1 _16347_/A sky130_fd_sc_hd__and3_1
XFILLER_0_51_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15320__A2_N _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15144_ _15041_/Y _15043_/X _15298_/A _15143_/X vssd1 vssd1 vccd1 vccd1 _15298_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_50_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12356_ _13155_/A _12784_/A vssd1 vssd1 vccd1 vccd1 _12359_/A sky130_fd_sc_hd__and2_1
XFILLER_0_65_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11307_ fanout58/X v0z[20] fanout17/X _11306_/X vssd1 vssd1 vccd1 vccd1 _11307_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15075_ _15075_/A _15075_/B vssd1 vssd1 vccd1 vccd1 _15082_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19952_ _19951_/A _19951_/B _20247_/D vssd1 vssd1 vccd1 vccd1 _19955_/D sky130_fd_sc_hd__o21a_1
XFILLER_0_77_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12287_ _12294_/C _12294_/D _12287_/C vssd1 vssd1 vccd1 vccd1 _12288_/C sky130_fd_sc_hd__and3b_1
XFILLER_0_121_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14026_ _14027_/A _14663_/D _14027_/C _14027_/D vssd1 vssd1 vccd1 vccd1 _14026_/X
+ sky130_fd_sc_hd__and4_1
X_18903_ _18899_/X _18901_/Y _18737_/X _18740_/X vssd1 vssd1 vccd1 vccd1 _18904_/B
+ sky130_fd_sc_hd__a211o_1
X_11238_ _21718_/D t1x[3] v2z[3] _11459_/B2 _11237_/X vssd1 vssd1 vccd1 vccd1 _11238_/X
+ sky130_fd_sc_hd__a221o_2
X_19883_ _19885_/A _19885_/B _19885_/C _19885_/D vssd1 vssd1 vccd1 vccd1 _19883_/Y
+ sky130_fd_sc_hd__o22ai_1
XANTENNA__13745__A _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18834_ _18834_/A _18834_/B vssd1 vssd1 vccd1 vccd1 _18837_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__16759__C _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11169_ hold266/X fanout51/X fanout49/X hold304/A vssd1 vssd1 vccd1 vccd1 _11169_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16282__A2 _16284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_clk_i_A _21806_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18765_ _18644_/A _18643_/B _18641_/X vssd1 vssd1 vccd1 vccd1 _18780_/A sky130_fd_sc_hd__a21o_1
X_15977_ _16196_/A _15978_/B _15975_/Y _16101_/A vssd1 vssd1 vccd1 vccd1 _15979_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17716_ _17607_/A _17715_/A _17617_/B _17850_/A _17715_/Y vssd1 vssd1 vccd1 vccd1
+ _17718_/C sky130_fd_sc_hd__o32ai_4
XANTENNA__19432__A _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14928_ _15153_/B _15155_/C _15829_/C _15954_/D vssd1 vssd1 vccd1 vccd1 _14930_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18696_ _19185_/D _19008_/D _19013_/C _19179_/C vssd1 vssd1 vccd1 vccd1 _18853_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__19220__A2 _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17647_ _17648_/A _17648_/B vssd1 vssd1 vccd1 vccd1 _17647_/X sky130_fd_sc_hd__and2_1
X_14859_ _14859_/A _15368_/D _14859_/C _14976_/A vssd1 vssd1 vccd1 vccd1 _14976_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_72_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15793__A1 _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17578_ _17575_/X _17576_/Y _17466_/C _17465_/Y vssd1 vssd1 vccd1 vccd1 _17580_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_9_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19317_ _19317_/A _19317_/B vssd1 vssd1 vccd1 vccd1 _19318_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_45_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16529_ _17300_/C _17520_/D _17504_/C _17490_/A vssd1 vssd1 vccd1 vccd1 _16530_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_58_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11204__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_940 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18731__A1 _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18731__B2 _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19248_ _19248_/A _19248_/B _19248_/C vssd1 vssd1 vccd1 vccd1 _19248_/X sky130_fd_sc_hd__and3_1
XFILLER_0_143_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12246__D _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19179_ _19650_/D _19493_/D _19179_/C vssd1 vssd1 vccd1 vccd1 _19179_/X sky130_fd_sc_hd__and3_1
XFILLER_0_131_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15838__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16204__A1_N _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11031__A1 hold270/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21210_ _21305_/A _21283_/B _21305_/B _21311_/A vssd1 vssd1 vccd1 vccd1 _21212_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_143_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11582__A2 _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21141_ _21141_/A _21247_/B vssd1 vssd1 vccd1 vccd1 _21415_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15854__B _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21072_ _20952_/B _20953_/Y _21228_/A _21071_/X vssd1 vssd1 vccd1 vccd1 _21228_/B
+ sky130_fd_sc_hd__a211oi_2
Xfanout503 _21743_/Q vssd1 vssd1 vccd1 vccd1 _13173_/C sky130_fd_sc_hd__buf_4
Xfanout514 _21741_/Q vssd1 vssd1 vccd1 vccd1 _15695_/A sky130_fd_sc_hd__buf_4
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout525 _14027_/A vssd1 vssd1 vccd1 vccd1 _12444_/B sky130_fd_sc_hd__buf_4
Xfanout536 _13867_/A vssd1 vssd1 vccd1 vccd1 _12642_/A sky130_fd_sc_hd__buf_4
XANTENNA_fanout395_A _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12531__A1 _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout547 _21734_/Q vssd1 vssd1 vccd1 vccd1 _15159_/D sky130_fd_sc_hd__clkbuf_8
X_20023_ _20164_/B _20021_/Y _19887_/Y _19925_/A vssd1 vssd1 vccd1 vccd1 _20024_/B
+ sky130_fd_sc_hd__o211ai_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16031__A _16031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout558 _21731_/Q vssd1 vssd1 vccd1 vccd1 _13556_/A sky130_fd_sc_hd__clkbuf_8
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout569 _12403_/B vssd1 vssd1 vccd1 vccd1 _14312_/D sky130_fd_sc_hd__clkbuf_4
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout562_A _14463_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21974_ _21974_/CLK _21974_/D vssd1 vssd1 vccd1 vccd1 hold296/A sky130_fd_sc_hd__dfxtp_1
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20925_ _20925_/A _21097_/B vssd1 vssd1 vccd1 vccd1 _20936_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_90_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14036__A1 _21741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20856_ _20856_/A _20856_/B vssd1 vssd1 vccd1 vccd1 _20877_/A sky130_fd_sc_hd__nand2_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20787_ _21034_/A _20787_/B vssd1 vssd1 vccd1 vccd1 _20788_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11270__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11270__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19278__A2 _19751_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_106_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12210_ _12207_/B _12207_/C _12207_/A vssd1 vssd1 vccd1 vccd1 _12210_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11022__A1 hold234/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21408_ hold124/X _21407_/X _21421_/S vssd1 vssd1 vccd1 vccd1 _21944_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_115_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13190_ _13051_/A _13051_/C _13051_/B vssd1 vssd1 vccd1 vccd1 _13191_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_33_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12770__A1 _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12141_ _12141_/A _12141_/B _12141_/C vssd1 vssd1 vccd1 vccd1 _12148_/A sky130_fd_sc_hd__nand3_1
X_21339_ hold193/X _21421_/S _21337_/Y _21338_/Y vssd1 vssd1 vccd1 vccd1 _21920_/D
+ sky130_fd_sc_hd__o22a_1
XANTENNA__12770__B2 _12771_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12072_ _12080_/A _12073_/A vssd1 vssd1 vccd1 vccd1 _12083_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_124_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20045__B1 _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15900_ _16031_/A _15901_/B vssd1 vssd1 vccd1 vccd1 _15902_/A sky130_fd_sc_hd__nand2_1
X_11023_ mstream_o[97] hold258/X _11027_/S vssd1 vssd1 vccd1 vccd1 hold259/A sky130_fd_sc_hd__mux2_1
X_16880_ _16881_/A _16881_/B vssd1 vssd1 vccd1 vccd1 _16880_/X sky130_fd_sc_hd__and2_1
XFILLER_0_95_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15831_ _15961_/D _16404_/B _15832_/C _15832_/D vssd1 vssd1 vccd1 vccd1 _15833_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_21_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15780__A _16036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18550_ _18550_/A _18550_/B vssd1 vssd1 vccd1 vccd1 _18551_/B sky130_fd_sc_hd__and2_1
X_15762_ _15763_/A _15763_/B vssd1 vssd1 vccd1 vccd1 _16034_/A sky130_fd_sc_hd__and2_2
XTAP_3430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12974_ _13102_/A vssd1 vssd1 vccd1 vccd1 _12976_/C sky130_fd_sc_hd__inv_2
XTAP_3441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_475 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17501_ _17490_/A _17741_/B _17397_/B _17395_/X vssd1 vssd1 vccd1 vccd1 _17510_/A
+ sky130_fd_sc_hd__a31o_1
Xclkbuf_2_1__f_clk_i clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 _21806_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14713_ _14713_/A _14713_/B _16173_/B vssd1 vssd1 vccd1 vccd1 _14848_/B sky130_fd_sc_hd__nand3_2
XTAP_3474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18481_ _18481_/A _18481_/B vssd1 vssd1 vccd1 vccd1 _18491_/A sky130_fd_sc_hd__nor2_1
X_11925_ _11924_/B _11924_/C _11924_/A vssd1 vssd1 vccd1 vccd1 _11928_/B sky130_fd_sc_hd__a21bo_1
XTAP_3485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15693_ _15605_/B _15693_/B vssd1 vssd1 vccd1 vccd1 _15737_/A sky130_fd_sc_hd__nand2b_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_1_clk_i _21822_/CLK vssd1 vssd1 vccd1 vccd1 _21974_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_3496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17764__A2 _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17432_ _17336_/A _17335_/A _17335_/B vssd1 vssd1 vccd1 vccd1 _17439_/A sky130_fd_sc_hd__o21ba_1
X_14644_ _14482_/B _14484_/B _14800_/A _14643_/Y vssd1 vssd1 vccd1 vccd1 _14800_/B
+ sky130_fd_sc_hd__a211oi_1
X_11856_ _11816_/A _11816_/B _11816_/C vssd1 vssd1 vccd1 vccd1 _11857_/C sky130_fd_sc_hd__a21o_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17203__C _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10807_ _10807_/A _10807_/B vssd1 vssd1 vccd1 vccd1 _11065_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14575_ _14575_/A _14575_/B vssd1 vssd1 vccd1 vccd1 _14576_/B sky130_fd_sc_hd__xnor2_4
X_17363_ _17363_/A _17363_/B vssd1 vssd1 vccd1 vccd1 _17365_/B sky130_fd_sc_hd__nand2_2
X_11787_ _11787_/A _11787_/B vssd1 vssd1 vccd1 vccd1 _11788_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_131_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20845__B _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19102_ _19101_/B _19101_/C _19101_/A vssd1 vssd1 vccd1 vccd1 _19103_/C sky130_fd_sc_hd__a21o_1
X_16314_ _16374_/A _16314_/B _16406_/B _16314_/D vssd1 vssd1 vccd1 vccd1 _16400_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__11261__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13526_ _13545_/B vssd1 vssd1 vccd1 vccd1 _13676_/A sky130_fd_sc_hd__inv_2
XFILLER_0_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17294_ _17294_/A _17294_/B vssd1 vssd1 vccd1 vccd1 _17297_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19033_ _18894_/D _18895_/B _19031_/Y _19032_/X vssd1 vssd1 vccd1 vccd1 _19035_/B
+ sky130_fd_sc_hd__a211o_1
XANTENNA__20564__C _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16245_ _16352_/A _16243_/Y _16123_/A _16127_/A vssd1 vssd1 vccd1 vccd1 _16245_/X
+ sky130_fd_sc_hd__a211o_1
X_13457_ _15076_/B _14212_/D _14384_/D _15076_/A vssd1 vssd1 vccd1 vccd1 _13461_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12408_ _12408_/A _12408_/B vssd1 vssd1 vccd1 vccd1 _12410_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_88_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16176_ _16176_/A _16176_/B vssd1 vssd1 vccd1 vccd1 _16178_/A sky130_fd_sc_hd__or2_1
XANTENNA__13459__B _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13388_ _13388_/A _13388_/B vssd1 vssd1 vccd1 vccd1 _13390_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_88_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20861__A _20991_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15127_ _15127_/A _15127_/B vssd1 vssd1 vccd1 vccd1 _15135_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12339_ _12416_/A _12338_/C _12338_/A vssd1 vssd1 vccd1 vccd1 _12375_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15058_ _15059_/B _15059_/A vssd1 vssd1 vccd1 vccd1 _15058_/Y sky130_fd_sc_hd__nand2b_1
X_19935_ _19777_/A _19777_/B _19775_/Y vssd1 vssd1 vccd1 vccd1 _19937_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_142_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18050__B _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12513__A1 _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14009_ _13845_/Y _13847_/Y _14007_/Y _14008_/Y vssd1 vssd1 vccd1 vccd1 _14131_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12513__B2 _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19866_ _20101_/A _20101_/B _19866_/C _19866_/D vssd1 vssd1 vccd1 vccd1 _19867_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_128_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18817_ _18817_/A _18817_/B _18815_/X _18816_/Y vssd1 vssd1 vccd1 vccd1 _18817_/X
+ sky130_fd_sc_hd__or4bb_4
X_19797_ _19656_/A _19656_/B _19659_/A vssd1 vssd1 vccd1 vccd1 _19939_/A sky130_fd_sc_hd__a21o_1
XANTENNA__13625__D _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21536__A0 hold283/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18748_ _19686_/A _19068_/C _19238_/C _19686_/B vssd1 vssd1 vccd1 vccd1 _18751_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17204__A1 _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18679_ _18693_/B _18678_/B _18676_/Y _18677_/X vssd1 vssd1 vccd1 vccd1 _18679_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__20101__A _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20710_ _20710_/A _20710_/B vssd1 vssd1 vccd1 vccd1 _20712_/C sky130_fd_sc_hd__and2_1
XFILLER_0_53_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21690_ _22080_/CLK _21690_/D vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_558 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13777__B1 _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20641_ _20903_/B _20641_/B vssd1 vssd1 vccd1 vccd1 _20900_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_18_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout143_A _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20572_ _20572_/A _20707_/A _20572_/C vssd1 vssd1 vccd1 vccd1 _20707_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_117_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout310_A _21793_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout408_A _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20193__D _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13369__B _13369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12752__A1 _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12752__B2 _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21124_ _20964_/A _21014_/A _21232_/B _21123_/X vssd1 vssd1 vccd1 vccd1 _21238_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__19056__B _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout300 _21795_/Q vssd1 vssd1 vccd1 vccd1 _17621_/C sky130_fd_sc_hd__buf_4
XFILLER_0_111_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout311 _18851_/C vssd1 vssd1 vccd1 vccd1 _19185_/D sky130_fd_sc_hd__buf_4
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout322 _18859_/A vssd1 vssd1 vccd1 vccd1 _17146_/D sky130_fd_sc_hd__buf_4
Xfanout333 _21786_/Q vssd1 vssd1 vccd1 vccd1 _16409_/B sky130_fd_sc_hd__buf_4
X_21055_ _20776_/B _20911_/B _20776_/A vssd1 vssd1 vccd1 vccd1 _21172_/A sky130_fd_sc_hd__o21ba_1
Xfanout344 _14477_/C vssd1 vssd1 vccd1 vccd1 _14155_/C sky130_fd_sc_hd__buf_4
Xfanout355 hold326/X vssd1 vssd1 vccd1 vccd1 _13402_/D sky130_fd_sc_hd__clkbuf_8
Xfanout366 _14663_/D vssd1 vssd1 vccd1 vccd1 _14817_/D sky130_fd_sc_hd__buf_4
XANTENNA__12720__C _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20006_ _20003_/Y _20143_/A _20148_/C _21286_/A vssd1 vssd1 vccd1 vccd1 _20143_/B
+ sky130_fd_sc_hd__and4bb_1
Xfanout377 _14828_/B vssd1 vssd1 vccd1 vccd1 _14365_/C sky130_fd_sc_hd__buf_4
XANTENNA__11617__B _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout388 _15768_/A vssd1 vssd1 vccd1 vccd1 _16027_/A sky130_fd_sc_hd__clkbuf_8
Xfanout399 _21770_/Q vssd1 vssd1 vccd1 vccd1 _14993_/A sky130_fd_sc_hd__buf_2
XFILLER_0_119_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21527__A0 hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout56_A _10798_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14928__B _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21957_ _21963_/CLK _21957_/D vssd1 vssd1 vccd1 vccd1 hold260/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11710_ _12899_/B _12637_/A vssd1 vssd1 vccd1 vccd1 _11714_/A sky130_fd_sc_hd__nand2_1
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20908_ hold117/X fanout8/X _20906_/Y _11550_/A _20907_/Y vssd1 vssd1 vccd1 vccd1
+ _20908_/X sky130_fd_sc_hd__a221o_1
XANTENNA__11491__A1 _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12690_ _12686_/X _12688_/Y _12578_/B _12578_/Y vssd1 vssd1 vccd1 vccd1 _12692_/D
+ sky130_fd_sc_hd__o211a_2
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21888_ _21888_/CLK hold135/X vssd1 vssd1 vccd1 vccd1 hold134/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11641_ _11640_/B _11640_/C _11640_/A vssd1 vssd1 vccd1 vccd1 _11643_/B sky130_fd_sc_hd__a21o_1
X_20839_ _20971_/A vssd1 vssd1 vccd1 vccd1 _20841_/D sky130_fd_sc_hd__inv_2
XFILLER_0_37_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13232__A2 _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15509__A1 _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14360_ _14358_/X _14360_/B vssd1 vssd1 vccd1 vccd1 _14361_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_107_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11243__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11572_ _12109_/C _13556_/A _11571_/B _11568_/X vssd1 vssd1 vccd1 vccd1 _11821_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__14980__A2 _21755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14663__B _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13311_ _15076_/A _15076_/B _14386_/B _14384_/C vssd1 vssd1 vccd1 vccd1 _13455_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__18135__B _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14291_ _14291_/A _14291_/B _14291_/C vssd1 vssd1 vccd1 vccd1 _14294_/C sky130_fd_sc_hd__nor3_1
XFILLER_0_150_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21199__D _21853_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16030_ _16031_/A _16031_/B vssd1 vssd1 vccd1 vccd1 _16032_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_150_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13242_ _13242_/A _13242_/B vssd1 vssd1 vccd1 vccd1 _13243_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_609 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15775__A _16031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13173_ _13171_/Y _13308_/A _13173_/C _15217_/A vssd1 vssd1 vccd1 vccd1 _13308_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_21_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12124_ _12124_/A _12124_/B _12124_/C vssd1 vssd1 vccd1 vccd1 _12124_/X sky130_fd_sc_hd__or3_1
XFILLER_0_102_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17981_ _18120_/A _17981_/B vssd1 vssd1 vccd1 vccd1 _17982_/C sky130_fd_sc_hd__nand2_1
XANTENNA__12911__B _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19720_ _19719_/B _19719_/C _19719_/A vssd1 vssd1 vccd1 vccd1 _19721_/B sky130_fd_sc_hd__a21oi_1
X_16932_ _16873_/A _16873_/C _16873_/B vssd1 vssd1 vccd1 vccd1 _16933_/C sky130_fd_sc_hd__a21o_1
X_12055_ _12055_/A _12055_/B vssd1 vssd1 vccd1 vccd1 _12057_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11808__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11006_ mstream_o[80] hold68/X _11012_/S vssd1 vssd1 vccd1 vccd1 _21617_/D sky130_fd_sc_hd__mux2_1
X_19651_ _19653_/A vssd1 vssd1 vccd1 vccd1 _19818_/A sky130_fd_sc_hd__inv_2
X_16863_ _16863_/A _16863_/B _16863_/C vssd1 vssd1 vccd1 vccd1 _16923_/A sky130_fd_sc_hd__nand3_1
X_18602_ _18603_/A _18603_/B vssd1 vssd1 vccd1 vccd1 _18757_/B sky130_fd_sc_hd__nand2_1
X_15814_ _15815_/A _15815_/B _15815_/C vssd1 vssd1 vccd1 vccd1 _15816_/B sky130_fd_sc_hd__a21o_2
X_19582_ _19581_/B _19581_/C _19581_/A vssd1 vssd1 vccd1 vccd1 _19583_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_88_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16794_ _17141_/A _17141_/B _17223_/A _16860_/C vssd1 vssd1 vccd1 vccd1 _16797_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__19187__B2 _17854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18533_ _18534_/A _18687_/A _18534_/C vssd1 vssd1 vccd1 vccd1 _18536_/A sky130_fd_sc_hd__and3_1
X_15745_ _15607_/X _15612_/C _15743_/Y _15744_/X vssd1 vssd1 vccd1 vccd1 _15745_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_3260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13742__B _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12957_ _12957_/A _12957_/B vssd1 vssd1 vccd1 vccd1 _12957_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__12639__A _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11482__A1 _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18464_ _19686_/B _18769_/B _18464_/C _18464_/D vssd1 vssd1 vccd1 vccd1 _18465_/B
+ sky130_fd_sc_hd__nand4_2
X_11908_ _11840_/X _11841_/Y _11905_/A _11905_/Y vssd1 vssd1 vccd1 vccd1 _11909_/B
+ sky130_fd_sc_hd__a211o_1
X_15676_ _15676_/A _15802_/B vssd1 vssd1 vccd1 vccd1 _15678_/B sky130_fd_sc_hd__or2_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_260 hold262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12888_ _12887_/A _12887_/B _12887_/C vssd1 vssd1 vccd1 vccd1 _12889_/C sky130_fd_sc_hd__a21o_1
XANTENNA_271 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_282 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17415_ _17415_/A _17415_/B vssd1 vssd1 vccd1 vccd1 _17425_/A sky130_fd_sc_hd__and2_1
XANTENNA_293 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14627_ _14627_/A _14627_/B vssd1 vssd1 vccd1 vccd1 _14629_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18395_ _18389_/A _18240_/X _18389_/B vssd1 vssd1 vccd1 vccd1 _18395_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_8_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11839_ _11840_/A _11840_/B _11834_/A vssd1 vssd1 vccd1 vccd1 _11839_/Y sky130_fd_sc_hd__nor3b_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11234__A1 _21718_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11234__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17346_ _17345_/B _17345_/C _17345_/A vssd1 vssd1 vccd1 vccd1 _17348_/B sky130_fd_sc_hd__a21o_1
X_14558_ _14859_/A _15370_/B _14559_/C _14724_/A vssd1 vssd1 vccd1 vccd1 _14560_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13509_ _13509_/A _13509_/B vssd1 vssd1 vccd1 vccd1 _13511_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_141_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17277_ _17277_/A _17387_/A _20797_/A _21258_/A vssd1 vssd1 vccd1 vccd1 _17278_/A
+ sky130_fd_sc_hd__and4_1
X_14489_ _14489_/A _14489_/B vssd1 vssd1 vccd1 vccd1 _14491_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_114_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19016_ _19016_/A _19016_/B vssd1 vssd1 vccd1 vccd1 _19019_/A sky130_fd_sc_hd__xnor2_2
X_16228_ _16109_/Y _16111_/Y _16225_/Y _16226_/X vssd1 vssd1 vccd1 vccd1 _16228_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_141_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12734__A1 _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12734__B2 _13554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16159_ _16371_/A _16391_/B _21754_/Q _16380_/A vssd1 vssd1 vccd1 vccd1 _16163_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19662__A2 _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18870__B1 _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19918_ _19917_/B _19917_/C _19917_/A vssd1 vssd1 vccd1 vccd1 _19918_/Y sky130_fd_sc_hd__a21oi_2
X_19849_ _19849_/A _19849_/B vssd1 vssd1 vccd1 vccd1 _19857_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17976__A2 _19030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_1148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19178__A1 _19650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19178__B2 _19493_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21811_ _21816_/CLK _21811_/D vssd1 vssd1 vccd1 vccd1 hold324/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__17124__B _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout260_A _19823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout358_A _16391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11473__A1 _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21742_ _22005_/CLK _21742_/D vssd1 vssd1 vccd1 vccd1 _21742_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_93_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12268__B _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21673_ _21939_/CLK _21673_/D vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout525_A _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17778__C _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21288__A2 _21283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11225__A1 _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20624_ _20621_/Y _20622_/X _20445_/Y _20448_/Y vssd1 vssd1 vccd1 vccd1 _20624_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__11225__B2 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12422__B1 _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19350__A1 _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19350__B2 _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20555_ _20556_/A _20556_/B vssd1 vssd1 vccd1 vccd1 _20742_/B sky130_fd_sc_hd__or2_1
XFILLER_0_104_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19993__C _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17900__A2 _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14175__B1 _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14714__A2 _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13099__B _13394_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20486_ _20486_/A _20486_/B _20486_/C vssd1 vssd1 vccd1 vccd1 _20486_/X sky130_fd_sc_hd__and3_1
XFILLER_0_89_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20799__A1 _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16467__A2 _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14478__A1 _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16203__B _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21107_ _21107_/A _21107_/B vssd1 vssd1 vccd1 vccd1 _21108_/B sky130_fd_sc_hd__or2_1
Xfanout130 _21836_/Q vssd1 vssd1 vccd1 vccd1 _20103_/A sky130_fd_sc_hd__clkbuf_8
X_22087_ _22096_/CLK _22087_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[23] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_121_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout141 _20249_/A vssd1 vssd1 vccd1 vccd1 _17206_/B sky130_fd_sc_hd__buf_4
Xfanout152 _19092_/A vssd1 vssd1 vccd1 vccd1 _18319_/B sky130_fd_sc_hd__buf_4
X_21038_ _21209_/A vssd1 vssd1 vccd1 vccd1 _21040_/D sky130_fd_sc_hd__inv_2
Xfanout163 _17324_/D vssd1 vssd1 vccd1 vccd1 _19732_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout174 _18058_/A vssd1 vssd1 vccd1 vccd1 _19723_/A sky130_fd_sc_hd__buf_4
XFILLER_0_96_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout185 _21825_/Q vssd1 vssd1 vccd1 vccd1 _17666_/A sky130_fd_sc_hd__buf_4
Xfanout196 hold294/A vssd1 vssd1 vccd1 vccd1 _21171_/B sky130_fd_sc_hd__buf_4
X_13860_ _13860_/A _13997_/C vssd1 vssd1 vccd1 vccd1 _13861_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_69_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12811_ _12807_/X _12809_/Y _12697_/C _12697_/Y vssd1 vssd1 vccd1 vccd1 _12813_/C
+ sky130_fd_sc_hd__o211a_1
X_13791_ _13790_/B _13790_/C _13790_/A vssd1 vssd1 vccd1 vccd1 _13791_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_69_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15530_ _16305_/B _15911_/A _15911_/C _16196_/B vssd1 vssd1 vccd1 vccd1 _15533_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11464__A1 _17443_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ _12743_/A _12743_/B _12743_/C vssd1 vssd1 vccd1 vccd1 _12744_/B sky130_fd_sc_hd__a21oi_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12661__B1 _21765_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18392__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15461_ _15461_/A _15461_/B vssd1 vssd1 vccd1 vccd1 _15464_/C sky130_fd_sc_hd__xnor2_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ _12784_/A _14386_/B vssd1 vssd1 vccd1 vccd1 _12676_/A sky130_fd_sc_hd__and2_1
XFILLER_0_132_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14674__A _16173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18146__A _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17200_ _17619_/B _17621_/C _17300_/C _17520_/D vssd1 vssd1 vccd1 vccd1 _17281_/A
+ sky130_fd_sc_hd__and4_1
X_14412_ _14412_/A _14412_/B vssd1 vssd1 vccd1 vccd1 _14423_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__11216__A1 _11215_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16592__C _16743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11624_ _11833_/A _11833_/B _11833_/C vssd1 vssd1 vccd1 vccd1 _11834_/A sky130_fd_sc_hd__a21oi_1
X_18180_ _18181_/A _18181_/B _18181_/C vssd1 vssd1 vccd1 vccd1 _18183_/B sky130_fd_sc_hd__a21o_2
X_15392_ _16084_/A _15913_/B _15392_/C _15588_/A vssd1 vssd1 vccd1 vccd1 _15588_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_71_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17131_ _17089_/X _17122_/Y _17123_/X _17140_/A vssd1 vssd1 vccd1 vccd1 _17132_/C
+ sky130_fd_sc_hd__a211o_1
X_14343_ _14343_/A _14343_/B vssd1 vssd1 vccd1 vccd1 _14345_/B sky130_fd_sc_hd__xnor2_4
X_11555_ hold2/A _11555_/B vssd1 vssd1 vccd1 vccd1 _12291_/B sky130_fd_sc_hd__or2_4
XFILLER_0_135_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17200__D _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14274_ _14273_/B _14273_/C _14273_/A vssd1 vssd1 vccd1 vccd1 _14274_/Y sky130_fd_sc_hd__a21oi_2
X_17062_ _17016_/A _17016_/C _17016_/B vssd1 vssd1 vccd1 vccd1 _17068_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_40_507 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11486_ _11498_/A1 t1y[12] t0x[12] _11501_/B2 vssd1 vssd1 vccd1 vccd1 _11486_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_122_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16013_ _16015_/A vssd1 vssd1 vccd1 vccd1 _16143_/A sky130_fd_sc_hd__inv_2
X_13225_ fanout9/X _21355_/B vssd1 vssd1 vccd1 vccd1 _13225_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_33_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13156_ _13155_/A _13155_/C _13155_/D _13155_/B vssd1 vssd1 vccd1 vccd1 _13157_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12107_ _12229_/A _12155_/B _12246_/D _12269_/C vssd1 vssd1 vccd1 vccd1 _12110_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_97_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ _13085_/A _13085_/B _12961_/A _12961_/B vssd1 vssd1 vccd1 vccd1 _13087_/X
+ sky130_fd_sc_hd__o211a_1
X_17964_ _17964_/A _17964_/B vssd1 vssd1 vccd1 vccd1 _17966_/B sky130_fd_sc_hd__or2_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19705__A _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19703_ _19906_/A _20146_/B _19703_/C _19906_/C vssd1 vssd1 vccd1 vccd1 _19903_/A
+ sky130_fd_sc_hd__nand4_2
X_16915_ _16909_/A _16908_/C _16908_/B vssd1 vssd1 vccd1 vccd1 _16916_/B sky130_fd_sc_hd__a21o_1
X_12038_ _12268_/A _12530_/A vssd1 vssd1 vccd1 vccd1 _12040_/B sky130_fd_sc_hd__and2_1
X_17895_ _18030_/B _18767_/B _18616_/D _19664_/B vssd1 vssd1 vccd1 vccd1 _17895_/X
+ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_34_clk_i clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _22080_/CLK sky130_fd_sc_hd__clkbuf_16
X_19634_ _19634_/A _19634_/B vssd1 vssd1 vccd1 vccd1 _19787_/B sky130_fd_sc_hd__xnor2_2
X_16846_ _16826_/Y _16844_/X _16845_/Y _16776_/X vssd1 vssd1 vccd1 vccd1 _16851_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_79_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13472__B _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19565_ _20101_/B _19906_/D _19868_/B _20101_/A vssd1 vssd1 vccd1 vccd1 _19565_/X
+ sky130_fd_sc_hd__a22o_1
X_16777_ _16712_/B _16712_/C _16712_/D _16715_/B vssd1 vssd1 vccd1 vccd1 _16777_/X
+ sky130_fd_sc_hd__a22o_1
X_13989_ _13989_/A _13989_/B vssd1 vssd1 vccd1 vccd1 _13990_/B sky130_fd_sc_hd__or2_1
XFILLER_0_88_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18907__A1 _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18516_ _18516_/A _18516_/B _18516_/C _18516_/D vssd1 vssd1 vccd1 vccd1 _18516_/X
+ sky130_fd_sc_hd__or4_1
XANTENNA__18907__B2 _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15728_ _15595_/Y _15597_/Y _15725_/Y _15727_/X vssd1 vssd1 vccd1 vccd1 _15728_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11455__A1 _17557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19496_ _19496_/A _19496_/B vssd1 vssd1 vccd1 vccd1 _19497_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_87_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20586__A _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1094 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18447_ _18314_/D _18316_/A _18445_/X _18594_/B vssd1 vssd1 vccd1 vccd1 _18606_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_29_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15659_ _15796_/A vssd1 vssd1 vccd1 vccd1 _15661_/D sky130_fd_sc_hd__inv_2
XFILLER_0_150_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1078 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20190__A2 _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12404__B1 _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18378_ _18398_/B _18378_/B _18377_/C _18377_/D vssd1 vssd1 vccd1 vccd1 _18378_/X
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19332__A1 _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_28_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17329_ _17329_/A _17329_/B vssd1 vssd1 vccd1 vccd1 _17331_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_43_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16146__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16146__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_356 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20340_ _20340_/A _20340_/B vssd1 vssd1 vccd1 vccd1 _20343_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20271_ _20421_/A vssd1 vssd1 vccd1 vccd1 _20273_/D sky130_fd_sc_hd__inv_2
XFILLER_0_109_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout106_A _21841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22010_ _22013_/CLK _22010_/D vssd1 vssd1 vccd1 vccd1 hold181/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_59_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17646__A1 _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18843__B1 _13967_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12551__B _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout475_A _15093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16621__A2 _17334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13435__A2 _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout642_A _21329_/B1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19988__C _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18892__C _19060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20927__C _21816_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21725_ _21938_/CLK _21725_/D _21329_/B1 vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__dfrtp_4
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14494__A _14494_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21656_ _21934_/CLK _21656_/D vssd1 vssd1 vccd1 vccd1 hold86/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_75_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout19_A _11224_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19323__B2 _19636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11630__B _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20607_ _21087_/D _21311_/B _20605_/Y _20729_/A vssd1 vssd1 vccd1 vccd1 _20609_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_151_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21587_ _21888_/CLK _21587_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[50] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_151_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11340_ _15954_/D _11339_/X _11348_/S vssd1 vssd1 vccd1 vccd1 _21786_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_90_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20538_ _20539_/A _20539_/B vssd1 vssd1 vccd1 vccd1 _20540_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19509__B _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11271_ fanout58/X v0z[11] fanout17/X _11270_/X vssd1 vssd1 vccd1 vccd1 _11271_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_120_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20469_ _20470_/A _20470_/B vssd1 vssd1 vccd1 vccd1 _20471_/A sky130_fd_sc_hd__nor2_1
X_13010_ _13010_/A _13010_/B vssd1 vssd1 vccd1 vccd1 _13029_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17029__B _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12180__C _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16868__B _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14961_ _14795_/X _14797_/Y _14959_/X _14960_/Y vssd1 vssd1 vccd1 vccd1 _14964_/A
+ sky130_fd_sc_hd__o211a_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
X_16700_ _16669_/A _16669_/B _16669_/C vssd1 vssd1 vccd1 vccd1 _16701_/C sky130_fd_sc_hd__a21o_1
X_13912_ _14557_/B _13913_/C _14077_/B _14557_/A vssd1 vssd1 vccd1 vccd1 _13915_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16587__C _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17680_ _17564_/A _17564_/C _17564_/B vssd1 vssd1 vccd1 vccd1 _17681_/C sky130_fd_sc_hd__a21bo_1
X_14892_ _14892_/A _14892_/B vssd1 vssd1 vccd1 vccd1 _14893_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_57_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16612__A2 _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16631_ _16631_/A _16631_/B _16631_/C vssd1 vssd1 vccd1 vccd1 _16634_/B sky130_fd_sc_hd__nand3_4
X_13843_ _13844_/A _13844_/B vssd1 vssd1 vccd1 vccd1 _13843_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__12189__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14623__B2 _14463_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11437__A1 _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19350_ _20026_/B _20733_/C _20606_/D _20178_/D vssd1 vssd1 vccd1 vccd1 _19353_/C
+ sky130_fd_sc_hd__a22o_1
X_16562_ _16989_/C _17520_/B _16561_/C _16586_/A vssd1 vssd1 vccd1 vccd1 _16563_/C
+ sky130_fd_sc_hd__a22o_1
X_13774_ _15370_/B _13773_/X _13772_/X vssd1 vssd1 vccd1 vccd1 _13775_/B sky130_fd_sc_hd__a21bo_1
X_10986_ _10982_/A _10984_/B _10982_/B vssd1 vssd1 vccd1 vccd1 _10988_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_85_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18301_ _18302_/A _18302_/B vssd1 vssd1 vccd1 vccd1 _18453_/B sky130_fd_sc_hd__nand2_1
X_15513_ _15763_/A _16286_/B vssd1 vssd1 vccd1 vccd1 _15517_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19281_ _19432_/A _19753_/B _19281_/C _19427_/A vssd1 vssd1 vccd1 vccd1 _19427_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_69_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12725_ _13822_/B _14018_/C _12725_/C _12725_/D vssd1 vssd1 vccd1 vccd1 _12851_/B
+ sky130_fd_sc_hd__and4_1
X_16493_ _16493_/A _16493_/B _16493_/C vssd1 vssd1 vccd1 vccd1 _16493_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_29_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20172__A2 _20841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18232_ _18091_/B _18091_/Y _18229_/X _18231_/Y vssd1 vssd1 vccd1 vccd1 _18386_/A
+ sky130_fd_sc_hd__a211oi_4
X_15444_ _15311_/A _15449_/A _15310_/B _15306_/X vssd1 vssd1 vccd1 vccd1 _15446_/B
+ sky130_fd_sc_hd__o31ai_2
XFILLER_0_127_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12656_ _12652_/X _12653_/Y _12539_/X _12541_/X vssd1 vssd1 vccd1 vccd1 _12692_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18163_ _18250_/B _18163_/B vssd1 vssd1 vccd1 vccd1 _18225_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11607_ _13012_/B _12312_/A _11606_/C _11606_/D vssd1 vssd1 vccd1 vccd1 _11608_/B
+ sky130_fd_sc_hd__a22oi_1
X_15375_ _15375_/A _16177_/B vssd1 vssd1 vccd1 vccd1 _15376_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_5_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17325__B1 _17324_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12587_ _12604_/B _12587_/B _12585_/Y _12586_/X vssd1 vssd1 vccd1 vccd1 _12587_/X
+ sky130_fd_sc_hd__or4bb_4
XFILLER_0_68_1130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19865__A2 _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17114_ _17114_/A _17114_/B _17114_/C vssd1 vssd1 vccd1 vccd1 _17159_/A sky130_fd_sc_hd__and3_1
XFILLER_0_29_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14326_ _15155_/C _15159_/D _14477_/C _14635_/D vssd1 vssd1 vccd1 vccd1 _14474_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_29_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18094_ _18091_/Y _18092_/X _17956_/Y _17958_/X vssd1 vssd1 vccd1 vccd1 _18095_/C
+ sky130_fd_sc_hd__a211o_1
X_11538_ _11544_/A1 t2x[29] v1z[29] fanout20/X _11537_/X vssd1 vssd1 vccd1 vccd1 _11538_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13748__A _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17045_ _16994_/Y _17010_/X _17028_/Y _17038_/X vssd1 vssd1 vccd1 vccd1 _17046_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14257_ _14095_/A _14095_/C _14095_/B vssd1 vssd1 vccd1 vccd1 _14258_/C sky130_fd_sc_hd__a21bo_1
X_11469_ _11502_/A1 t2x[6] v1z[6] fanout18/X _11468_/X vssd1 vssd1 vccd1 vccd1 _11469_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13208_ _13230_/B _13209_/B _13209_/C _13209_/D vssd1 vssd1 vccd1 vccd1 _13208_/Y
+ sky130_fd_sc_hd__nor4_2
XANTENNA__13467__B _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14188_ _14186_/X _14188_/B vssd1 vssd1 vccd1 vccd1 _14189_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_96_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13139_ _13140_/A _13140_/B _13140_/C vssd1 vssd1 vccd1 vccd1 _13139_/X sky130_fd_sc_hd__and3_1
XFILLER_0_104_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13186__C _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18996_ _18995_/A _18995_/B _18708_/A vssd1 vssd1 vccd1 vccd1 _18999_/C sky130_fd_sc_hd__o21bai_2
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13114__B2 _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17947_ _17948_/A _17948_/B _17948_/C vssd1 vssd1 vccd1 vccd1 _17947_/Y sky130_fd_sc_hd__nor3_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18696__D _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11125__B1 _21422_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_139_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17878_ _17878_/A _17878_/B _17878_/C vssd1 vssd1 vccd1 vccd1 _17881_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16829_ _17041_/A _16899_/B _17141_/C _17493_/A vssd1 vssd1 vccd1 vccd1 _16833_/A
+ sky130_fd_sc_hd__and4_1
X_19617_ _19617_/A _19617_/B vssd1 vssd1 vccd1 vccd1 _19620_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_36_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14614__A1 _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13417__A2 _14516_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11207__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14614__B2 _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11428__A1 _21283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19548_ _21839_/Q _19692_/B _19548_/C _19700_/A vssd1 vssd1 vccd1 vccd1 _19700_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_152_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19479_ hold217/X _19478_/Y fanout4/X vssd1 vssd1 vccd1 vccd1 hold218/A sky130_fd_sc_hd__mux2_1
XFILLER_0_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21510_ hold233/X sstream_i[87] _21510_/S vssd1 vssd1 vccd1 vccd1 _22037_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21441_ hold295/X sstream_i[18] _21442_/S vssd1 vssd1 vccd1 vccd1 _21968_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13050__B1 _14077_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11600__A1 _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21372_ hold47/X fanout40/X _21371_/Y vssd1 vssd1 vccd1 vccd1 _21931_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20323_ _20181_/A _20328_/A _20180_/B _20176_/X vssd1 vssd1 vccd1 vccd1 _20325_/B
+ sky130_fd_sc_hd__o31ai_2
XFILLER_0_141_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14550__B1 _14548_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20254_ _20252_/Y _20254_/B vssd1 vssd1 vccd1 vccd1 _20255_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_40_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16969__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20185_ _20185_/A _20185_/B vssd1 vssd1 vccd1 vccd1 _20206_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11116__A0 _10959_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20926__A1 _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13824__C _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold268_A hold268/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20926__B2 _21267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18595__A2 _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15704__A1_N _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10840_ hold221/A hold80/A _10841_/B vssd1 vssd1 vccd1 vccd1 _10843_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11419__A1 _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14936__B _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19544__A1 _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12510_ _12510_/A _12510_/B vssd1 vssd1 vccd1 vccd1 _12517_/A sky130_fd_sc_hd__or2_1
X_13490_ _13491_/A _13491_/B _13491_/C _13491_/D vssd1 vssd1 vccd1 vccd1 _13490_/Y
+ sky130_fd_sc_hd__nor4_2
X_21708_ _22096_/CLK _21708_/D vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15030__A1 _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12441_ _12877_/B _12899_/B _12345_/B _12343_/X vssd1 vssd1 vccd1 vccd1 _12451_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_137_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21639_ _21722_/CLK _21639_/D fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[102]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_805 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15160_ _15162_/A vssd1 vssd1 vccd1 vccd1 _15315_/A sky130_fd_sc_hd__inv_2
XANTENNA__17858__A1 _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12372_ _11753_/B _11753_/Y _12369_/X _12371_/Y vssd1 vssd1 vccd1 vccd1 _12375_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_117_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14111_ _13948_/C _13947_/Y _14109_/X _14110_/X vssd1 vssd1 vccd1 vccd1 _14111_/Y
+ sky130_fd_sc_hd__o211ai_4
X_11323_ fanout59/X v0z[24] fanout18/X _11322_/X vssd1 vssd1 vccd1 vccd1 _11323_/X
+ sky130_fd_sc_hd__a31o_2
X_15091_ _15892_/A _15632_/B _15091_/C vssd1 vssd1 vccd1 vccd1 _15091_/X sky130_fd_sc_hd__and3_1
XFILLER_0_120_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14042_ _13881_/A _13880_/B _13878_/X vssd1 vssd1 vccd1 vccd1 _14043_/C sky130_fd_sc_hd__a21o_1
XANTENNA__21406__A2 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11254_ _11502_/A1 t1x[7] v2z[7] _11459_/B2 _11253_/X vssd1 vssd1 vccd1 vccd1 _11254_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_120_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18850_ _18851_/C _19179_/C _18848_/Y _19017_/A vssd1 vssd1 vccd1 vccd1 _18854_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_11185_ hold142/X fanout22/X _11184_/X vssd1 vssd1 vccd1 vccd1 _11185_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_140_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15097__A1 _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17801_ _17678_/A _17678_/C _17678_/B vssd1 vssd1 vccd1 vccd1 _17802_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18781_ _18925_/B _18780_/C _18780_/A vssd1 vssd1 vccd1 vccd1 _18781_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__11107__A0 _10892_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15993_ _15991_/B _15991_/C _15991_/A vssd1 vssd1 vccd1 vccd1 _15993_/Y sky130_fd_sc_hd__o21ai_2
X_17732_ _17732_/A _17732_/B vssd1 vssd1 vccd1 vccd1 _17734_/B sky130_fd_sc_hd__or2_2
X_14944_ _14944_/A _14944_/B vssd1 vssd1 vccd1 vccd1 _14967_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17663_ _17661_/X _17663_/B vssd1 vssd1 vccd1 vccd1 _17664_/B sky130_fd_sc_hd__nand2b_1
X_14875_ _15514_/B _16414_/B _16391_/B _15514_/A vssd1 vssd1 vccd1 vccd1 _14878_/C
+ sky130_fd_sc_hd__a22o_1
X_19402_ _19271_/Y _19275_/A _19400_/X _19401_/Y vssd1 vssd1 vccd1 vccd1 _19404_/A
+ sky130_fd_sc_hd__a211oi_1
X_16614_ _16613_/B _16613_/C _16613_/A vssd1 vssd1 vccd1 vccd1 _16615_/C sky130_fd_sc_hd__a21bo_1
X_13826_ _13985_/A _16404_/B _13670_/X _13671_/X _16399_/B vssd1 vssd1 vccd1 vccd1
+ _13828_/B sky130_fd_sc_hd__a32o_1
X_17594_ _17594_/A _17594_/B vssd1 vssd1 vccd1 vccd1 _17595_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_106_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19333_ _19493_/D _20841_/B vssd1 vssd1 vccd1 vccd1 _19334_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13750__B _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16545_ _16547_/A _16547_/B vssd1 vssd1 vccd1 vccd1 _16546_/A sky130_fd_sc_hd__or2_1
XFILLER_0_57_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13757_ _13758_/A _13758_/B _13758_/C vssd1 vssd1 vccd1 vccd1 _13757_/X sky130_fd_sc_hd__o21a_2
XFILLER_0_85_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10969_ hold76/A hold100/A vssd1 vssd1 vccd1 vccd1 _10971_/A sky130_fd_sc_hd__or2_1
XANTENNA__20145__A2 _21305_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16119__A _16119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14565__C _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11551__A _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_971 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19264_ _20650_/A _19906_/D _19264_/C _19264_/D vssd1 vssd1 vccd1 vccd1 _19266_/B
+ sky130_fd_sc_hd__nand4_2
X_12708_ _12708_/A _12708_/B _12825_/B vssd1 vssd1 vccd1 vccd1 _12708_/X sky130_fd_sc_hd__or3_1
XFILLER_0_156_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16476_ _16476_/A _16476_/B vssd1 vssd1 vccd1 vccd1 _16493_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13688_ _13690_/A _13690_/B _13690_/C vssd1 vssd1 vccd1 vccd1 _13689_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_85_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18215_ _18215_/A _18215_/B _18215_/C vssd1 vssd1 vccd1 vccd1 _18215_/Y sky130_fd_sc_hd__nand3_2
X_15427_ _15426_/A _15426_/B _15426_/C _15426_/D vssd1 vssd1 vccd1 vccd1 _15427_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_122_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19195_ _19064_/A _19063_/B _19061_/X vssd1 vssd1 vccd1 vccd1 _19195_/Y sky130_fd_sc_hd__a21oi_1
X_12639_ _12639_/A _13012_/B _12639_/C _12639_/D vssd1 vssd1 vccd1 vccd1 _12641_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_127_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20583__B _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18146_ _19051_/A _20317_/D _19068_/C _19238_/C vssd1 vssd1 vccd1 vccd1 _18293_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__15677__B _15678_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15358_ _12291_/B _15356_/X _15357_/X vssd1 vssd1 vccd1 vccd1 _15358_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold205 hold205/A vssd1 vssd1 vccd1 vccd1 hold205/X sky130_fd_sc_hd__dlygate4sd3_1
X_14309_ _14309_/A _14309_/B vssd1 vssd1 vccd1 vccd1 _14311_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_123_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18077_ _18077_/A _18077_/B _18077_/C vssd1 vssd1 vccd1 vccd1 _18077_/Y sky130_fd_sc_hd__nand3_2
X_15289_ _15290_/A _15290_/B vssd1 vssd1 vccd1 vccd1 _15289_/Y sky130_fd_sc_hd__nand2b_2
Xhold216 hold216/A vssd1 vssd1 vccd1 vccd1 hold216/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold227 hold227/A vssd1 vssd1 vccd1 vccd1 hold227/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 hold238/A vssd1 vssd1 vccd1 vccd1 hold238/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12138__A2 _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17028_ _17028_/A _17028_/B _17028_/C vssd1 vssd1 vccd1 vccd1 _17028_/Y sky130_fd_sc_hd__nand3_1
Xhold249 hold249/A vssd1 vssd1 vccd1 vccd1 hold249/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_1122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13925__B _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18979_ _18979_/A _18979_/B _18979_/C vssd1 vssd1 vccd1 vccd1 _18979_/Y sky130_fd_sc_hd__nor3_2
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12846__B1 _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21990_ _22020_/CLK _21990_/D vssd1 vssd1 vccd1 vccd1 hold183/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__20908__B2 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14621__A_N _14463_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20941_ _21056_/A _21169_/A hold264/A hold294/A vssd1 vssd1 vccd1 vccd1 _21054_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__16588__A1 _21825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16588__B2 _16734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout173_A _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17413__A _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20872_ _20872_/A _20872_/B _20872_/C vssd1 vssd1 vccd1 vccd1 _20872_/X sky130_fd_sc_hd__and3_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19331__C _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15260__A1 _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18445__A2_N _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout340_A _14635_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout438_A _14712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20774__A _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15563__A2 _15386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout605_A _11459_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21424_ hold224/X sstream_i[1] _21442_/S vssd1 vssd1 vccd1 vccd1 _21951_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19059__B _19060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21355_ _21720_/D _21355_/B vssd1 vssd1 vccd1 vccd1 _21355_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_32_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13326__A1 _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18898__B _19230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20306_ _20206_/A _20206_/B _20204_/X vssd1 vssd1 vccd1 vccd1 _20354_/A sky130_fd_sc_hd__o21a_1
XANTENNA__13326__B2 _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21286_ _21286_/A _21286_/B vssd1 vssd1 vccd1 vccd1 _21287_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20237_ _20237_/A _20381_/B vssd1 vssd1 vccd1 vccd1 _20239_/B sky130_fd_sc_hd__xor2_2
XANTENNA_fanout86_A _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17307__B _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20168_ _20168_/A _20168_/B vssd1 vssd1 vccd1 vccd1 _20208_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14826__A1 _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14826__B2 _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13554__C _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12990_ _13858_/A _13012_/B _12878_/X _12877_/X _13152_/C vssd1 vssd1 vccd1 vccd1
+ _12995_/A sky130_fd_sc_hd__a32o_1
X_20099_ _20091_/A _19956_/B _20087_/B _19961_/C vssd1 vssd1 vccd1 vccd1 _20116_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12301__A2 _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11941_ _11941_/A _11941_/B _11941_/C vssd1 vssd1 vccd1 vccd1 _11941_/X sky130_fd_sc_hd__and3_2
XTAP_3645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21572__A1 _11051_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17323__A _17417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14660_ _14660_/A _14660_/B vssd1 vssd1 vccd1 vccd1 _14670_/A sky130_fd_sc_hd__xor2_2
XTAP_2933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11872_ _11870_/A _11870_/Y _11871_/Y _11822_/X vssd1 vssd1 vccd1 vccd1 _11872_/Y
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__14054__A2 _14212_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__22068__RESET_B fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_1059 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13611_ _14557_/A _14557_/B _14218_/B _14873_/B vssd1 vssd1 vccd1 vccd1 _13613_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_95_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10823_ hold74/A hold90/A vssd1 vssd1 vccd1 vccd1 _11050_/B sky130_fd_sc_hd__nor2_1
XTAP_2988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14591_ _14591_/A _14591_/B vssd1 vssd1 vccd1 vccd1 _14592_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__20127__A2 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16330_ _16331_/A _16331_/B vssd1 vssd1 vccd1 vccd1 _16330_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_109_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13542_ _13538_/A _13539_/X _13383_/X _13385_/Y vssd1 vssd1 vccd1 vccd1 _13542_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17977__B _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18585__A1_N _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12186__B _12242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19895__D _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16261_ _16151_/B _16261_/B vssd1 vssd1 vccd1 vccd1 _16261_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_129_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13473_ _14089_/A _14087_/A _15370_/B _15098_/B vssd1 vssd1 vccd1 vccd1 _13475_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_125_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18000_ _17999_/B _17999_/C _17999_/A vssd1 vssd1 vccd1 vccd1 _18002_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_70_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15212_ hold20/X hold39/X fanout4/X vssd1 vssd1 vccd1 vccd1 _21875_/D sky130_fd_sc_hd__mux2_1
XANTENNA__21088__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12424_ _12512_/A _15768_/A _12421_/Y _12423_/B vssd1 vssd1 vccd1 vccd1 _12425_/B
+ sky130_fd_sc_hd__a22oi_1
X_16192_ _16038_/A _16038_/B _16079_/X vssd1 vssd1 vccd1 vccd1 _16193_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_129_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11576__B1 _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15143_ _15253_/B _15141_/X _15006_/X _15012_/C vssd1 vssd1 vccd1 vccd1 _15143_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_125_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12355_ _12355_/A _12355_/B vssd1 vssd1 vccd1 vccd1 _12364_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_121_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16105__C _16396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21632__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11306_ _11224_/A t1x[20] v2z[20] _11223_/A _11305_/X vssd1 vssd1 vccd1 vccd1 _11306_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_61_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15074_ _14968_/A _14965_/X _14966_/Y _14969_/X vssd1 vssd1 vccd1 vccd1 _15196_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11328__A0 _14635_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12286_ _12286_/A _12286_/B _12286_/C vssd1 vssd1 vccd1 vccd1 _12287_/C sky130_fd_sc_hd__or3_1
X_19951_ _19951_/A _19951_/B _20247_/D vssd1 vssd1 vccd1 vccd1 _20087_/A sky130_fd_sc_hd__nand3_2
X_14025_ _14659_/A _14817_/D _14027_/C _14027_/D vssd1 vssd1 vccd1 vccd1 _14025_/X
+ sky130_fd_sc_hd__a22o_1
X_11237_ _11122_/A t2y[3] t0y[3] _11123_/A vssd1 vssd1 vccd1 vccd1 _11237_/X sky130_fd_sc_hd__a22o_1
X_18902_ _18737_/X _18740_/X _18899_/X _18901_/Y vssd1 vssd1 vccd1 vccd1 _18902_/X
+ sky130_fd_sc_hd__o211a_1
X_19882_ _19879_/X _19880_/Y _19756_/B _19758_/B vssd1 vssd1 vccd1 vccd1 _19885_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_120_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11343__A3 fanout20/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13745__B _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18833_ _18834_/A _18833_/B _18833_/C vssd1 vssd1 vccd1 vccd1 _18999_/A sky130_fd_sc_hd__or3_1
X_11168_ _13017_/A _11167_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21739_/D sky130_fd_sc_hd__mux2_1
XANTENNA__16759__D _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11546__A _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18764_ _18760_/Y _18761_/X _18604_/Y _18607_/X vssd1 vssd1 vccd1 vccd1 _18822_/B
+ sky130_fd_sc_hd__a211oi_2
X_15976_ _16196_/B _16305_/B _16396_/B _15976_/D vssd1 vssd1 vccd1 vccd1 _16101_/A
+ sky130_fd_sc_hd__and4_1
X_11099_ _11063_/X hold173/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21693_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_136_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17715_ _17715_/A _17715_/B vssd1 vssd1 vccd1 vccd1 _17715_/Y sky130_fd_sc_hd__nor2_1
X_14927_ _15153_/B _15829_/C _15954_/D _15155_/C vssd1 vssd1 vccd1 vccd1 _14930_/C
+ sky130_fd_sc_hd__a22o_1
X_18695_ _18698_/D vssd1 vssd1 vccd1 vccd1 _18695_/Y sky130_fd_sc_hd__inv_2
XANTENNA__19432__B _19751_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14857__A _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17646_ _17525_/A _18624_/A _17528_/B _17526_/X vssd1 vssd1 vccd1 vccd1 _17648_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_37_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14858_ _14859_/A _15368_/D _14859_/C _14976_/A vssd1 vssd1 vccd1 vccd1 _14860_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19508__A1 _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13809_ _13806_/X _13807_/Y _13548_/Y _13551_/X vssd1 vssd1 vccd1 vccd1 _13809_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_147_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13253__B1 _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17577_ _17466_/C _17465_/Y _17575_/X _17576_/Y vssd1 vssd1 vccd1 vccd1 _17580_/C
+ sky130_fd_sc_hd__o211ai_4
X_14789_ _15153_/B _15978_/B _14790_/C _14946_/A vssd1 vssd1 vccd1 vccd1 _14791_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21315__A1 _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19316_ _19316_/A _19316_/B vssd1 vssd1 vccd1 vccd1 _19317_/B sky130_fd_sc_hd__and2_1
X_16528_ _17300_/C _17504_/C _17490_/A _17520_/D vssd1 vssd1 vccd1 vccd1 _16530_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_46_727 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18731__A2 _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19247_ _19246_/A _19246_/B _19246_/C vssd1 vssd1 vccd1 vccd1 _19248_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_155_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16459_ _17041_/A _17013_/C _17013_/D _16899_/B vssd1 vssd1 vccd1 vccd1 _16459_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19178_ _19650_/D _19013_/C _19179_/C _19493_/D vssd1 vssd1 vccd1 vccd1 _19178_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_147_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18129_ _18129_/A _18129_/B vssd1 vssd1 vccd1 vccd1 _18230_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_42_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21140_ _21138_/A _21026_/B _21138_/B _21025_/B _21137_/Y vssd1 vssd1 vccd1 vccd1
+ _21247_/B sky130_fd_sc_hd__o311a_1
XFILLER_0_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11319__B1 _11318_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18247__A1 _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21071_ _21068_/X _21069_/Y _20913_/Y _20917_/A vssd1 vssd1 vccd1 vccd1 _21071_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout504 _21743_/Q vssd1 vssd1 vccd1 vccd1 _14365_/A sky130_fd_sc_hd__buf_4
XFILLER_0_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout515 _13018_/B vssd1 vssd1 vccd1 vccd1 _13157_/A sky130_fd_sc_hd__buf_4
XANTENNA__16258__B1 _10978_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20022_ _19887_/Y _19925_/A _20164_/B _20021_/Y vssd1 vssd1 vccd1 vccd1 _20024_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__12531__A2 _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout526 _14027_/A vssd1 vssd1 vccd1 vccd1 _13013_/A sky130_fd_sc_hd__clkbuf_2
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout537 _15439_/D vssd1 vssd1 vccd1 vccd1 _13867_/A sky130_fd_sc_hd__buf_4
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout548 _12639_/A vssd1 vssd1 vccd1 vccd1 _12528_/B sky130_fd_sc_hd__buf_4
Xfanout559 _14621_/D vssd1 vssd1 vccd1 vccd1 _14138_/A sky130_fd_sc_hd__buf_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20005__A1_N _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout290_A _17874_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout388_A _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19747__A1 _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11786__A2_N _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21973_ _22016_/CLK _21973_/D vssd1 vssd1 vccd1 vccd1 hold291/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout555_A _14774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13671__A _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20924_ _20924_/A _21264_/A _20924_/C _21097_/A vssd1 vssd1 vccd1 vccd1 _21097_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_96_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15233__A1 _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14036__A2 _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15233__B2 _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20855_ _20855_/A _20855_/B vssd1 vssd1 vccd1 vccd1 _20856_/B sky130_fd_sc_hd__or2_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14992__B1 _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20786_ _20786_/A _20786_/B vssd1 vssd1 vccd1 vccd1 _20787_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_996 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21407_ _15888_/Y _20769_/Y _21407_/S vssd1 vssd1 vccd1 vccd1 _21407_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_150_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12140_ _12139_/B _12139_/C _12139_/A vssd1 vssd1 vccd1 vccd1 _12141_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_60_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21338_ _21407_/S _12493_/B _21421_/S vssd1 vssd1 vccd1 vccd1 _21338_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__12770__A2 _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12071_ _12071_/A _12071_/B vssd1 vssd1 vccd1 vccd1 _12080_/A sky130_fd_sc_hd__or2_1
XFILLER_0_102_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21269_ _21269_/A _21269_/B vssd1 vssd1 vccd1 vccd1 _21271_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12750__A _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20045__A1 _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11022_ mstream_o[96] hold234/X _11027_/S vssd1 vssd1 vccd1 vccd1 _21633_/D sky130_fd_sc_hd__mux2_1
XANTENNA__20045__B2 _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15830_ _15959_/A vssd1 vssd1 vccd1 vccd1 _15832_/D sky130_fd_sc_hd__inv_2
XTAP_3420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15761_ hold78/X _15760_/X fanout2/X vssd1 vssd1 vccd1 vccd1 _21879_/D sky130_fd_sc_hd__mux2_1
X_12973_ _14312_/D _13822_/B _14176_/C _13402_/D vssd1 vssd1 vccd1 vccd1 _13102_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17500_ _17500_/A _17500_/B vssd1 vssd1 vccd1 vccd1 _17513_/A sky130_fd_sc_hd__xnor2_1
XTAP_3453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14712_ _14712_/A _14712_/B _16173_/B vssd1 vssd1 vccd1 vccd1 _14712_/X sky130_fd_sc_hd__and3_1
XTAP_3464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18480_ _18477_/Y _18478_/X _18323_/X _18325_/X vssd1 vssd1 vccd1 vccd1 _18516_/B
+ sky130_fd_sc_hd__a211oi_2
X_11924_ _11924_/A _11924_/B _11924_/C vssd1 vssd1 vccd1 vccd1 _11999_/A sky130_fd_sc_hd__nand3_1
X_15692_ _15689_/Y _15690_/X _15528_/Y _15567_/X vssd1 vssd1 vccd1 vccd1 _15741_/B
+ sky130_fd_sc_hd__o211a_1
XTAP_3475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17431_ _17417_/A _19432_/A _17326_/B _17324_/X vssd1 vssd1 vccd1 vccd1 _17441_/A
+ sky130_fd_sc_hd__a31o_1
X_14643_ _14642_/B _14642_/C _14631_/Y vssd1 vssd1 vccd1 vccd1 _14643_/Y sky130_fd_sc_hd__a21boi_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ _11854_/B _11854_/C _11854_/A vssd1 vssd1 vccd1 vccd1 _11857_/B sky130_fd_sc_hd__a21bo_1
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17203__D _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10806_ hold88/A hold34/A vssd1 vssd1 vccd1 vccd1 _10807_/B sky130_fd_sc_hd__or2_1
X_17362_ _17362_/A _17362_/B vssd1 vssd1 vccd1 vccd1 _17365_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14574_ _14575_/B _14575_/A vssd1 vssd1 vccd1 vccd1 _14574_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_67_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11786_ _12223_/A _12751_/B _11625_/X _11626_/Y vssd1 vssd1 vccd1 vccd1 _11787_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_144_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19101_ _19101_/A _19101_/B _19101_/C vssd1 vssd1 vccd1 vccd1 _19103_/B sky130_fd_sc_hd__nand3_2
X_16313_ _16374_/A _16406_/B _16314_/D _16314_/B vssd1 vssd1 vccd1 vccd1 _16315_/A
+ sky130_fd_sc_hd__a22o_1
X_13525_ _13525_/A _13985_/A _16399_/B _16409_/B vssd1 vssd1 vccd1 vccd1 _13545_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__20845__C _21853_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17293_ _17293_/A _17293_/B vssd1 vssd1 vccd1 vccd1 _17294_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19032_ _19650_/D _19201_/B _19032_/C _19032_/D vssd1 vssd1 vccd1 vccd1 _19032_/X
+ sky130_fd_sc_hd__and4_1
X_16244_ _16123_/A _16127_/A _16352_/A _16243_/Y vssd1 vssd1 vccd1 vccd1 _16352_/B
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_153_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13456_ _14716_/A _14384_/D _13322_/B _13320_/X vssd1 vssd1 vccd1 vccd1 _13464_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_955 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12407_ _12408_/A _12408_/B vssd1 vssd1 vccd1 vccd1 _12521_/A sky130_fd_sc_hd__nand2_1
X_16175_ _16284_/A _16286_/B _16284_/B vssd1 vssd1 vccd1 vccd1 _16176_/B sky130_fd_sc_hd__and3_1
XANTENNA__13459__C _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13387_ _13388_/A _13388_/B vssd1 vssd1 vccd1 vccd1 _13387_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_437 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11040__S _21721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20861__B _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15126_ _15126_/A _15126_/B vssd1 vssd1 vccd1 vccd1 _15140_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_10_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12338_ _12338_/A _12416_/A _12338_/C vssd1 vssd1 vccd1 vccd1 _12416_/B sky130_fd_sc_hd__nand3_1
X_15057_ _14897_/A _14897_/B _14895_/Y vssd1 vssd1 vccd1 vccd1 _15059_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19934_ _19934_/A _19934_/B vssd1 vssd1 vccd1 vccd1 _19937_/A sky130_fd_sc_hd__xnor2_1
X_12269_ _12269_/A _12269_/B _12269_/C _12269_/D vssd1 vssd1 vccd1 vccd1 _12269_/X
+ sky130_fd_sc_hd__and4_1
XANTENNA__12660__A _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14008_ _14004_/X _14005_/Y _13842_/A _13843_/Y vssd1 vssd1 vccd1 vccd1 _14008_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__18050__C _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12513__A2 _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19865_ _20101_/B _21153_/B _19866_/D _20101_/A vssd1 vssd1 vccd1 vccd1 _19867_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18816_ _18812_/X _18814_/Y _18664_/B _18664_/Y vssd1 vssd1 vccd1 vccd1 _18816_/Y
+ sky130_fd_sc_hd__o211ai_2
X_19796_ _19796_/A _19796_/B vssd1 vssd1 vccd1 vccd1 _19944_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_128_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15959_ _15959_/A _15959_/B vssd1 vssd1 vccd1 vccd1 _15960_/B sky130_fd_sc_hd__nor2_2
X_18747_ _19686_/A _18769_/B _18618_/A _18617_/A vssd1 vssd1 vccd1 vccd1 _18752_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__13474__B1 _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17204__A2 _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18678_ _18693_/B _18678_/B _18676_/Y _18677_/X vssd1 vssd1 vccd1 vccd1 _18678_/X
+ sky130_fd_sc_hd__or4bb_2
XFILLER_0_77_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13922__C _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20101__B _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13226__B1 _11061_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17629_ _17629_/A _17629_/B _17629_/C vssd1 vssd1 vccd1 vccd1 _17630_/C sky130_fd_sc_hd__and3_1
XANTENNA__17898__A _19823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13777__A1 _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20640_ _20903_/B _20641_/B vssd1 vssd1 vccd1 vccd1 _20640_/X sky130_fd_sc_hd__and2b_1
XANTENNA__13777__B2 _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18165__B1 _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21213__A _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20571_ _20571_/A _20571_/B _20571_/C vssd1 vssd1 vccd1 vccd1 _20572_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_116_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout136_A _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14726__B1 _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout303_A _17086_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_1014 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12752__A2 _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19337__B _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21123_ _21232_/A _21122_/B _21236_/B _21122_/D vssd1 vssd1 vccd1 vccd1 _21123_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_1058 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19056__C _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout301 _21795_/Q vssd1 vssd1 vccd1 vccd1 _18849_/A sky130_fd_sc_hd__clkbuf_8
Xfanout312 _21793_/Q vssd1 vssd1 vccd1 vccd1 _18851_/C sky130_fd_sc_hd__buf_4
XANTENNA__19968__A1 _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21054_ _21054_/A _21054_/B vssd1 vssd1 vccd1 vccd1 _21064_/A sky130_fd_sc_hd__or2_1
Xfanout323 _18859_/A vssd1 vssd1 vccd1 vccd1 _17387_/A sky130_fd_sc_hd__buf_4
Xfanout334 _16084_/C vssd1 vssd1 vccd1 vccd1 _15829_/C sky130_fd_sc_hd__buf_4
Xfanout345 _21782_/Q vssd1 vssd1 vccd1 vccd1 _14477_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__11712__B1 _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout356 _14176_/C vssd1 vssd1 vccd1 vccd1 _13858_/C sky130_fd_sc_hd__buf_6
X_20005_ _20148_/C _21286_/A _20003_/Y _20143_/A vssd1 vssd1 vccd1 vccd1 _20007_/B
+ sky130_fd_sc_hd__o2bb2a_1
Xfanout367 _15916_/B vssd1 vssd1 vccd1 vccd1 _14663_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__12720__D _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout378 _16284_/A vssd1 vssd1 vccd1 vccd1 _15931_/B sky130_fd_sc_hd__buf_4
Xfanout389 _21772_/Q vssd1 vssd1 vccd1 vccd1 _15768_/A sky130_fd_sc_hd__buf_6
XANTENNA__11617__C _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14928__C _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21956_ _21963_/CLK _21956_/D vssd1 vssd1 vccd1 vccd1 hold231/A sky130_fd_sc_hd__dfxtp_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20907_ _21142_/A _21409_/B vssd1 vssd1 vccd1 vccd1 _20907_/Y sky130_fd_sc_hd__nor2_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21887_ _22106_/CLK _21887_/D vssd1 vssd1 vccd1 vccd1 hold223/A sky130_fd_sc_hd__dfxtp_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _11640_/A _11640_/B _11640_/C vssd1 vssd1 vccd1 vccd1 _11643_/A sky130_fd_sc_hd__nand3_1
X_20838_ _21199_/A _20838_/B _20838_/C _20838_/D vssd1 vssd1 vccd1 vccd1 _20971_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_126_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15509__A2 _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11571_ _11568_/X _11571_/B vssd1 vssd1 vccd1 vccd1 _11865_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_91_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20769_ _20900_/B _20769_/B vssd1 vssd1 vccd1 vccd1 _20769_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_64_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13310_ _15076_/B _14386_/B _14384_/C _15076_/A vssd1 vssd1 vccd1 vccd1 _13310_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_80_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18135__C _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14290_ _14290_/A _14290_/B vssd1 vssd1 vccd1 vccd1 _14290_/X sky130_fd_sc_hd__or2_1
XFILLER_0_64_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13241_ _13242_/A _13242_/B vssd1 vssd1 vccd1 vccd1 _13241_/X sky130_fd_sc_hd__or2_1
XFILLER_0_21_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18432__A _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20266__A1 _21261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13172_ _15076_/A _15076_/B _14365_/D _14386_/B vssd1 vssd1 vccd1 vccd1 _13308_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_60_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11951__B1 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12123_ _12124_/A _12124_/B _12124_/C vssd1 vssd1 vccd1 vccd1 _12123_/Y sky130_fd_sc_hd__nor3_1
X_17980_ _17980_/A _17980_/B _17980_/C vssd1 vssd1 vccd1 vccd1 _17981_/B sky130_fd_sc_hd__or3_1
XFILLER_0_62_1169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12911__C _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16931_ _16930_/B _16930_/C _16930_/A vssd1 vssd1 vccd1 vccd1 _16933_/B sky130_fd_sc_hd__a21bo_1
X_12054_ _12781_/D _12214_/C _12046_/B _12044_/X vssd1 vssd1 vccd1 vccd1 _12057_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__11808__B _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11005_ mstream_o[79] hold24/X _11005_/S vssd1 vssd1 vccd1 vccd1 _21616_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_74_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16862_ _17141_/A _16860_/C _16917_/C _17141_/B vssd1 vssd1 vccd1 vccd1 _16863_/C
+ sky130_fd_sc_hd__a22o_1
X_19650_ _18849_/A _20178_/B _20721_/C _19650_/D vssd1 vssd1 vccd1 vccd1 _19653_/A
+ sky130_fd_sc_hd__and4b_2
XFILLER_0_102_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_15813_ _15813_/A _15813_/B vssd1 vssd1 vccd1 vccd1 _15815_/C sky130_fd_sc_hd__xnor2_1
X_18601_ _18757_/A _18601_/B vssd1 vssd1 vccd1 vccd1 _18603_/B sky130_fd_sc_hd__and2_1
X_19581_ _19581_/A _19581_/B _19581_/C vssd1 vssd1 vccd1 vccd1 _19583_/B sky130_fd_sc_hd__nand3_1
X_16793_ _16790_/A _16789_/C _16789_/A vssd1 vssd1 vccd1 vccd1 _17165_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_137_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18532_ _18684_/B _18530_/Y _18380_/Y _18382_/Y vssd1 vssd1 vccd1 vccd1 _18534_/C
+ sky130_fd_sc_hd__a211o_1
X_15744_ _15741_/X _15742_/Y _15612_/A _15612_/Y vssd1 vssd1 vccd1 vccd1 _15744_/X
+ sky130_fd_sc_hd__a211o_1
XTAP_3250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13742__C _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12956_ _12824_/A _12824_/B _13091_/A _12950_/B vssd1 vssd1 vccd1 vccd1 _12956_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_133_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12639__B _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18463_ _19686_/B _18769_/B _18464_/C _18464_/D vssd1 vssd1 vccd1 vccd1 _18465_/A
+ sky130_fd_sc_hd__a22o_1
X_11907_ _11907_/A vssd1 vssd1 vccd1 vccd1 _12496_/A sky130_fd_sc_hd__inv_2
X_15675_ _15802_/A _16377_/B _15808_/C _15675_/D vssd1 vssd1 vccd1 vccd1 _15802_/B
+ sky130_fd_sc_hd__and4b_1
XANTENNA__14557__D _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_250 hold262/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12887_ _12887_/A _12887_/B _12887_/C vssd1 vssd1 vccd1 vccd1 _13010_/A sky130_fd_sc_hd__nand3_1
XANTENNA_261 hold262/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_272 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17414_ _17619_/B _17636_/B _17413_/C _17413_/D vssd1 vssd1 vccd1 vccd1 _17415_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14626_ _14467_/A _14466_/A _14466_/B _14462_/B _14462_/A vssd1 vssd1 vccd1 vccd1
+ _14627_/B sky130_fd_sc_hd__o32ai_4
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_283 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18394_ _18394_/A _18394_/B _18394_/C vssd1 vssd1 vccd1 vccd1 _18394_/Y sky130_fd_sc_hd__nor3_2
X_11838_ _11805_/X _11806_/Y _11836_/A _11836_/Y vssd1 vssd1 vccd1 vccd1 _11840_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA_294 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18147__B1 _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17345_ _17345_/A _17345_/B _17345_/C vssd1 vssd1 vccd1 vccd1 _17348_/A sky130_fd_sc_hd__nand3_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14557_ _14557_/A _14557_/B _15510_/B _14557_/D vssd1 vssd1 vccd1 vccd1 _14724_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12431__A1 _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11769_ _11685_/A _11685_/C _11685_/B vssd1 vssd1 vccd1 vccd1 _11770_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13508_ _13508_/A _13508_/B vssd1 vssd1 vccd1 vccd1 _13511_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_130_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17276_ _17277_/A _20797_/A _21258_/A _17387_/A vssd1 vssd1 vccd1 vccd1 _17279_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14488_ _14647_/B _14488_/B vssd1 vssd1 vccd1 vccd1 _14491_/A sky130_fd_sc_hd__nand2b_2
X_19015_ _19185_/D _19181_/B vssd1 vssd1 vccd1 vccd1 _19016_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_71_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16227_ _16109_/Y _16111_/Y _16225_/Y _16226_/X vssd1 vssd1 vccd1 vccd1 _16227_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_114_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13439_ _13439_/A _13439_/B vssd1 vssd1 vccd1 vccd1 _13449_/A sky130_fd_sc_hd__and2_1
XFILLER_0_70_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12734__A2 _13269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16158_ _16158_/A _16324_/B vssd1 vssd1 vccd1 vccd1 _16169_/A sky130_fd_sc_hd__or2_1
XFILLER_0_144_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15109_ _15107_/Y _15250_/B _15012_/B _15011_/Y vssd1 vssd1 vccd1 vccd1 _15147_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_122_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16089_ _16089_/A _16089_/B vssd1 vssd1 vccd1 vccd1 _16091_/B sky130_fd_sc_hd__or2_1
XANTENNA__18870__B2 _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19917_ _19917_/A _19917_/B _19917_/C vssd1 vssd1 vccd1 vccd1 _19917_/X sky130_fd_sc_hd__and3_2
XFILLER_0_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19848_ _19961_/A _20381_/A vssd1 vssd1 vccd1 vccd1 _20237_/A sky130_fd_sc_hd__nor2_2
X_19779_ _19779_/A _19779_/B _19779_/C vssd1 vssd1 vccd1 vccd1 _19780_/B sky130_fd_sc_hd__nand3_1
XANTENNA__19178__A2 _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13998__A1 _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21810_ _21816_/CLK _21810_/D vssd1 vssd1 vccd1 vccd1 hold331/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__17124__C _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21741_ _22021_/CLK _21741_/D vssd1 vssd1 vccd1 vccd1 _21741_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_66_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout253_A _18166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21672_ _21939_/CLK _21672_/D vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17778__D _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12422__A1 _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20623_ _20445_/Y _20448_/Y _20621_/Y _20622_/X vssd1 vssd1 vccd1 vccd1 _20623_/X
+ sky130_fd_sc_hd__a211o_2
XANTENNA_fanout420_A _21765_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12422__B2 _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12565__A _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15579__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout518_A _21740_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19350__A2 _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20554_ _20554_/A _20554_/B vssd1 vssd1 vccd1 vccd1 _20556_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_144_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14175__A1 _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14175__B2 _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20485_ _20486_/A _20486_/B _20486_/C vssd1 vssd1 vccd1 vccd1 _20485_/Y sky130_fd_sc_hd__a21oi_4
XANTENNA__13099__C _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20799__A2 _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_0_clk_i _21822_/CLK vssd1 vssd1 vccd1 vccd1 _21767_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_121_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14478__A2 _15174_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21106_ _21107_/A _21107_/B vssd1 vssd1 vccd1 vccd1 _21222_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16203__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_22086_ _22096_/CLK _22086_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[22] sky130_fd_sc_hd__dfrtp_4
Xfanout120 _20562_/B vssd1 vssd1 vccd1 vccd1 _20146_/B sky130_fd_sc_hd__buf_6
Xfanout131 _20774_/B vssd1 vssd1 vccd1 vccd1 _17520_/D sky130_fd_sc_hd__buf_4
Xfanout142 _21833_/Q vssd1 vssd1 vccd1 vccd1 _20249_/A sky130_fd_sc_hd__clkbuf_4
X_21037_ _21151_/A _21301_/A _21283_/A _21264_/B vssd1 vssd1 vccd1 vccd1 _21209_/A
+ sky130_fd_sc_hd__and4_1
Xfanout153 _19092_/A vssd1 vssd1 vccd1 vccd1 _19972_/A sky130_fd_sc_hd__buf_6
XFILLER_0_121_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout164 _21829_/Q vssd1 vssd1 vccd1 vccd1 _17324_/D sky130_fd_sc_hd__clkbuf_4
XANTENNA__15427__A1 _15426_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout175 _21827_/Q vssd1 vssd1 vccd1 vccd1 _18058_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__16500__A _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout186 _21824_/Q vssd1 vssd1 vccd1 vccd1 _17145_/A sky130_fd_sc_hd__buf_4
XFILLER_0_22_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout197 _21258_/B vssd1 vssd1 vccd1 vccd1 _20249_/B sky130_fd_sc_hd__buf_4
XFILLER_0_96_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12810_ _12697_/C _12697_/Y _12807_/X _12809_/Y vssd1 vssd1 vccd1 vccd1 _12813_/B
+ sky130_fd_sc_hd__a211oi_4
X_13790_ _13790_/A _13790_/B _13790_/C vssd1 vssd1 vccd1 vccd1 _13790_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__14020__A _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_1069 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12741_ _12741_/A _12741_/B vssd1 vssd1 vccd1 vccd1 _12743_/C sky130_fd_sc_hd__xnor2_2
X_21939_ _21939_/CLK _21939_/D vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_97_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12661__A1 _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12661__B2 _13018_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18427__A _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15460_ _15461_/A _15461_/B vssd1 vssd1 vccd1 vccd1 _15460_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14938__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ _12672_/A _12672_/B vssd1 vssd1 vccd1 vccd1 _12681_/A sky130_fd_sc_hd__nor2_1
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14674__B _14828_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14411_ _14409_/X _14411_/B vssd1 vssd1 vccd1 vccd1 _14412_/B sky130_fd_sc_hd__and2b_1
XANTENNA__18146__B _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16592__D _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ _11623_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _11833_/C sky130_fd_sc_hd__xnor2_1
X_15391_ _16084_/A _15913_/B _15392_/C _15588_/A vssd1 vssd1 vccd1 vccd1 _15393_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13610__B1 _14873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17130_ _17130_/A _17130_/B vssd1 vssd1 vccd1 vccd1 _17132_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_37_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14342_ _14343_/B _14343_/A vssd1 vssd1 vccd1 vccd1 _14453_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_108_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11554_ hold2/A _11555_/B vssd1 vssd1 vccd1 vccd1 fanout9/A sky130_fd_sc_hd__nor2_4
XFILLER_0_123_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15786__A _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17061_ _17025_/A _17025_/C _17025_/B vssd1 vssd1 vccd1 vccd1 _17073_/B sky130_fd_sc_hd__a21o_1
X_14273_ _14273_/A _14273_/B _14273_/C vssd1 vssd1 vccd1 vccd1 _14273_/X sky130_fd_sc_hd__and3_1
XFILLER_0_123_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11485_ _11484_/X _18624_/A _11521_/S vssd1 vssd1 vccd1 vccd1 _21833_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_40_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16012_ _16014_/A _16014_/B vssd1 vssd1 vccd1 vccd1 _16015_/A sky130_fd_sc_hd__or2_1
XFILLER_0_21_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13224_ _13224_/A _13518_/B vssd1 vssd1 vccd1 vccd1 _21355_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_33_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_1042 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13155_ _13155_/A _13155_/B _13155_/C _13155_/D vssd1 vssd1 vccd1 vccd1 _13298_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_104_1221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _12106_/A _12106_/B vssd1 vssd1 vccd1 vccd1 _12112_/A sky130_fd_sc_hd__xnor2_1
X_17963_ _17962_/B _17962_/C _17962_/A vssd1 vssd1 vccd1 vccd1 _17964_/B sky130_fd_sc_hd__o21a_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ _12961_/A _12961_/B _13085_/A _13085_/B vssd1 vssd1 vccd1 vccd1 _13223_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_104_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19702_ _20146_/B _19703_/C _19906_/C _19906_/A vssd1 vssd1 vccd1 vccd1 _19705_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16914_ _17372_/A _16914_/B vssd1 vssd1 vccd1 vccd1 _17171_/A sky130_fd_sc_hd__xor2_4
X_12037_ _12261_/A _12269_/B _12637_/B _12639_/A vssd1 vssd1 vccd1 vccd1 _12040_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19801__B1 _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17894_ _18030_/B _19664_/B _18616_/D vssd1 vssd1 vccd1 vccd1 _17894_/X sky130_fd_sc_hd__and3_1
XFILLER_0_109_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21028__A _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19633_ _19634_/A _19634_/B vssd1 vssd1 vccd1 vccd1 _19633_/X sky130_fd_sc_hd__and2b_1
X_16845_ _16756_/Y _16757_/X _16783_/B _16776_/D vssd1 vssd1 vccd1 vccd1 _16845_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
X_16776_ _16756_/Y _16757_/X _16783_/B _16776_/D vssd1 vssd1 vccd1 vccd1 _16776_/X
+ sky130_fd_sc_hd__and4bb_2
X_19564_ _19436_/A _19435_/B _19433_/X vssd1 vssd1 vccd1 vccd1 _19581_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_137_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13988_ _13989_/A _13989_/B vssd1 vssd1 vccd1 vccd1 _14149_/B sky130_fd_sc_hd__nand2_1
XANTENNA__18907__A2 _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15727_ _15727_/A _15727_/B _15727_/C vssd1 vssd1 vccd1 vccd1 _15727_/X sky130_fd_sc_hd__and3_1
XFILLER_0_88_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18515_ _18516_/A _18516_/B _18516_/C _18516_/D vssd1 vssd1 vccd1 vccd1 _18515_/Y
+ sky130_fd_sc_hd__nor4_1
XTAP_3080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12939_ _12938_/B _12938_/C _12938_/A vssd1 vssd1 vccd1 vccd1 _12939_/X sky130_fd_sc_hd__a21o_1
XTAP_3091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19495_ _18849_/A _20178_/B _21261_/B _18849_/B vssd1 vssd1 vccd1 vccd1 _19496_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12088__C _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15658_ _15791_/A _15916_/B _16040_/C _16396_/A vssd1 vssd1 vccd1 vccd1 _15796_/A
+ sky130_fd_sc_hd__and4_1
X_18446_ _18443_/Y _18594_/A _19051_/A _19240_/B vssd1 vssd1 vccd1 vccd1 _18594_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_34_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14609_ _14596_/A _14596_/B _14594_/Y vssd1 vssd1 vccd1 vccd1 _14758_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_146_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18377_ _18398_/B _18378_/B _18377_/C _18377_/D vssd1 vssd1 vccd1 vccd1 _18377_/X
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__12404__A1 _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15589_ _16374_/A _15717_/C _15976_/D _16087_/A vssd1 vssd1 vccd1 vccd1 _15593_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__12404__B2 _12403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17328_ _17329_/A _17329_/B vssd1 vssd1 vccd1 vccd1 _17427_/A sky130_fd_sc_hd__nand2b_2
XFILLER_0_71_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10966__A1 _10965_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17259_ _17256_/X _17257_/Y _16657_/C _16656_/Y vssd1 vssd1 vccd1 vccd1 _17260_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_109_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20270_ _20416_/A _20416_/B _20270_/C _20924_/A vssd1 vssd1 vccd1 vccd1 _20421_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_11_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17646__A2 _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18843__B2 _11550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15657__A1 _15916_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12551__C _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_985 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17416__A _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19652__A1_N _19650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout370_A _12402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout468_A _14698_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20777__A _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18892__D _19051_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout635_A _21776_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21724_ _21724_/CLK _21724_/D _21422_/A vssd1 vssd1 vccd1 vccd1 _21724_/Q sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20927__D _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_1157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21655_ _21888_/CLK _21655_/D vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20606_ _21261_/A _20863_/C _21283_/B _20606_/D vssd1 vssd1 vccd1 vccd1 _20729_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_90_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21586_ _21888_/CLK _21586_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[49] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_7_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20537_ _20918_/A _20404_/B _20788_/A vssd1 vssd1 vccd1 vccd1 _20539_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_104_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ _11502_/A1 t1x[11] v2z[11] _11501_/B2 _11269_/X vssd1 vssd1 vccd1 vccd1 _11270_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20468_ _20468_/A _20468_/B vssd1 vssd1 vccd1 vccd1 _20470_/B sky130_fd_sc_hd__or2_1
XFILLER_0_127_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11639__A _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20399_ _20399_/A _20399_/B vssd1 vssd1 vccd1 vccd1 _20401_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__17029__C _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13123__A2 _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12180__D _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14960_ _14956_/X _14957_/Y _14793_/B _14795_/B vssd1 vssd1 vccd1 vccd1 _14960_/Y
+ sky130_fd_sc_hd__o211ai_2
X_22069_ _22069_/CLK _22069_/D fanout639/X vssd1 vssd1 vccd1 vccd1 mstream_o[5] sky130_fd_sc_hd__dfrtp_4
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
X_13911_ _14848_/A _14077_/B _13772_/X _13773_/X _15370_/B vssd1 vssd1 vccd1 vccd1
+ _13916_/A sky130_fd_sc_hd__a32o_1
XANTENNA__16587__D _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14891_ _14892_/B _14892_/A vssd1 vssd1 vccd1 vccd1 _14891_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_57_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16630_ _16629_/B _16629_/C _16629_/A vssd1 vssd1 vccd1 vccd1 _16631_/C sky130_fd_sc_hd__a21bo_1
X_13842_ _13842_/A _13842_/B vssd1 vssd1 vccd1 vccd1 _13844_/B sky130_fd_sc_hd__and2_1
XFILLER_0_134_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12189__B _12269_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_1236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16561_ _21830_/Q _17520_/B _16561_/C _16586_/A vssd1 vssd1 vccd1 vccd1 _16586_/B
+ sky130_fd_sc_hd__nand4_2
X_13773_ _14713_/A _14713_/B _14234_/C vssd1 vssd1 vccd1 vccd1 _13773_/X sky130_fd_sc_hd__and3_1
XFILLER_0_58_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10985_ mstream_o[62] _10984_/Y _11005_/S vssd1 vssd1 vccd1 vccd1 _21599_/D sky130_fd_sc_hd__mux2_1
X_15512_ _15375_/A _16177_/B _15376_/A _15374_/B vssd1 vssd1 vccd1 vccd1 _15518_/A
+ sky130_fd_sc_hd__a31o_1
X_18300_ _18453_/A _18300_/B vssd1 vssd1 vccd1 vccd1 _18302_/B sky130_fd_sc_hd__and2_1
XFILLER_0_84_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12724_ _13975_/B _13258_/C _13258_/D _13682_/C vssd1 vssd1 vccd1 vccd1 _12725_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_29_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19280_ _19432_/A _19753_/B _19281_/C _19427_/A vssd1 vssd1 vccd1 vccd1 _19282_/B
+ sky130_fd_sc_hd__a22o_1
X_16492_ _16771_/A _16771_/B vssd1 vssd1 vccd1 vccd1 _16492_/X sky130_fd_sc_hd__and2_1
XFILLER_0_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18231_ _18230_/B _18230_/C _18230_/A vssd1 vssd1 vccd1 vccd1 _18231_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_128_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15443_ _15443_/A _15443_/B vssd1 vssd1 vccd1 vccd1 _15446_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__17996__A _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12655_ _12539_/X _12541_/X _12652_/X _12653_/Y vssd1 vssd1 vccd1 vccd1 _12655_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18162_ _18250_/A _18160_/Y _18017_/X _18020_/X vssd1 vssd1 vccd1 vccd1 _18163_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11606_ _13012_/B _12312_/A _11606_/C _11606_/D vssd1 vssd1 vccd1 vccd1 _11612_/B
+ sky130_fd_sc_hd__and4_1
X_15374_ _15374_/A _15374_/B vssd1 vssd1 vccd1 vccd1 _15376_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_142_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17325__A1 _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12586_ _12583_/X _12584_/Y _12475_/C _12475_/Y vssd1 vssd1 vccd1 vccd1 _12586_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_81_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17325__B2 _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14139__A1 _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11070__A0 _10867_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17113_ _17081_/A _17081_/C _17081_/B vssd1 vssd1 vccd1 vccd1 _17114_/C sky130_fd_sc_hd__o21bai_1
XFILLER_0_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14325_ _15155_/C _14477_/C _14635_/D _15159_/D vssd1 vssd1 vccd1 vccd1 _14328_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21311__A _21311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18093_ _17956_/Y _17958_/X _18091_/Y _18092_/X vssd1 vssd1 vccd1 vccd1 _18095_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11537_ _11089_/B t1y[29] t0x[29] _11543_/B2 vssd1 vssd1 vccd1 vccd1 _11537_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_151_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17044_ _17044_/A _17044_/B vssd1 vssd1 vccd1 vccd1 _17046_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14256_ _14255_/B _14255_/C _14255_/A vssd1 vssd1 vccd1 vccd1 _14258_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_29_1159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13748__B _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11468_ _11123_/A t1y[6] t0x[6] _21724_/D vssd1 vssd1 vccd1 vccd1 _11468_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_1_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11549__A _11549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13207_ _13204_/X _13205_/Y _13067_/B _13066_/Y vssd1 vssd1 vccd1 vccd1 _13209_/D
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_21_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14187_ _14183_/X _14185_/Y _14023_/X _14026_/X vssd1 vssd1 vccd1 vccd1 _14188_/B
+ sky130_fd_sc_hd__a211o_1
X_11399_ _11124_/A hold265/X fanout47/X hold153/X vssd1 vssd1 vccd1 vccd1 _11399_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15639__A1 _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ _12997_/A _12997_/C _12997_/B vssd1 vssd1 vccd1 vccd1 _13140_/C sky130_fd_sc_hd__a21bo_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13186__D _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18995_ _18995_/A _18995_/B _18708_/A vssd1 vssd1 vccd1 vccd1 _19160_/B sky130_fd_sc_hd__or3b_2
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13764__A _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13114__A2 _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ _12929_/B _12928_/Y _13067_/X _13068_/Y vssd1 vssd1 vccd1 vccd1 _13072_/B
+ sky130_fd_sc_hd__o211a_2
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17946_ _17942_/X _17944_/Y _17805_/B _17805_/Y vssd1 vssd1 vccd1 vccd1 _17948_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17877_ _18006_/B _17876_/C _17876_/A vssd1 vssd1 vccd1 vccd1 _17878_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_136_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19616_ _19616_/A _19616_/B vssd1 vssd1 vccd1 vccd1 _19617_/B sky130_fd_sc_hd__xnor2_4
X_16828_ _16828_/A _16828_/B vssd1 vssd1 vccd1 vccd1 _16836_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__14614__A2 _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19547_ _21839_/Q _19692_/B _19548_/C _19700_/A vssd1 vssd1 vccd1 vccd1 _19549_/B
+ sky130_fd_sc_hd__a22o_1
X_16759_ _17041_/A _16899_/B _17123_/C _17282_/A vssd1 vssd1 vccd1 vccd1 _16759_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_48_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19601__D _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19478_ _20770_/B _19476_/Y _19477_/X vssd1 vssd1 vccd1 vccd1 _19478_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21360__A2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18429_ _18849_/A _19223_/B _18429_/C _18429_/D vssd1 vssd1 vccd1 vccd1 _18430_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_1_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21440_ hold279/X sstream_i[17] _21489_/S vssd1 vssd1 vccd1 vccd1 _21967_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13050__A1 _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_942 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13050__B2 _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21371_ _21420_/S _18842_/B _21370_/Y vssd1 vssd1 vccd1 vccd1 _21371_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11600__A2 _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout216_A _21040_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20322_ _20322_/A _20466_/B vssd1 vssd1 vccd1 vccd1 _20325_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_102_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19069__A1 _19379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20253_ _20253_/A _20253_/B vssd1 vssd1 vccd1 vccd1 _20254_/B sky130_fd_sc_hd__nand2_1
XANTENNA__16969__B _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12561__B1 _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20184_ _20184_/A _20184_/B vssd1 vssd1 vccd1 vccd1 _20185_/B sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout585_A _11447_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16688__C _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17146__A _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20387__B1 _21258_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20926__A2 _21046_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14936__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout31_A _21490_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21707_ _22096_/CLK _21707_/D vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15030__A2 _14873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12440_ _12436_/X _12437_/Y _12331_/X _12333_/X vssd1 vssd1 vccd1 vccd1 _12475_/B
+ sky130_fd_sc_hd__a211oi_2
X_21638_ _21682_/CLK _21638_/D fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[101]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11052__A0 _11051_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15318__B1 _15976_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17858__A2 _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_clk_i clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _22096_/CLK sky130_fd_sc_hd__clkbuf_16
X_12371_ _12370_/B _12370_/C _12370_/A vssd1 vssd1 vccd1 vccd1 _12371_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_151_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21569_ mstream_o[32] _11043_/X _21579_/S vssd1 vssd1 vccd1 vccd1 _22096_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_35_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14110_ _14132_/B _14109_/B _14107_/X _14108_/Y vssd1 vssd1 vccd1 vccd1 _14110_/X
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_22_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11322_ _11544_/A1 t1x[24] v2z[24] _11223_/A _11321_/X vssd1 vssd1 vccd1 vccd1 _11322_/X
+ sky130_fd_sc_hd__a221o_2
X_15090_ _15632_/B _15091_/C _15001_/B _15892_/A vssd1 vssd1 vccd1 vccd1 _15090_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14041_ _14040_/B _14040_/C _14040_/A vssd1 vssd1 vccd1 vccd1 _14043_/B sky130_fd_sc_hd__a21o_1
X_11253_ _11122_/A t2y[7] t0y[7] _11123_/A vssd1 vssd1 vccd1 vccd1 _11253_/X sky130_fd_sc_hd__a22o_1
XANTENNA__12552__B1 _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11184_ hold301/X fanout51/X fanout47/X hold246/A vssd1 vssd1 vccd1 vccd1 _11184_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15097__A2 _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17800_ _17799_/B _17799_/C _17799_/A vssd1 vssd1 vccd1 vccd1 _17802_/B sky130_fd_sc_hd__a21o_1
X_15992_ _15992_/A vssd1 vssd1 vccd1 vccd1 _15992_/Y sky130_fd_sc_hd__inv_2
X_18780_ _18780_/A _18925_/B _18780_/C vssd1 vssd1 vccd1 vccd1 _18780_/X sky130_fd_sc_hd__and3_1
XFILLER_0_59_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14943_ _14944_/A _14944_/B vssd1 vssd1 vccd1 vccd1 _14943_/Y sky130_fd_sc_hd__nor2_1
X_17731_ _17865_/B _17731_/B vssd1 vssd1 vccd1 vccd1 _17734_/A sky130_fd_sc_hd__or2_1
XANTENNA__20378__B1 _21399_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11308__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14874_ _14874_/A _14874_/B vssd1 vssd1 vccd1 vccd1 _14881_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17662_ _17777_/B _17660_/X _17552_/X _17555_/A vssd1 vssd1 vccd1 vccd1 _17663_/B
+ sky130_fd_sc_hd__a211o_1
X_19401_ _19400_/B _19400_/C _19400_/A vssd1 vssd1 vccd1 vccd1 _19401_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13825_ _13827_/A _13979_/B vssd1 vssd1 vccd1 vccd1 _13828_/A sky130_fd_sc_hd__or2_1
XANTENNA__21088__A1_N _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16613_ _16613_/A _16613_/B _16613_/C vssd1 vssd1 vccd1 vccd1 _16625_/A sky130_fd_sc_hd__nand3_1
X_17593_ _17593_/A _17593_/B vssd1 vssd1 vccd1 vccd1 _17594_/B sky130_fd_sc_hd__nand2_1
X_16544_ _16544_/A _16544_/B vssd1 vssd1 vccd1 vccd1 _16547_/B sky130_fd_sc_hd__xnor2_1
X_19332_ _20838_/C _19331_/X _19330_/X vssd1 vssd1 vccd1 vccd1 _19334_/A sky130_fd_sc_hd__a21bo_1
X_13756_ _13756_/A _13756_/B vssd1 vssd1 vccd1 vccd1 _13758_/C sky130_fd_sc_hd__xor2_1
X_10968_ _10959_/A _10958_/Y _10967_/C _10967_/X _10961_/X vssd1 vssd1 vccd1 vccd1
+ _10972_/A sky130_fd_sc_hd__a311o_2
XANTENNA__21342__A2 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11551__B _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ _12825_/C _12707_/B vssd1 vssd1 vccd1 vccd1 _12957_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__14565__D _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16475_ _16476_/A _16476_/B vssd1 vssd1 vccd1 vccd1 _16475_/X sky130_fd_sc_hd__and2_1
XANTENNA__11291__B1 _11290_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19263_ _20650_/A _19906_/D _19264_/C _19264_/D vssd1 vssd1 vccd1 vccd1 _19266_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13687_ _13687_/A _13687_/B vssd1 vssd1 vccd1 vccd1 _13690_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10899_ _10899_/A _10899_/B vssd1 vssd1 vccd1 vccd1 _10902_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_156_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15426_ _15426_/A _15426_/B _15426_/C _15426_/D vssd1 vssd1 vccd1 vccd1 _15426_/Y
+ sky130_fd_sc_hd__nor4_4
X_18214_ _18215_/A _18215_/B _18215_/C vssd1 vssd1 vccd1 vccd1 _18214_/X sky130_fd_sc_hd__and3_1
XFILLER_0_66_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19194_ _19194_/A _19194_/B vssd1 vssd1 vccd1 vccd1 _19214_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_54_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12638_ _12637_/A _13152_/C _13152_/D _12750_/A vssd1 vssd1 vccd1 vccd1 _12639_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15309__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15357_ _21720_/Q hold167/A _10934_/Y fanout5/X vssd1 vssd1 vccd1 vccd1 _15357_/X
+ sky130_fd_sc_hd__a22o_1
X_18145_ _18032_/A _18031_/A _18031_/B vssd1 vssd1 vccd1 vccd1 _18150_/A sky130_fd_sc_hd__a21boi_2
X_12569_ _12460_/A _12460_/C _12460_/B vssd1 vssd1 vccd1 vccd1 _12570_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_41_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14308_ _14463_/D _15698_/B vssd1 vssd1 vccd1 vccd1 _14309_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_53_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18076_ _18077_/A _18077_/B _18077_/C vssd1 vssd1 vccd1 vccd1 _18076_/X sky130_fd_sc_hd__and3_1
X_15288_ _15288_/A _15288_/B vssd1 vssd1 vccd1 vccd1 _15290_/B sky130_fd_sc_hd__xnor2_1
Xhold206 hold206/A vssd1 vssd1 vccd1 vccd1 hold206/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold217 hold217/A vssd1 vssd1 vccd1 vccd1 hold217/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold228 hold228/A vssd1 vssd1 vccd1 vccd1 hold228/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_106_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17027_ _17028_/A _17028_/B _17028_/C vssd1 vssd1 vccd1 vccd1 _17038_/A sky130_fd_sc_hd__and3_1
X_14239_ _14237_/X _14239_/B vssd1 vssd1 vccd1 vccd1 _14240_/B sky130_fd_sc_hd__and2b_1
Xhold239 hold239/A vssd1 vssd1 vccd1 vccd1 hold239/X sky130_fd_sc_hd__buf_4
XFILLER_0_81_1150 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16285__A1 _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18978_ _18974_/X _18976_/Y _18813_/B _18813_/Y vssd1 vssd1 vccd1 vccd1 _18979_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17929_ _21824_/Q _19092_/C vssd1 vssd1 vccd1 vccd1 _17932_/A sky130_fd_sc_hd__and2_1
XANTENNA__12846__A1 _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16037__A1 _16036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20908__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19181__A _19337_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20940_ _21169_/A hold264/A hold294/A _21056_/A vssd1 vssd1 vccd1 vccd1 _20944_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16588__A2 _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20871_ _20872_/A _20872_/B _20872_/C vssd1 vssd1 vccd1 vccd1 _20871_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17413__B _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout166_A _21828_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21333__A2 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20541__B1 _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20774__B _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21423_ hold225/X sstream_i[0] _21442_/S vssd1 vssd1 vccd1 vccd1 _21950_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16045__A _16380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_934 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21354_ hold155/X fanout40/X _21353_/X vssd1 vssd1 vccd1 vccd1 _21925_/D sky130_fd_sc_hd__a21o_1
XFILLER_0_60_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13326__A2 _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20305_ _20302_/Y _20303_/X _20123_/Y _20162_/Y vssd1 vssd1 vccd1 vccd1 _20355_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_141_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18898__C _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21285_ _21285_/A _21285_/B vssd1 vssd1 vccd1 vccd1 _21300_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11337__B2 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20236_ _20386_/B _20236_/B vssd1 vssd1 vccd1 vccd1 _20381_/B sky130_fd_sc_hd__or2_2
X_20167_ _20167_/A _20167_/B vssd1 vssd1 vccd1 vccd1 _20210_/A sky130_fd_sc_hd__or2_1
XANTENNA__14826__A2 _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout79_A _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20098_ _20098_/A _20098_/B vssd1 vssd1 vccd1 vccd1 _20119_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13554__D _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17225__B1 _17324_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11940_ _11940_/A _11940_/B vssd1 vssd1 vccd1 vccd1 _11941_/C sky130_fd_sc_hd__xor2_1
XTAP_3635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17323__B _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11871_ _11823_/A _11823_/B _11823_/C vssd1 vssd1 vccd1 vccd1 _11871_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_58_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13610_ _14557_/B _14218_/B _14873_/B _14557_/A vssd1 vssd1 vccd1 vccd1 _13613_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_2967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10822_ hold74/A hold90/A vssd1 vssd1 vccd1 vccd1 _11050_/A sky130_fd_sc_hd__and2_1
XTAP_2978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14590_ _14591_/B _14591_/A vssd1 vssd1 vccd1 vccd1 _14590_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13541_ _13383_/X _13385_/Y _13538_/A _13539_/X vssd1 vssd1 vccd1 vccd1 _13541_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17977__C _19030_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12186__C _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16260_ _16152_/A _16152_/B _16193_/B vssd1 vssd1 vccd1 vccd1 _16300_/A sky130_fd_sc_hd__o21ai_1
X_13472_ _14572_/A _14234_/C vssd1 vssd1 vccd1 vccd1 _13475_/A sky130_fd_sc_hd__and2_1
XANTENNA__13014__A1 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14211__B1 _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__B2 _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15211_ _21720_/Q hold38/X _10926_/X fanout5/X _15210_/Y vssd1 vssd1 vccd1 vccd1
+ hold39/A sky130_fd_sc_hd__a221o_1
X_12423_ _12510_/A _12423_/B _12512_/A _15768_/A vssd1 vssd1 vccd1 vccd1 _12510_/B
+ sky130_fd_sc_hd__and4b_1
X_16191_ _16191_/A _16303_/B _16191_/C vssd1 vssd1 vccd1 vccd1 _16193_/B sky130_fd_sc_hd__or3_2
XANTENNA__21088__B2 _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11576__A1 _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11576__B2 _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15142_ _15006_/X _15012_/C _15253_/B _15141_/X vssd1 vssd1 vccd1 vccd1 _15298_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_2_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12354_ _12354_/A _12354_/B vssd1 vssd1 vccd1 vccd1 _12355_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15794__A _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11305_ _11325_/A1 t2y[20] t0y[20] _21723_/D vssd1 vssd1 vccd1 vccd1 _11305_/X sky130_fd_sc_hd__a22o_1
XANTENNA__16105__D _16418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15073_ _14942_/A _14942_/B _14943_/Y vssd1 vssd1 vccd1 vccd1 _15201_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19950_ _19950_/A _19950_/B vssd1 vssd1 vccd1 vccd1 _19958_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12285_ _12082_/X _12284_/Y _12081_/X vssd1 vssd1 vccd1 vccd1 _12288_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__11328__A1 _11327_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14024_ _14508_/A _14024_/B _15808_/C _14354_/C vssd1 vssd1 vccd1 vccd1 _14027_/D
+ sky130_fd_sc_hd__nand4_1
X_18901_ _19373_/B _19227_/D _18901_/C _18901_/D vssd1 vssd1 vccd1 vccd1 _18901_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11236_ _12268_/A _11235_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21760_/D sky130_fd_sc_hd__mux2_1
X_19881_ _19756_/B _19758_/B _19879_/X _19880_/Y vssd1 vssd1 vccd1 vccd1 _19885_/C
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__16267__A1 _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18832_ _18833_/B _18833_/C vssd1 vssd1 vccd1 vccd1 _18834_/B sky130_fd_sc_hd__nor2_2
X_11167_ hold170/X fanout23/X _11166_/X vssd1 vssd1 vccd1 vccd1 _11167_/X sky130_fd_sc_hd__a21o_1
XANTENNA__14203__A _14203_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15018__B _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18763_ _18604_/Y _18607_/X _18760_/Y _18761_/X vssd1 vssd1 vccd1 vccd1 _18763_/Y
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__11546__B _11555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15975_ _15978_/D vssd1 vssd1 vccd1 vccd1 _15975_/Y sky130_fd_sc_hd__inv_2
X_11098_ _11061_/X hold33/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21692_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17714_ _17715_/A _17715_/B vssd1 vssd1 vccd1 vccd1 _17850_/A sky130_fd_sc_hd__and2_2
XFILLER_0_26_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14926_ _14844_/A _14844_/C _14844_/B vssd1 vssd1 vccd1 vccd1 _14968_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17767__A1 _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18694_ _19185_/D _19013_/C _19179_/C _19008_/D vssd1 vssd1 vccd1 vccd1 _18698_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19124__B1_N _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11500__A1 _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14857__B _21765_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17767__B2 _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17645_ _17645_/A _17645_/B vssd1 vssd1 vccd1 vccd1 _17648_/A sky130_fd_sc_hd__xor2_2
X_14857_ _15076_/A _21765_/Q _21755_/Q _16380_/B vssd1 vssd1 vccd1 vccd1 _14976_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__11562__A _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19508__A2 _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15034__A _15933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13808_ _13548_/Y _13551_/X _13806_/X _13807_/Y vssd1 vssd1 vccd1 vccd1 _13818_/B
+ sky130_fd_sc_hd__a211o_1
X_14788_ _15702_/D _15579_/D _15717_/C _15976_/D vssd1 vssd1 vccd1 vccd1 _14946_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__13253__A1 _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17576_ _17575_/A _17575_/B _17575_/C _17575_/D vssd1 vssd1 vccd1 vccd1 _17576_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_97_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13253__B2 _14463_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21315__A2 _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14450__B1 _10886_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20034__A2_N _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11264__A0 _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19315_ _19316_/A _19316_/B vssd1 vssd1 vccd1 vccd1 _19317_/A sky130_fd_sc_hd__nor2_1
X_13739_ _13581_/A _13581_/Y _13736_/Y _13737_/X vssd1 vssd1 vccd1 vccd1 _13739_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_86_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16527_ _17636_/B _17282_/A vssd1 vssd1 vccd1 vccd1 _16531_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_156_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14873__A _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19246_ _19246_/A _19246_/B _19246_/C vssd1 vssd1 vccd1 vccd1 _19248_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_73_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16458_ _17206_/B _17019_/C vssd1 vssd1 vccd1 vccd1 _16462_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_115_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21079__A1 _21291_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15409_ _15412_/D vssd1 vssd1 vccd1 vccd1 _15409_/Y sky130_fd_sc_hd__inv_2
XANTENNA__21079__B2 _21293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16389_ _16321_/A _16320_/Y _16318_/X vssd1 vssd1 vccd1 vccd1 _16390_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19177_ _19083_/A _19083_/B _19082_/A vssd1 vssd1 vccd1 vccd1 _19216_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_83_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18128_ _18129_/A _18129_/B vssd1 vssd1 vccd1 vccd1 _18128_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18059_ _19438_/A _19438_/B _18640_/B _19092_/C vssd1 vssd1 vccd1 vccd1 _18061_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_44_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11319__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21070_ _20913_/Y _20917_/A _21068_/X _21069_/Y vssd1 vssd1 vccd1 vccd1 _21228_/A
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__18247__A2 _21358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout505 _16374_/A vssd1 vssd1 vccd1 vccd1 _16084_/A sky130_fd_sc_hd__buf_4
XANTENNA__16258__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20021_ _19985_/Y _20164_/A _20168_/B _20020_/D vssd1 vssd1 vccd1 vccd1 _20021_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
Xfanout516 _13875_/B vssd1 vssd1 vccd1 vccd1 _13018_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__16258__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout527 _21738_/Q vssd1 vssd1 vccd1 vccd1 _14027_/A sky130_fd_sc_hd__clkbuf_8
Xfanout538 _15439_/D vssd1 vssd1 vccd1 vccd1 _15153_/B sky130_fd_sc_hd__clkbuf_8
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout549 _13860_/A vssd1 vssd1 vccd1 vccd1 _12639_/A sky130_fd_sc_hd__clkbuf_8
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout283_A _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21972_ _21974_/CLK _21972_/D vssd1 vssd1 vccd1 vccd1 hold297/A sky130_fd_sc_hd__dfxtp_1
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13671__B _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20923_ _20924_/A _21264_/A _20924_/C _21097_/A vssd1 vssd1 vccd1 vccd1 _20925_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout450_A _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_1112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout548_A _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20854_ _20855_/A _20855_/B vssd1 vssd1 vccd1 vccd1 _20856_/A sky130_fd_sc_hd__nand2_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11255__B1 _11254_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14992__A1 _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20785_ _20786_/A _20786_/B vssd1 vssd1 vccd1 vccd1 _20785_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_14_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_638 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21406_ hold112/X _21381_/B _21405_/X vssd1 vssd1 vccd1 vccd1 _21943_/D sky130_fd_sc_hd__a21o_1
XANTENNA__12622__A2_N _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21337_ _21349_/A _21337_/B vssd1 vssd1 vccd1 vccd1 _21337_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12070_ _12070_/A _12118_/A vssd1 vssd1 vccd1 vccd1 _12071_/B sky130_fd_sc_hd__nor2_1
X_21268_ _21187_/Y _21231_/B _21186_/A vssd1 vssd1 vccd1 vccd1 _21269_/B sky130_fd_sc_hd__o21a_1
XANTENNA__12750__B _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11021_ mstream_o[95] hold6/X _11027_/S vssd1 vssd1 vccd1 vccd1 _21632_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11647__A _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20045__A2 _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20219_ _20070_/A _20070_/B _20068_/X vssd1 vssd1 vccd1 vccd1 _20220_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__14023__A _14508_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21199_ _21199_/A _21199_/B _21293_/B _21853_/Q vssd1 vssd1 vccd1 vccd1 _21287_/A
+ sky130_fd_sc_hd__nand4_2
X_15760_ _16363_/A hold112/X _10950_/Y fanout5/X _15759_/Y vssd1 vssd1 vccd1 vccd1
+ _15760_/X sky130_fd_sc_hd__a221o_1
XANTENNA__17334__A _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12972_ _13218_/A _12972_/B vssd1 vssd1 vccd1 vccd1 _13077_/A sky130_fd_sc_hd__nor2_1
XTAP_3421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14711_ _14711_/A _14711_/B vssd1 vssd1 vccd1 vccd1 _14739_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_87_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11923_ _11923_/A _11923_/B vssd1 vssd1 vccd1 vccd1 _11924_/C sky130_fd_sc_hd__xnor2_1
X_15691_ _15528_/Y _15567_/X _15689_/Y _15690_/X vssd1 vssd1 vccd1 vccd1 _15741_/A
+ sky130_fd_sc_hd__a211oi_4
XTAP_3454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14642_ _14631_/Y _14642_/B _14642_/C vssd1 vssd1 vccd1 vccd1 _14800_/A sky130_fd_sc_hd__and3b_1
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17430_ _17426_/X _17427_/Y _17312_/X _17314_/X vssd1 vssd1 vccd1 vccd1 _17466_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11854_ _11854_/A _11854_/B _11854_/C vssd1 vssd1 vccd1 vccd1 _11928_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_86_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ _10807_/A vssd1 vssd1 vccd1 vccd1 _10805_/Y sky130_fd_sc_hd__inv_2
X_14573_ _14419_/A _14419_/B _14974_/A vssd1 vssd1 vccd1 vccd1 _14575_/B sky130_fd_sc_hd__a21oi_2
X_17361_ _17382_/B _17360_/B _17360_/C _17360_/D vssd1 vssd1 vccd1 vccd1 _17362_/B
+ sky130_fd_sc_hd__o22a_1
XANTENNA__14693__A _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11785_ _11784_/A _11784_/C _11784_/B vssd1 vssd1 vccd1 vccd1 _11788_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_28_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19100_ _19099_/B _19099_/C _19099_/A vssd1 vssd1 vccd1 vccd1 _19101_/C sky130_fd_sc_hd__a21o_1
X_16312_ _16312_/A _16312_/B vssd1 vssd1 vccd1 vccd1 _16316_/A sky130_fd_sc_hd__nor2_1
X_13524_ _13525_/A _16399_/B _16409_/B _13394_/A vssd1 vssd1 vccd1 vccd1 _13545_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_67_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20845__D _20845_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17292_ _17293_/A _17293_/B vssd1 vssd1 vccd1 vccd1 _17292_/X sky130_fd_sc_hd__and2b_1
X_16243_ _16347_/B _16241_/X _16128_/A _16128_/Y vssd1 vssd1 vccd1 vccd1 _16243_/Y
+ sky130_fd_sc_hd__o211ai_2
X_19031_ _19650_/D _19201_/B _19032_/C _19032_/D vssd1 vssd1 vccd1 vccd1 _19031_/Y
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_152_221 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13455_ _13455_/A _13455_/B vssd1 vssd1 vccd1 vccd1 _13466_/A sky130_fd_sc_hd__or2_1
XFILLER_0_42_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12406_ _12406_/A _12406_/B vssd1 vssd1 vccd1 vccd1 _12408_/B sky130_fd_sc_hd__xnor2_1
X_16174_ _16284_/A _16286_/B _16284_/B vssd1 vssd1 vccd1 vccd1 _16176_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13386_ _13386_/A _13386_/B vssd1 vssd1 vccd1 vccd1 _13388_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13459__D _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15125_ _15126_/A _15126_/B vssd1 vssd1 vccd1 vccd1 _15328_/B sky130_fd_sc_hd__or2_1
XANTENNA__20861__C _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12337_ _12338_/A _12416_/A _12338_/C vssd1 vssd1 vccd1 vccd1 _12375_/A sky130_fd_sc_hd__and3_1
XFILLER_0_107_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15056_ _15056_/A _15056_/B vssd1 vssd1 vccd1 vccd1 _15059_/A sky130_fd_sc_hd__xor2_1
X_19933_ _19934_/A _19934_/B vssd1 vssd1 vccd1 vccd1 _20072_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12268_ _12268_/A _12268_/B vssd1 vssd1 vccd1 vccd1 _12268_/X sky130_fd_sc_hd__or2_1
XANTENNA__12660__B _13018_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14007_ _14007_/A vssd1 vssd1 vccd1 vccd1 _14007_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13171__B1 _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11219_ _14250_/B _11218_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21756_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18050__D _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19864_ _19737_/A _19737_/C _19737_/B vssd1 vssd1 vccd1 vccd1 _19879_/A sky130_fd_sc_hd__a21bo_1
X_12199_ _12199_/A _12199_/B _12199_/C vssd1 vssd1 vccd1 vccd1 _12200_/B sky130_fd_sc_hd__or3_1
X_18815_ _18664_/B _18664_/Y _18812_/X _18814_/Y vssd1 vssd1 vccd1 vccd1 _18815_/X
+ sky130_fd_sc_hd__a211o_2
X_19795_ hold126/X _19794_/X fanout4/X vssd1 vssd1 vccd1 vccd1 hold127/A sky130_fd_sc_hd__mux2_1
XFILLER_0_128_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18746_ _19686_/B _19529_/B _19068_/C _19238_/C _18598_/X vssd1 vssd1 vccd1 vccd1
+ _18755_/A sky130_fd_sc_hd__a41o_1
X_15958_ _15958_/A _16089_/B vssd1 vssd1 vccd1 vccd1 _15960_/A sky130_fd_sc_hd__or2_2
XANTENNA__13474__A1 _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13474__B2 _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14909_ _14909_/A _14909_/B vssd1 vssd1 vccd1 vccd1 _14910_/B sky130_fd_sc_hd__and2_1
XFILLER_0_78_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18677_ _18674_/X _18675_/Y _18521_/C _18520_/Y vssd1 vssd1 vccd1 vccd1 _18677_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13922__D _14234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15889_ _16363_/A hold124/X _10959_/Y fanout5/X vssd1 vssd1 vccd1 vccd1 _15889_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20101__C _21816_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17628_ _17629_/A _17629_/B _17629_/C vssd1 vssd1 vccd1 vccd1 _17630_/B sky130_fd_sc_hd__a21oi_4
XFILLER_0_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13226__A1 _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17898__B _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13226__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13777__A2 _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17559_ _17559_/A _17559_/B _17559_/C vssd1 vssd1 vccd1 vccd1 _17562_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18165__A1 _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18165__B2 _19230_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21213__B _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20570_ _20571_/A _20571_/B _20571_/C vssd1 vssd1 vccd1 vccd1 _20707_/A sky130_fd_sc_hd__a21o_1
XANTENNA__16307__B _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14726__A1 _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19229_ _19230_/A _19382_/B _19230_/C _19230_/D vssd1 vssd1 vccd1 vccd1 _19229_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14726__B2 _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13012__A _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout129_A _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19665__A1 _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19337__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21122_ _21232_/A _21122_/B _21236_/B _21122_/D vssd1 vssd1 vccd1 vccd1 _21232_/B
+ sky130_fd_sc_hd__nor4_1
XFILLER_0_100_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16042__B _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19056__D _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout302 _21795_/Q vssd1 vssd1 vccd1 vccd1 _19493_/D sky130_fd_sc_hd__buf_2
XANTENNA_fanout498_A _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21053_ _21207_/B _21053_/B vssd1 vssd1 vccd1 vccd1 _21069_/A sky130_fd_sc_hd__and2_1
Xfanout313 _17141_/C vssd1 vssd1 vccd1 vccd1 _17145_/B sky130_fd_sc_hd__buf_4
Xfanout324 _18859_/A vssd1 vssd1 vccd1 vccd1 _18703_/A sky130_fd_sc_hd__clkbuf_8
Xfanout335 _16399_/B vssd1 vssd1 vccd1 vccd1 _16084_/C sky130_fd_sc_hd__buf_4
Xfanout346 _16396_/B vssd1 vssd1 vccd1 vccd1 _15717_/C sky130_fd_sc_hd__buf_4
Xfanout357 _16391_/A vssd1 vssd1 vccd1 vccd1 _15653_/C sky130_fd_sc_hd__buf_4
XANTENNA__11712__B2 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20004_ _20689_/A _20562_/B _20924_/A _21305_/A vssd1 vssd1 vccd1 vccd1 _20143_/A
+ sky130_fd_sc_hd__and4_1
Xfanout368 _15916_/B vssd1 vssd1 vccd1 vccd1 _16371_/A sky130_fd_sc_hd__buf_4
XANTENNA__19353__B _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout379 _14828_/B vssd1 vssd1 vccd1 vccd1 _16284_/A sky130_fd_sc_hd__buf_2
XANTENNA__11617__D _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19196__A3 _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14928__D _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21955_ _21963_/CLK _21955_/D vssd1 vssd1 vccd1 vccd1 hold255/A sky130_fd_sc_hd__dfxtp_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_115_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20906_ _20906_/A _20906_/B vssd1 vssd1 vccd1 vccd1 _20906_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21886_ _21926_/CLK _21886_/D vssd1 vssd1 vccd1 vccd1 hold194/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_96_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21404__A _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20837_ _21199_/A _21286_/B _21296_/B _20838_/B vssd1 vssd1 vccd1 vccd1 _20841_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11930__A _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11570_ _12229_/A _12528_/B _12619_/A _12155_/B vssd1 vssd1 vccd1 vccd1 _11571_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11243__A3 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20768_ _20900_/A _20645_/B _20640_/X vssd1 vssd1 vccd1 vccd1 _20769_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14663__D _14663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18135__D _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14018__A _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18713__A _19337_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11141__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20699_ _20699_/A _20699_/B _20699_/C vssd1 vssd1 vccd1 vccd1 _20700_/A sky130_fd_sc_hd__and3_1
XFILLER_0_134_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13240_ _13240_/A _13240_/B vssd1 vssd1 vccd1 vccd1 _13242_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_126_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18432__B _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20266__A2 _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13171_ _15076_/B _13034_/D _14386_/B _15076_/A vssd1 vssd1 vccd1 vccd1 _13171_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_60_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11951__A1 _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12122_ _12066_/X _12085_/Y _12115_/A _12114_/Y vssd1 vssd1 vccd1 vccd1 _12124_/C
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__11951__B2 _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19408__A1 _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19408__B2 _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12911__D _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16930_ _16930_/A _16930_/B _16930_/C vssd1 vssd1 vccd1 vccd1 _16982_/A sky130_fd_sc_hd__nand3_1
X_12053_ _12053_/A _12053_/B _12053_/C vssd1 vssd1 vccd1 vccd1 _12066_/A sky130_fd_sc_hd__and3_1
XANTENNA__13295__C _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11004_ mstream_o[78] hold10/X _11005_/S vssd1 vssd1 vccd1 vccd1 _21615_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_99_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15791__B _15916_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16861_ _17145_/A _16968_/C vssd1 vssd1 vccd1 vccd1 _16863_/B sky130_fd_sc_hd__and2_1
X_18600_ _18597_/Y _18598_/X _18464_/D _18465_/B vssd1 vssd1 vccd1 vccd1 _18601_/B
+ sky130_fd_sc_hd__o211ai_1
X_15812_ _15813_/A _15813_/B vssd1 vssd1 vccd1 vccd1 _15940_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_137_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17064__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19580_ _19581_/A _19581_/B _19581_/C vssd1 vssd1 vccd1 vccd1 _19580_/X sky130_fd_sc_hd__and3_1
XANTENNA__13456__A1 _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16792_ _16792_/A _16792_/B vssd1 vssd1 vccd1 vccd1 _17372_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_137_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18531_ _18380_/Y _18382_/Y _18684_/B _18530_/Y vssd1 vssd1 vccd1 vccd1 _18687_/A
+ sky130_fd_sc_hd__o211ai_4
X_15743_ _15612_/A _15612_/Y _15741_/X _15742_/Y vssd1 vssd1 vccd1 vccd1 _15743_/Y
+ sky130_fd_sc_hd__o211ai_4
XTAP_3240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12955_ hold221/X _12954_/X fanout3/X vssd1 vssd1 vccd1 vccd1 _21860_/D sky130_fd_sc_hd__mux2_1
XTAP_3251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13742__D _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11316__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11906_ _11905_/A _11905_/Y _11840_/X _11841_/Y vssd1 vssd1 vccd1 vccd1 _11907_/A
+ sky130_fd_sc_hd__o211a_1
XTAP_3284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18462_ _19695_/A _19686_/A _18767_/B _18616_/D vssd1 vssd1 vccd1 vccd1 _18464_/D
+ sky130_fd_sc_hd__nand4_4
X_15674_ _15933_/C _16377_/B _15672_/Y _15802_/A vssd1 vssd1 vccd1 vccd1 _15676_/A
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_3295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_240 hold309/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12886_ _12877_/A _13157_/B _12757_/X _12756_/X _13155_/C vssd1 vssd1 vccd1 vccd1
+ _12887_/C sky130_fd_sc_hd__a32o_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_251 _21825_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_262 hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17413_ _17619_/B _20910_/A _17413_/C _17413_/D vssd1 vssd1 vccd1 vccd1 _17415_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA_273 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14625_ _14625_/A _14625_/B vssd1 vssd1 vccd1 vccd1 _14627_/A sky130_fd_sc_hd__xnor2_1
X_11837_ _11836_/A _11836_/Y _11805_/X _11806_/Y vssd1 vssd1 vccd1 vccd1 _11840_/A
+ sky130_fd_sc_hd__a211oi_4
XANTENNA_284 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18393_ hold34/X _18392_/X fanout2/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__mux2_1
XFILLER_0_28_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_295 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15441__A2_N _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18147__A1 _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18147__B2 _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14556_ _14557_/B _15510_/B _14557_/D _14557_/A vssd1 vssd1 vccd1 vccd1 _14559_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17344_ _17343_/A _17343_/B _17343_/C vssd1 vssd1 vccd1 vccd1 _17345_/C sky130_fd_sc_hd__a21o_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ _11767_/A _11767_/C _11767_/B vssd1 vssd1 vccd1 vccd1 _11772_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_82_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12431__A2 _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13507_ _13503_/Y _13505_/X _13248_/Y _13251_/Y vssd1 vssd1 vccd1 vccd1 _13508_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_83_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14487_ _14647_/A _14485_/Y _14331_/B _14333_/B vssd1 vssd1 vccd1 vccd1 _14488_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_15_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17275_ _17197_/A _17197_/B _17198_/A _17195_/X vssd1 vssd1 vccd1 vccd1 _17366_/A
+ sky130_fd_sc_hd__a31oi_4
X_11699_ _11699_/A _12318_/A _11699_/C vssd1 vssd1 vccd1 vccd1 _12318_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_114_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19014_ _19179_/C _19013_/X _19012_/X vssd1 vssd1 vccd1 vccd1 _19016_/A sky130_fd_sc_hd__a21bo_1
X_16226_ _16226_/A _16226_/B _16226_/C vssd1 vssd1 vccd1 vccd1 _16226_/X sky130_fd_sc_hd__and3_1
X_13438_ _14024_/B _14537_/A _13437_/C _13437_/D vssd1 vssd1 vccd1 vccd1 _13439_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16157_ _16418_/A _16377_/A _16157_/C _16157_/D vssd1 vssd1 vccd1 vccd1 _16324_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__17658__B1 _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13369_ fanout9/X _13369_/B vssd1 vssd1 vccd1 vccd1 _13369_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15108_ _15108_/A _15108_/B _15254_/B _15108_/D vssd1 vssd1 vccd1 vccd1 _15250_/B
+ sky130_fd_sc_hd__or4_2
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16088_ _16088_/A _16201_/B vssd1 vssd1 vccd1 vccd1 _16091_/A sky130_fd_sc_hd__or2_1
XFILLER_0_11_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18870__A2 _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15039_ _14833_/A _14833_/C _14833_/B vssd1 vssd1 vccd1 vccd1 _15040_/C sky130_fd_sc_hd__a21bo_1
X_19916_ _19914_/A _19914_/B _19914_/C vssd1 vssd1 vccd1 vccd1 _19917_/C sky130_fd_sc_hd__a21o_1
X_19847_ _19847_/A _19847_/B vssd1 vssd1 vccd1 vccd1 _19847_/X sky130_fd_sc_hd__or2_1
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19778_ _19779_/A _19779_/B _19779_/C vssd1 vssd1 vccd1 vccd1 _19942_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_39_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18729_ _18569_/Y _18572_/X _18846_/A _18728_/X vssd1 vssd1 vccd1 vccd1 _18846_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__17124__D _17141_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21740_ _22021_/CLK _21740_/D vssd1 vssd1 vccd1 vccd1 _21740_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_94_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21671_ _21906_/CLK _21671_/D vssd1 vssd1 vccd1 vccd1 hold69/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__18138__A1 _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout246_A _21807_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20622_ _20621_/B _20621_/C _20621_/A vssd1 vssd1 vccd1 vccd1 _20622_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_129_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12422__A2 _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12565__B _12785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20553_ _20554_/A _20554_/B vssd1 vssd1 vccd1 vccd1 _20742_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_85_1115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout413_A _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15372__A1 _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14175__A2 _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15372__B2 _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20484_ _20484_/A _20484_/B vssd1 vssd1 vccd1 vccd1 _20486_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_6_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15892__A _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21105_ _21105_/A _21105_/B vssd1 vssd1 vccd1 vccd1 _21107_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__20006__C _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16203__D _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22085_ _22096_/CLK _22085_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[21] sky130_fd_sc_hd__dfrtp_4
Xfanout110 _19692_/C vssd1 vssd1 vccd1 vccd1 _20416_/A sky130_fd_sc_hd__buf_4
Xfanout121 _21838_/Q vssd1 vssd1 vccd1 vccd1 _20562_/B sky130_fd_sc_hd__buf_4
XFILLER_0_121_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout132 _19087_/B vssd1 vssd1 vccd1 vccd1 _20774_/B sky130_fd_sc_hd__buf_4
XFILLER_0_100_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21036_ _21301_/A _21283_/A _21264_/B _21151_/A vssd1 vssd1 vccd1 vccd1 _21040_/C
+ sky130_fd_sc_hd__a22o_1
Xfanout143 _18624_/A vssd1 vssd1 vccd1 vccd1 _20650_/A sky130_fd_sc_hd__clkbuf_8
Xfanout154 _21831_/Q vssd1 vssd1 vccd1 vccd1 _19092_/A sky130_fd_sc_hd__buf_4
Xfanout165 _16813_/A vssd1 vssd1 vccd1 vccd1 _17029_/A sky130_fd_sc_hd__buf_4
Xfanout176 _16734_/B vssd1 vssd1 vccd1 vccd1 _17129_/B sky130_fd_sc_hd__buf_4
XANTENNA__16500__B _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11161__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15427__A2 _15426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout187 _21824_/Q vssd1 vssd1 vccd1 vccd1 _19445_/A sky130_fd_sc_hd__buf_4
XANTENNA__13438__A1 _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout198 hold264/A vssd1 vssd1 vccd1 vccd1 _21258_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout61_A _10791_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11449__A0 _11448_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14020__B _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12740_ _12741_/A _12741_/B vssd1 vssd1 vccd1 vccd1 _12868_/B sky130_fd_sc_hd__nand2_1
X_21938_ _21938_/CLK _21938_/D vssd1 vssd1 vccd1 vccd1 hold87/A sky130_fd_sc_hd__dfxtp_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12661__A2 _12771_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18427__B _18873_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ _13155_/A _12781_/D _12668_/Y _12669_/X vssd1 vssd1 vccd1 vccd1 _12672_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__14938__B2 _14774_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21869_ _21942_/CLK _21869_/D vssd1 vssd1 vccd1 vccd1 hold157/A sky130_fd_sc_hd__dfxtp_1
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12756__A _14024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14410_ _14409_/B _14554_/B _14409_/A vssd1 vssd1 vccd1 vccd1 _14411_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_33_1250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14674__C _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18146__C _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11622_ _11623_/A _11623_/B vssd1 vssd1 vccd1 vccd1 _11672_/A sky130_fd_sc_hd__or2_1
XFILLER_0_155_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15390_ _15717_/B _16196_/B _15911_/A _15911_/C vssd1 vssd1 vccd1 vccd1 _15588_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13610__A1 _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13610__B2 _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14341_ _14341_/A _14341_/B vssd1 vssd1 vccd1 vccd1 _14343_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_107_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11553_ _21412_/A _11551_/Y _21329_/B1 vssd1 vssd1 vccd1 vccd1 _11553_/Y sky130_fd_sc_hd__o21ai_4
XFILLER_0_65_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17060_ _17038_/A _17038_/C _17038_/B vssd1 vssd1 vccd1 vccd1 _17060_/Y sky130_fd_sc_hd__o21ai_1
X_14272_ _14268_/X _14269_/Y _14107_/X _14109_/X vssd1 vssd1 vccd1 vccd1 _14273_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_123_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11484_ _11502_/A1 t2x[11] v1z[11] fanout20/X _11483_/X vssd1 vssd1 vccd1 vccd1 _11484_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_52_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16011_ _16011_/A _16011_/B vssd1 vssd1 vccd1 vccd1 _16014_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_123_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13223_ _13223_/A _13365_/A vssd1 vssd1 vccd1 vccd1 _13518_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13154_ _13154_/A _13154_/B vssd1 vssd1 vccd1 vccd1 _13162_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_1054 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_103_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12105_ _12106_/A _12106_/B vssd1 vssd1 vccd1 vccd1 _12120_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_104_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17962_ _17962_/A _17962_/B _17962_/C vssd1 vssd1 vccd1 vccd1 _17964_/A sky130_fd_sc_hd__nor3_2
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13085_ _13085_/A _13085_/B vssd1 vssd1 vccd1 vccd1 _13088_/B sky130_fd_sc_hd__nor2_2
X_19701_ _20103_/A _19906_/C _19565_/X _19566_/X _19868_/B vssd1 vssd1 vccd1 vccd1
+ _19706_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_100_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16913_ _16912_/A _16912_/B _17372_/B vssd1 vssd1 vccd1 vccd1 _16914_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__18065__B1 _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12036_ _12036_/A _12036_/B _12036_/C vssd1 vssd1 vccd1 vccd1 _12036_/X sky130_fd_sc_hd__and3_1
XANTENNA__19801__A1 _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17893_ _18008_/A _18769_/B vssd1 vssd1 vccd1 vccd1 _17897_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19801__B2 _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11152__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19632_ _19634_/B _19634_/A vssd1 vssd1 vccd1 vccd1 _19632_/Y sky130_fd_sc_hd__nand2b_1
X_16844_ _16844_/A _16844_/B _16849_/C _16844_/D vssd1 vssd1 vccd1 vccd1 _16844_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_18_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11554__B _11555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19563_ _19563_/A _19563_/B vssd1 vssd1 vccd1 vccd1 _19583_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_88_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16775_ _16783_/A _16773_/Y _16764_/X _16770_/X vssd1 vssd1 vccd1 vccd1 _16776_/D
+ sky130_fd_sc_hd__a211o_1
X_13987_ _13987_/A vssd1 vssd1 vccd1 vccd1 _13989_/B sky130_fd_sc_hd__inv_2
XFILLER_0_34_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19565__B1 _19868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11046__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18514_ _18510_/X _18512_/Y _18363_/B _18363_/Y vssd1 vssd1 vccd1 vccd1 _18516_/D
+ sky130_fd_sc_hd__o211a_1
X_15726_ _15727_/A _15727_/B _15727_/C vssd1 vssd1 vccd1 vccd1 _15726_/X sky130_fd_sc_hd__a21o_1
XTAP_3070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17522__A _17619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19494_ _19496_/A vssd1 vssd1 vccd1 vccd1 _19658_/A sky130_fd_sc_hd__inv_2
X_12938_ _12938_/A _12938_/B _12938_/C vssd1 vssd1 vccd1 vccd1 _12938_/Y sky130_fd_sc_hd__nand3_4
XTAP_3092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_778 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14929__A1 _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18445_ _19051_/A _19240_/B _18443_/Y _18594_/A vssd1 vssd1 vccd1 vccd1 _18445_/X
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12088__D _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15657_ _15916_/B _16040_/C _16396_/A _15791_/A vssd1 vssd1 vccd1 vccd1 _15661_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15051__B1 _15050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ _12869_/A _12869_/B _12869_/C vssd1 vssd1 vccd1 vccd1 _12869_/X sky130_fd_sc_hd__and3_2
XFILLER_0_8_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_1069 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14608_ _14608_/A _14608_/B vssd1 vssd1 vccd1 vccd1 _14759_/A sky130_fd_sc_hd__or2_2
X_18376_ _18373_/X _18374_/Y _18225_/B _18224_/Y vssd1 vssd1 vccd1 vccd1 _18377_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12404__A2 _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15588_ _15588_/A _15588_/B vssd1 vssd1 vccd1 vccd1 _15596_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17327_ _17327_/A _17327_/B vssd1 vssd1 vccd1 vccd1 _17329_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_71_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14539_ _15373_/B _16268_/B _16266_/C _14698_/A vssd1 vssd1 vccd1 vccd1 _14543_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17258_ _16657_/C _16656_/Y _17256_/X _17257_/Y vssd1 vssd1 vccd1 vccd1 _17363_/A
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_109_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16209_ _16209_/A _16209_/B vssd1 vssd1 vccd1 vccd1 _16211_/B sky130_fd_sc_hd__or2_1
XFILLER_0_3_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17189_ _16549_/A _16548_/B _16546_/A vssd1 vssd1 vccd1 vccd1 _17191_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_12_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18843__A2 fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11391__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12551__D _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17416__B _20249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11143__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12340__A1 _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15217__A _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout363_A _21778_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20777__B _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17031__A1 _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21723_ _21845_/CLK _21723_/D fanout639/X vssd1 vssd1 vccd1 vccd1 _21723_/Q sky130_fd_sc_hd__dfrtp_1
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11851__B1 _12637_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__16048__A _16273_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout628_A _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21654_ _21888_/CLK _21654_/D vssd1 vssd1 vccd1 vccd1 hold143/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__11911__C _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20605_ _20608_/D vssd1 vssd1 vccd1 vccd1 _20605_/Y sky130_fd_sc_hd__inv_2
XANTENNA__11603__B1 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21585_ _21888_/CLK _21585_/D fanout640/X vssd1 vssd1 vccd1 vccd1 mstream_o[48] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_90_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1081 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20536_ _20536_/A _20665_/B vssd1 vssd1 vccd1 vccd1 _20539_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_117_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16542__B1 _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20467_ _20466_/A _20466_/B _20466_/C vssd1 vssd1 vccd1 vccd1 _20468_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_132_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11639__B _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20398_ _20398_/A _20398_/B vssd1 vssd1 vccd1 vccd1 _20399_/B sky130_fd_sc_hd__xor2_1
XANTENNA__17029__D _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11382__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16511__A _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14856__B1 _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22068_ _22069_/CLK _22068_/D fanout639/X vssd1 vssd1 vccd1 vccd1 mstream_o[4] sky130_fd_sc_hd__dfrtp_4
XANTENNA__11134__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13910_ _13910_/A _13910_/B vssd1 vssd1 vccd1 vccd1 _13919_/A sky130_fd_sc_hd__nand2_1
X_21019_ _20886_/X _20888_/Y _21129_/B _21018_/X vssd1 vssd1 vccd1 vccd1 _21135_/A
+ sky130_fd_sc_hd__a211oi_2
X_14890_ _14739_/A _14739_/B _14737_/Y vssd1 vssd1 vccd1 vccd1 _14892_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__13573__C _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1003 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10893__A1 _10892_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13841_ _13838_/Y _13839_/X _13707_/D _13708_/B vssd1 vssd1 vccd1 vccd1 _13842_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_134_1215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13772_ _14713_/B _14234_/C _15370_/B _14713_/A vssd1 vssd1 vccd1 vccd1 _13772_/X
+ sky130_fd_sc_hd__a22o_1
X_16560_ _16813_/A _16743_/B _17223_/A _16860_/C vssd1 vssd1 vccd1 vccd1 _16586_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__12095__B1 _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10984_ _10984_/A _10984_/B vssd1 vssd1 vccd1 vccd1 _10984_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_70_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15511_ _15511_/A _15670_/B vssd1 vssd1 vccd1 vccd1 _15519_/A sky130_fd_sc_hd__nand2_1
X_12723_ _12851_/A vssd1 vssd1 vccd1 vccd1 _12725_/C sky130_fd_sc_hd__inv_2
XFILLER_0_57_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16491_ _16495_/B _16491_/B vssd1 vssd1 vccd1 vccd1 _16771_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_155_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_759 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18230_ _18230_/A _18230_/B _18230_/C vssd1 vssd1 vccd1 vccd1 _18230_/Y sky130_fd_sc_hd__nand3_2
X_15442_ _15442_/A _15442_/B vssd1 vssd1 vccd1 vccd1 _15443_/B sky130_fd_sc_hd__nor2_1
XANTENNA__21626__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12654_ _12539_/X _12541_/X _12652_/X _12653_/Y vssd1 vssd1 vccd1 vccd1 _12692_/A
+ sky130_fd_sc_hd__o211a_2
XANTENNA__17996__B _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11605_ _11612_/A vssd1 vssd1 vccd1 vccd1 _11606_/D sky130_fd_sc_hd__inv_2
XFILLER_0_143_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18161_ _18017_/X _18020_/X _18250_/A _18160_/Y vssd1 vssd1 vccd1 vccd1 _18250_/B
+ sky130_fd_sc_hd__o211ai_1
X_15373_ _15373_/A _15373_/B _16286_/B _16027_/B vssd1 vssd1 vccd1 vccd1 _15374_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_108_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12585_ _12475_/C _12475_/Y _12583_/X _12584_/Y vssd1 vssd1 vccd1 vccd1 _12585_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_136_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17325__A2 _19430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17112_ _17046_/A _17046_/C _17046_/B vssd1 vssd1 vccd1 vccd1 _17114_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__15411__A1_N _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14324_ _15155_/C _15788_/B _14175_/X _14176_/X _15112_/D vssd1 vssd1 vccd1 vccd1
+ _14329_/A sky130_fd_sc_hd__a32o_1
X_11536_ _11535_/X _19179_/C _11545_/S vssd1 vssd1 vccd1 vccd1 _21850_/D sky130_fd_sc_hd__mux2_1
XANTENNA__21311__B _21311_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18092_ _18091_/B _18091_/C _18091_/A vssd1 vssd1 vccd1 vccd1 _18092_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_41_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_987 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14255_ _14255_/A _14255_/B _14255_/C vssd1 vssd1 vccd1 vccd1 _14258_/A sky130_fd_sc_hd__nand3_1
X_17043_ _17044_/A _17044_/B vssd1 vssd1 vccd1 vccd1 _17049_/A sky130_fd_sc_hd__nor2_1
X_11467_ _11466_/X _18058_/A _11470_/S vssd1 vssd1 vccd1 vccd1 _21827_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13748__C _14212_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18901__A _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13206_ _13067_/B _13066_/Y _13204_/X _13205_/Y vssd1 vssd1 vccd1 vccd1 _13209_/C
+ sky130_fd_sc_hd__o211a_4
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14186_ _14023_/X _14026_/X _14183_/X _14185_/Y vssd1 vssd1 vccd1 vccd1 _14186_/X
+ sky130_fd_sc_hd__o211a_1
X_11398_ _11397_/X _18166_/A _11401_/S vssd1 vssd1 vccd1 vccd1 _21804_/D sky130_fd_sc_hd__mux2_1
XANTENNA__11373__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13137_ _13136_/B _13136_/C _13136_/A vssd1 vssd1 vccd1 vccd1 _13140_/B sky130_fd_sc_hd__a21o_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18994_ _19155_/B _18992_/Y _18830_/B _18833_/B vssd1 vssd1 vccd1 vccd1 _18995_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13764__B _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13068_ _13067_/B _13067_/C _13067_/A vssd1 vssd1 vccd1 vccd1 _13068_/Y sky130_fd_sc_hd__o21ai_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17945_ _17805_/B _17805_/Y _17942_/X _17944_/Y vssd1 vssd1 vccd1 vccd1 _17948_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_29_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_1051 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12019_ _12019_/A _12019_/B vssd1 vssd1 vccd1 vccd1 _12070_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_40_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19732__A _19732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17876_ _17876_/A _18006_/B _17876_/C vssd1 vssd1 vccd1 vccd1 _17878_/B sky130_fd_sc_hd__nand3_1
X_19615_ _19616_/B _19616_/A vssd1 vssd1 vccd1 vccd1 _19615_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_136_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16827_ _16754_/Y _16824_/X _16823_/X _16809_/X vssd1 vssd1 vccd1 vccd1 _16844_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__14876__A _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16794__C _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19546_ _19906_/A _20146_/B _19705_/B _19546_/D vssd1 vssd1 vccd1 vccd1 _19700_/A
+ sky130_fd_sc_hd__nand4_2
X_16758_ _16758_/A _16758_/B vssd1 vssd1 vccd1 vccd1 _16765_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_45_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15709_ _15709_/A _15709_/B vssd1 vssd1 vccd1 vccd1 _15712_/B sky130_fd_sc_hd__xnor2_2
X_19477_ hold111/A fanout7/X _14605_/B _19636_/A vssd1 vssd1 vccd1 vccd1 _19477_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_16689_ _17145_/A _17223_/A vssd1 vssd1 vccd1 vccd1 _16691_/B sky130_fd_sc_hd__and2_1
XFILLER_0_29_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18428_ _18849_/A _19223_/B _18429_/C _18429_/D vssd1 vssd1 vccd1 vccd1 _18430_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18359_ _18209_/A _18209_/C _18209_/B vssd1 vssd1 vccd1 vccd1 _18360_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__19179__A _19650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13050__A2 _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21370_ _21420_/S _13967_/X _21421_/S vssd1 vssd1 vccd1 vccd1 _21370_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_976 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20321_ _20321_/A _20321_/B _20321_/C vssd1 vssd1 vccd1 vccd1 _20466_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_3_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout111_A _21267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19069__A2 _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout209_A _21815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20252_ _20253_/A _20253_/B vssd1 vssd1 vccd1 vccd1 _20252_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_3_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11364__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12561__A1 _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12561__B2 _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20183_ _20184_/A _20184_/B vssd1 vssd1 vccd1 vccd1 _20183_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_0_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18029__B1 _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16688__D _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17146__B _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout480_A _14217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout578_A _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20387__A1 _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20387__B2 _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10875__A1 _10874_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11625__D _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14936__D _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15015__B1 _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1075 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21706_ _22096_/CLK _21706_/D vssd1 vssd1 vccd1 vccd1 hold168/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout24_A _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21412__A _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21637_ _21722_/CLK _21637_/D fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[100]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__19089__A _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15410__A _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12370_ _12370_/A _12370_/B _12370_/C vssd1 vssd1 vccd1 vccd1 _12370_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__20311__A1 _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21568_ mstream_o[31] hold67/X _21568_/S vssd1 vssd1 vccd1 vccd1 _22095_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_117_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11321_ _11325_/A1 t2y[24] t0y[24] _21723_/D vssd1 vssd1 vccd1 vccd1 _11321_/X sky130_fd_sc_hd__a22o_1
X_20519_ _20774_/B _21258_/B _21171_/B _20774_/A vssd1 vssd1 vccd1 vccd1 _20523_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14026__A _14027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21499_ hold303/X sstream_i[76] _21510_/S vssd1 vssd1 vccd1 vccd1 _22026_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14040_ _14040_/A _14040_/B _14040_/C vssd1 vssd1 vccd1 vccd1 _14043_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_105_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11252_ _12229_/A _11251_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21764_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_31_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11355__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12552__A1 _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17337__A _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12552__B2 _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11183_ _13034_/D _11182_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21744_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15991_ _15991_/A _15991_/B _15991_/C vssd1 vssd1 vccd1 vccd1 _15992_/A sky130_fd_sc_hd__or3_2
XFILLER_0_98_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17730_ _18851_/C _19060_/B _17865_/A _17728_/Y vssd1 vssd1 vccd1 vccd1 _17731_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14942_ _14942_/A _14942_/B vssd1 vssd1 vccd1 vccd1 _14944_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__20378__B2 _11550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18797__A2_N _19753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17661_ _17552_/X _17555_/A _17777_/B _17660_/X vssd1 vssd1 vccd1 vccd1 _17661_/X
+ sky130_fd_sc_hd__o211a_1
X_14873_ _16027_/A _14873_/B vssd1 vssd1 vccd1 vccd1 _14874_/B sky130_fd_sc_hd__nand2_1
X_19400_ _19400_/A _19400_/B _19400_/C vssd1 vssd1 vccd1 vccd1 _19400_/X sky130_fd_sc_hd__and3_1
X_16612_ _21822_/Q _17657_/A _17334_/B _21823_/Q vssd1 vssd1 vccd1 vccd1 _16613_/C
+ sky130_fd_sc_hd__a22o_1
X_13824_ _13979_/A _16404_/B _13983_/B _13824_/D vssd1 vssd1 vccd1 vccd1 _13979_/B
+ sky130_fd_sc_hd__and4b_1
X_17592_ _17705_/B _17592_/B vssd1 vssd1 vccd1 vccd1 _17595_/A sky130_fd_sc_hd__xnor2_4
XFILLER_0_106_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19331_ _19487_/B _19650_/D _20838_/D vssd1 vssd1 vccd1 vccd1 _19331_/X sky130_fd_sc_hd__and3_1
X_16543_ _16541_/X _16543_/B vssd1 vssd1 vccd1 vccd1 _16544_/B sky130_fd_sc_hd__and2b_1
X_13755_ _13756_/A _13756_/B vssd1 vssd1 vccd1 vccd1 _13755_/X sky130_fd_sc_hd__or2_1
X_10967_ hold208/A hold226/A _10967_/C vssd1 vssd1 vccd1 vccd1 _10967_/X sky130_fd_sc_hd__and3_1
XFILLER_0_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11324__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19262_ _19972_/A _20394_/B _19262_/C _19414_/C vssd1 vssd1 vccd1 vccd1 _19264_/D
+ sky130_fd_sc_hd__nand4_4
X_12706_ _12825_/A _12596_/B _12831_/D vssd1 vssd1 vccd1 vccd1 _12707_/B sky130_fd_sc_hd__o21ba_1
X_16474_ _16474_/A _16474_/B vssd1 vssd1 vccd1 vccd1 _16476_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_57_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13686_ _13687_/A _13687_/B vssd1 vssd1 vccd1 vccd1 _13686_/Y sky130_fd_sc_hd__nand2_1
X_10898_ hold216/A hold217/A hold243/A hold252/A vssd1 vssd1 vccd1 vccd1 _10899_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18213_ _18212_/A _18212_/B _18212_/C vssd1 vssd1 vccd1 vccd1 _18215_/C sky130_fd_sc_hd__a21o_1
X_15425_ _15422_/X _15423_/Y _15283_/Y _15285_/Y vssd1 vssd1 vccd1 vccd1 _15426_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19193_ _19194_/B vssd1 vssd1 vccd1 vccd1 _19193_/Y sky130_fd_sc_hd__inv_2
X_12637_ _12637_/A _12637_/B _13152_/C _13152_/D vssd1 vssd1 vccd1 vccd1 _12639_/C
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18144_ _18144_/A _18144_/B vssd1 vssd1 vccd1 vccd1 _18152_/A sky130_fd_sc_hd__nand2_2
XANTENNA__15309__B2 _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15356_ _15492_/B _15356_/B vssd1 vssd1 vccd1 vccd1 _15356_/X sky130_fd_sc_hd__xor2_4
XFILLER_0_81_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12568_ _12567_/B _12567_/C _12567_/A vssd1 vssd1 vccd1 vccd1 _12570_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_81_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14307_ _16084_/C _14306_/X _14305_/X vssd1 vssd1 vccd1 vccd1 _14309_/A sky130_fd_sc_hd__a21bo_2
X_11519_ _21723_/D t1y[23] t0x[23] _11223_/A vssd1 vssd1 vccd1 vccd1 _11519_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18075_ _18074_/A _18074_/B _18074_/C vssd1 vssd1 vccd1 vccd1 _18077_/C sky130_fd_sc_hd__a21o_1
X_15287_ _15288_/A _15288_/B vssd1 vssd1 vccd1 vccd1 _15287_/Y sky130_fd_sc_hd__nand2b_2
XFILLER_0_41_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12499_ _12296_/X _12497_/Y _12498_/Y vssd1 vssd1 vccd1 vccd1 _12600_/A sky130_fd_sc_hd__a21o_2
Xhold207 hold207/A vssd1 vssd1 vccd1 vccd1 hold207/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold218 hold218/A vssd1 vssd1 vccd1 vccd1 hold218/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17026_ _17025_/B _17025_/C _17025_/A vssd1 vssd1 vccd1 vccd1 _17028_/C sky130_fd_sc_hd__a21bo_1
Xhold229 hold229/A vssd1 vssd1 vccd1 vccd1 hold229/X sky130_fd_sc_hd__dlygate4sd3_1
X_14238_ _14237_/B _14403_/B _14237_/A vssd1 vssd1 vccd1 vccd1 _14239_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_106_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1162 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14169_ _14301_/B _14168_/B _14303_/A _14168_/D vssd1 vssd1 vccd1 vccd1 _14170_/B
+ sky130_fd_sc_hd__o22a_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18977_ _18813_/B _18813_/Y _18974_/X _18976_/Y vssd1 vssd1 vccd1 vccd1 _18979_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17928_ _17928_/A _17928_/B vssd1 vssd1 vccd1 vccd1 _17937_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__12846__A2 _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18431__B1 _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17859_ _17980_/B _17859_/B vssd1 vssd1 vccd1 vccd1 _17869_/A sky130_fd_sc_hd__or2_1
XANTENNA__19181__B _19181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20870_ _20872_/A _20872_/B _20872_/C vssd1 vssd1 vccd1 vccd1 _20870_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19529_ _19686_/B _19529_/B _20265_/D vssd1 vssd1 vccd1 vccd1 _19529_/X sky130_fd_sc_hd__and3_1
XFILLER_0_53_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout159_A _16743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11282__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16745__B1 _17013_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20541__A1 _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20541__B2 _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20774__C _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16326__A _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout326_A hold319/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21422_ _21422_/A sstream_o sstream_i[114] vssd1 vssd1 vccd1 vccd1 _21422_/X sky130_fd_sc_hd__and3_1
XANTENNA__11034__A1 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_998 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16045__B _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21353_ _21412_/A _17970_/X _21421_/S _21352_/Y vssd1 vssd1 vccd1 vccd1 _21353_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20847__A2_N _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20304_ _20123_/Y _20162_/Y _20302_/Y _20303_/X vssd1 vssd1 vccd1 vccd1 _20355_/C
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_142_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout1 fanout2/X vssd1 vssd1 vccd1 vccd1 fanout1/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21284_ _21226_/A _21225_/B _21225_/A vssd1 vssd1 vccd1 vccd1 _21285_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1079 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20235_ _20235_/A _20235_/B vssd1 vssd1 vccd1 vccd1 _20236_/B sky130_fd_sc_hd__and2_1
X_20166_ _20166_/A _20166_/B vssd1 vssd1 vccd1 vccd1 _20212_/A sky130_fd_sc_hd__xnor2_2
X_20097_ _20097_/A _20097_/B vssd1 vssd1 vccd1 vccd1 _20121_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__17225__A1 _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17225__B2 _17417_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15787__A1 _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11870_ _11870_/A _11870_/B _11870_/C vssd1 vssd1 vccd1 vccd1 _11870_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_54_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10821_ _10821_/A _10821_/B vssd1 vssd1 vccd1 vccd1 _11053_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_39_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20999_ _20999_/A _20999_/B _20999_/C vssd1 vssd1 vccd1 vccd1 _20999_/X sky130_fd_sc_hd__and3_1
XFILLER_0_138_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11144__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13540_ _13383_/X _13385_/Y _13538_/A _13539_/X vssd1 vssd1 vccd1 vccd1 _13540_/Y
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__11273__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17977__D _19199_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__21142__A _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13471_ _13471_/A _13471_/B vssd1 vssd1 vccd1 vccd1 _13480_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_94_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12186__D _12246_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14211__A1 _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13014__A2 _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_943 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14211__B2 _14384_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11025__A1 hold256/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15210_ fanout9/X _15210_/B vssd1 vssd1 vccd1 vccd1 _15210_/Y sky130_fd_sc_hd__nor2_1
X_12422_ _12639_/A _12319_/C _12420_/D _12530_/A vssd1 vssd1 vccd1 vccd1 _12423_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16190_ _16303_/B _16191_/C _16191_/A vssd1 vssd1 vccd1 vccd1 _16193_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_35_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11576__A2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15141_ _15253_/A _15140_/C _15140_/A vssd1 vssd1 vccd1 vccd1 _15141_/X sky130_fd_sc_hd__a21o_1
X_12353_ _13155_/B _13157_/A _12780_/A _12780_/B vssd1 vssd1 vccd1 vccd1 _12354_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_129_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11304_ _13258_/D _11303_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21777_/D sky130_fd_sc_hd__mux2_1
X_15072_ hold205/X _15071_/X fanout4/A vssd1 vssd1 vccd1 vccd1 _21874_/D sky130_fd_sc_hd__mux2_1
X_12284_ _12130_/Y _12283_/X _12129_/Y vssd1 vssd1 vccd1 vccd1 _12284_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_22_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14023_ _14508_/A _14813_/A _15808_/C _14817_/C vssd1 vssd1 vccd1 vccd1 _14023_/X
+ sky130_fd_sc_hd__and4_1
X_18900_ _19373_/B _19057_/D _18901_/C _18901_/D vssd1 vssd1 vccd1 vccd1 _18900_/X
+ sky130_fd_sc_hd__and4_1
X_11235_ fanout59/X v0z[2] fanout19/X _11234_/X vssd1 vssd1 vccd1 vccd1 _11235_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19880_ _19879_/B _19879_/C _19879_/A vssd1 vssd1 vccd1 vccd1 _19880_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18831_ _18830_/B _18830_/C _18830_/A vssd1 vssd1 vccd1 vccd1 _18833_/C sky130_fd_sc_hd__o21a_1
XFILLER_0_105_1180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11166_ hold254/X _11126_/A fanout47/X hold312/X vssd1 vssd1 vccd1 vccd1 _11166_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18762_ _18604_/Y _18607_/X _18760_/Y _18761_/X vssd1 vssd1 vccd1 vccd1 _18822_/A
+ sky130_fd_sc_hd__o211a_1
X_15974_ _16305_/B _16396_/B _16418_/B _16196_/B vssd1 vssd1 vccd1 vccd1 _15978_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11097_ _11059_/Y hold19/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21691_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12004__A _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17713_ _17830_/B _17705_/X _17837_/A _17710_/B vssd1 vssd1 vccd1 vccd1 _17832_/A
+ sky130_fd_sc_hd__o22a_2
X_14925_ _14925_/A _14925_/B vssd1 vssd1 vccd1 vccd1 _14970_/A sky130_fd_sc_hd__nor2_1
X_18693_ _18693_/A _18693_/B vssd1 vssd1 vccd1 vccd1 _18830_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_26_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17767__A2 _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold90 hold90/A vssd1 vssd1 vccd1 vccd1 hold90/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11843__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14857__C _21755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17644_ _18319_/B _17642_/X _17643_/X vssd1 vssd1 vccd1 vccd1 _17645_/B sky130_fd_sc_hd__a21bo_1
X_14856_ _14557_/B _21755_/Q _16380_/B _12771_/C vssd1 vssd1 vccd1 vccd1 _14859_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__20771__A1 _11550_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20771__B2 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13807_ _13804_/X _13805_/X _13652_/C _13652_/Y vssd1 vssd1 vccd1 vccd1 _13807_/Y
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__11562__B _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15034__B _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17575_ _17575_/A _17575_/B _17575_/C _17575_/D vssd1 vssd1 vccd1 vccd1 _17575_/X
+ sky130_fd_sc_hd__or4_2
X_14787_ _15702_/D _15717_/C _15976_/D _15579_/D vssd1 vssd1 vccd1 vccd1 _14790_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13253__A2 _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14450__A1 _21725_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11054__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11999_ _11999_/A _11999_/B _11999_/C vssd1 vssd1 vccd1 vccd1 _12011_/A sky130_fd_sc_hd__nand3_2
XANTENNA__14450__B2 fanout6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19314_ _19152_/A _19152_/C _19152_/B vssd1 vssd1 vccd1 vccd1 _19316_/B sky130_fd_sc_hd__a21boi_1
X_16526_ _16525_/A _16525_/B _16525_/C vssd1 vssd1 vccd1 vccd1 _16532_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_46_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13738_ _13581_/A _13581_/Y _13736_/Y _13737_/X vssd1 vssd1 vccd1 vccd1 _13800_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_85_364 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14873__B _14873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19245_ _19073_/A _19073_/C _19073_/B vssd1 vssd1 vccd1 vccd1 _19246_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_129_989 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16457_ _16703_/A _16703_/B vssd1 vssd1 vccd1 vccd1 _16493_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13669_ _13669_/A _13669_/B vssd1 vssd1 vccd1 vccd1 _13702_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_42_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12674__A _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15408_ _15931_/B _16396_/A _16266_/C _15931_/A vssd1 vssd1 vccd1 vccd1 _15412_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18064__C _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19176_ _19176_/A _19176_/B vssd1 vssd1 vccd1 vccd1 _19218_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_147_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16388_ _16388_/A _16388_/B vssd1 vssd1 vccd1 vccd1 _16390_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18127_ _18121_/B _18127_/B _18127_/C vssd1 vssd1 vccd1 vccd1 _18129_/B sky130_fd_sc_hd__and3b_1
X_15339_ _15338_/B _15338_/C _15338_/A vssd1 vssd1 vccd1 vccd1 _15340_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18058_ _18058_/A _19703_/C vssd1 vssd1 vccd1 vccd1 _18062_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17009_ _17002_/A _17002_/C _17002_/B vssd1 vssd1 vccd1 vccd1 _17009_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_1_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout506 _21743_/Q vssd1 vssd1 vccd1 vccd1 _16374_/A sky130_fd_sc_hd__buf_4
X_20020_ _19985_/Y _20164_/A _20168_/B _20020_/D vssd1 vssd1 vccd1 vccd1 _20164_/B
+ sky130_fd_sc_hd__and4bb_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout517 _21740_/Q vssd1 vssd1 vccd1 vccd1 _13875_/B sky130_fd_sc_hd__buf_4
Xfanout528 _14659_/A vssd1 vssd1 vccd1 vccd1 _15702_/D sky130_fd_sc_hd__buf_4
XFILLER_0_10_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout539 _21736_/Q vssd1 vssd1 vccd1 vccd1 _15439_/D sky130_fd_sc_hd__buf_4
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21971_ _21974_/CLK _21971_/D vssd1 vssd1 vccd1 vccd1 hold302/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_83_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_32_clk_i clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _22105_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_154_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout276_A _18008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20922_ _21151_/A _21301_/A _21305_/A _21153_/B vssd1 vssd1 vccd1 vccd1 _21097_/A
+ sky130_fd_sc_hd__nand4_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13671__C _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20853_ _20853_/A vssd1 vssd1 vccd1 vccd1 _20855_/B sky130_fd_sc_hd__inv_2
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11255__A1 fanout59/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20784_ _20784_/A _20784_/B vssd1 vssd1 vccd1 vccd1 _20786_/B sky130_fd_sc_hd__and2_1
XFILLER_0_77_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_1240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout610_A _21718_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21405_ _21720_/D _20645_/X _21421_/S _21404_/Y vssd1 vssd1 vccd1 vccd1 _21405_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__15895__A _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18271__A _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_968 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21336_ hold132/X _21381_/B _21334_/Y _21335_/Y vssd1 vssd1 vccd1 vccd1 _21919_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18891__B1 _19051_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13704__B1 _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21267_ _21267_/A hold294/A vssd1 vssd1 vccd1 vccd1 _21269_/A sky130_fd_sc_hd__nand2_1
XANTENNA_fanout91_A _21844_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11020_ mstream_o[94] hold46/X _11027_/S vssd1 vssd1 vccd1 vccd1 _21631_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_25_1163 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20218_ _20218_/A _20218_/B vssd1 vssd1 vccd1 vccd1 _20220_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__11647__B _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21198_ _21199_/A _21293_/B _21853_/Q _21199_/B vssd1 vssd1 vccd1 vccd1 _21200_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_2_0__f_clk_i_A clkbuf_0_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14023__B _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20149_ _20149_/A _20281_/B vssd1 vssd1 vccd1 vccd1 _20151_/B sky130_fd_sc_hd__or2_1
XTAP_3400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12971_ _12971_/A _12971_/B _12971_/C vssd1 vssd1 vccd1 vccd1 _12972_/B sky130_fd_sc_hd__and3_1
XANTENNA__17334__B _17334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14710_ _14690_/A _14690_/B _14709_/A _14709_/B vssd1 vssd1 vccd1 vccd1 _14710_/Y
+ sky130_fd_sc_hd__a211oi_2
XTAP_3444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11494__A1 _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11922_ _11922_/A _11922_/B vssd1 vssd1 vccd1 vccd1 _11923_/B sky130_fd_sc_hd__nor2_1
X_15690_ _15689_/B _15689_/C _15689_/A vssd1 vssd1 vccd1 vccd1 _15690_/X sky130_fd_sc_hd__o21a_1
XTAP_3455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14641_ _14640_/B _14640_/C _14640_/A vssd1 vssd1 vccd1 vccd1 _14642_/C sky130_fd_sc_hd__a21o_1
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11853_ _11853_/A _11853_/B vssd1 vssd1 vccd1 vccd1 _11854_/C sky130_fd_sc_hd__xor2_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_1150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10804_ hold88/A hold34/A vssd1 vssd1 vccd1 vccd1 _10807_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11246__A1 _11549_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17360_ _17382_/B _17360_/B _17360_/C _17360_/D vssd1 vssd1 vccd1 vccd1 _17362_/A
+ sky130_fd_sc_hd__nor4_2
X_14572_ _14572_/A _14572_/B vssd1 vssd1 vccd1 vccd1 _14974_/A sky130_fd_sc_hd__and2_2
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11246__B2 _21724_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11784_ _11784_/A _11784_/B _11784_/C vssd1 vssd1 vccd1 vccd1 _11788_/A sky130_fd_sc_hd__nand3_1
XANTENNA__14693__B _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16311_ _16310_/B _16311_/B vssd1 vssd1 vccd1 vccd1 _16312_/B sky130_fd_sc_hd__and2b_1
XANTENNA__12994__A1 _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13523_ _13523_/A _13523_/B vssd1 vssd1 vccd1 vccd1 _13656_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_32_1156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17291_ _17188_/A _17188_/B _17186_/X vssd1 vssd1 vccd1 vccd1 _17293_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_126_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19030_ _20032_/D _19810_/D _19030_/C _21847_/Q vssd1 vssd1 vccd1 vccd1 _19032_/D
+ sky130_fd_sc_hd__nand4_1
X_16242_ _16128_/A _16128_/Y _16347_/B _16241_/X vssd1 vssd1 vccd1 vccd1 _16352_/A
+ sky130_fd_sc_hd__a211o_1
X_13454_ _13450_/X _13451_/Y _13299_/X _13301_/X vssd1 vssd1 vccd1 vccd1 _13491_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_152_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20269__B1 _20924_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12405_ _12403_/X _12405_/B vssd1 vssd1 vccd1 vccd1 _12406_/B sky130_fd_sc_hd__and2b_1
X_16173_ _16173_/A _16173_/B vssd1 vssd1 vccd1 vccd1 _16284_/B sky130_fd_sc_hd__and2_1
X_13385_ _13386_/A _13386_/B vssd1 vssd1 vccd1 vccd1 _13385_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_134_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15124_ _15328_/A _15124_/B vssd1 vssd1 vccd1 vccd1 _15126_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_133_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20861__D _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12336_ _12336_/A _12336_/B _12336_/C vssd1 vssd1 vccd1 vccd1 _12338_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_107_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15055_ _15055_/A _15055_/B vssd1 vssd1 vccd1 vccd1 _15056_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12267_ _12267_/A _12269_/D _12267_/C _12267_/D vssd1 vssd1 vccd1 vccd1 _12267_/Y
+ sky130_fd_sc_hd__nand4_1
X_19932_ _19932_/A _19932_/B vssd1 vssd1 vccd1 vccd1 _19934_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14214__A _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13171__A1 _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12660__C _21765_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14006_ _13842_/A _13843_/Y _14004_/X _14005_/Y vssd1 vssd1 vccd1 vccd1 _14007_/A
+ sky130_fd_sc_hd__a211oi_2
X_11218_ hold201/X fanout22/X _11217_/X vssd1 vssd1 vccd1 vccd1 _11218_/X sky130_fd_sc_hd__a21o_1
XANTENNA__13171__B2 _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19863_ _19863_/A _19863_/B _19863_/C vssd1 vssd1 vccd1 vccd1 _19885_/B sky130_fd_sc_hd__and3_2
XFILLER_0_128_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12198_ _12199_/A _12199_/B _12199_/C vssd1 vssd1 vccd1 vccd1 _12207_/A sky130_fd_sc_hd__o21ai_2
XANTENNA__11049__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17525__A _17525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18814_ _18813_/B _18813_/C _18813_/A vssd1 vssd1 vccd1 vccd1 _18814_/Y sky130_fd_sc_hd__a21oi_1
X_11149_ hold182/X fanout23/X _11148_/X vssd1 vssd1 vccd1 vccd1 _11149_/X sky130_fd_sc_hd__a21o_1
X_19794_ hold174/A fanout8/X _14918_/Y _11550_/B _19793_/Y vssd1 vssd1 vccd1 vccd1
+ _19794_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18745_ _18745_/A _18745_/B vssd1 vssd1 vccd1 vccd1 _18758_/A sky130_fd_sc_hd__xnor2_1
X_15957_ _16092_/D _21787_/Q _15957_/C _15957_/D vssd1 vssd1 vccd1 vccd1 _16089_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_37_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12669__A _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13474__A2 _15370_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14908_ _14909_/A _14909_/B vssd1 vssd1 vccd1 vccd1 _14910_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11485__A1 _18624_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18059__C _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18676_ _18521_/C _18520_/Y _18674_/X _18675_/Y vssd1 vssd1 vccd1 vccd1 _18676_/Y
+ sky130_fd_sc_hd__o211ai_2
X_15888_ _15888_/A _15888_/B vssd1 vssd1 vccd1 vccd1 _15888_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_53_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17627_ _17627_/A _17627_/B vssd1 vssd1 vccd1 vccd1 _17629_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__20101__D _21817_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14839_ _14840_/A _14840_/B _14840_/C vssd1 vssd1 vccd1 vccd1 _14839_/X sky130_fd_sc_hd__and3_1
XANTENNA__11237__A1 _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11237__B2 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17558_ _19123_/B _17670_/B _20270_/C _19123_/A vssd1 vssd1 vccd1 vccd1 _17559_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18165__A2 _18929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16509_ _16507_/X _16508_/Y _17096_/A _16860_/C vssd1 vssd1 vccd1 vccd1 _16668_/A
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_156_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17489_ _17489_/A _17489_/B vssd1 vssd1 vccd1 vccd1 _17584_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_46_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11512__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19228_ _19230_/A _19382_/B _19230_/C _19230_/D vssd1 vssd1 vccd1 vccd1 _19228_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13012__B _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19159_ _19159_/A _19159_/B vssd1 vssd1 vccd1 vccd1 _19162_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_54_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17125__B1 _17141_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_1190 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19665__A2 _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21121_ _21236_/A _21119_/X _21003_/Y _21005_/X vssd1 vssd1 vccd1 vccd1 _21122_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA__19337__D _19337_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21052_ _21052_/A _21052_/B vssd1 vssd1 vccd1 vccd1 _21053_/B sky130_fd_sc_hd__nand2_1
Xfanout303 _17086_/C vssd1 vssd1 vccd1 vccd1 _17019_/C sky130_fd_sc_hd__buf_4
XFILLER_0_10_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout314 _21792_/Q vssd1 vssd1 vccd1 vccd1 _17141_/C sky130_fd_sc_hd__clkbuf_4
Xfanout325 _21790_/Q vssd1 vssd1 vccd1 vccd1 _18859_/A sky130_fd_sc_hd__buf_6
XANTENNA_fanout393_A _15892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout336 _21785_/Q vssd1 vssd1 vccd1 vccd1 _16399_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_10_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11712__A2 _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20003_ _20562_/B _20924_/A _19868_/B _20689_/A vssd1 vssd1 vccd1 vccd1 _20003_/Y
+ sky130_fd_sc_hd__a22oi_1
Xfanout347 _21782_/Q vssd1 vssd1 vccd1 vccd1 _16396_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__16977__C _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout358 _16391_/A vssd1 vssd1 vccd1 vccd1 _15911_/A sky130_fd_sc_hd__buf_2
Xfanout369 _21777_/Q vssd1 vssd1 vccd1 vccd1 _15916_/B sky130_fd_sc_hd__buf_2
XFILLER_0_94_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout560_A _21731_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18928__A1 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18928__B2 _21833_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11476__A1 _18789_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19050__B1 _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21954_ _21963_/CLK _21954_/D vssd1 vssd1 vccd1 vccd1 hold249/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__19196__A4 _21847_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21391__S _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17600__A1 _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20905_ _20904_/A _20904_/B _20904_/C _20904_/D _20899_/Y vssd1 vssd1 vccd1 vccd1
+ _21026_/B sky130_fd_sc_hd__a41oi_4
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21885_ _21945_/CLK _21885_/D vssd1 vssd1 vccd1 vccd1 hold232/A sky130_fd_sc_hd__dfxtp_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11228__A1 _11227_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20836_ _20836_/A _20836_/B vssd1 vssd1 vccd1 vccd1 _20881_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11930__B _12897_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20767_ _20903_/A _20904_/A vssd1 vssd1 vccd1 vccd1 _20900_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_65_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11422__S _11446_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_518 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20698_ _20698_/A _20698_/B _20698_/C vssd1 vssd1 vccd1 vccd1 _20699_/C sky130_fd_sc_hd__nand3_1
XANTENNA__14018__B _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18713__B _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13170_ _13047_/A _13046_/B _13046_/A vssd1 vssd1 vccd1 vccd1 _13177_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__18432__C _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ _12127_/A _12121_/B vssd1 vssd1 vccd1 vccd1 _12124_/B sky130_fd_sc_hd__nand2_1
X_21319_ _21319_/A _21319_/B vssd1 vssd1 vccd1 vccd1 _21320_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__11951__A2 _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11658__A _12402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19825__A _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19408__A2 _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12052_ _11996_/A _11996_/C _11996_/B vssd1 vssd1 vccd1 vccd1 _12053_/C sky130_fd_sc_hd__a21o_1
XANTENNA__13295__D _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11003_ mstream_o[77] hold99/X _11005_/S vssd1 vssd1 vccd1 vccd1 _21614_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12900__A1 _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16860_ _17141_/A _17141_/B _16860_/C _16917_/C vssd1 vssd1 vccd1 vccd1 _16863_/A
+ sky130_fd_sc_hd__nand4_1
X_15811_ _15811_/A _15811_/B vssd1 vssd1 vccd1 vccd1 _15813_/B sky130_fd_sc_hd__xor2_1
XANTENNA__17064__B _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16791_ _16792_/A _16792_/B vssd1 vssd1 vccd1 vccd1 _17379_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13456__A2 _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15850__B1 _16418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18530_ _18529_/B _18529_/C _18529_/A vssd1 vssd1 vccd1 vccd1 _18530_/Y sky130_fd_sc_hd__o21ai_2
X_15742_ _15741_/A _15741_/B _15741_/C _15741_/D vssd1 vssd1 vccd1 vccd1 _15742_/Y
+ sky130_fd_sc_hd__o22ai_4
XTAP_3230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11467__A1 _18058_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12954_ _21725_/D hold96/X _11057_/Y fanout6/X _12953_/Y vssd1 vssd1 vccd1 vccd1
+ _12954_/X sky130_fd_sc_hd__a221o_1
XTAP_3252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18461_ _19695_/A _18929_/B _18616_/D _19686_/A vssd1 vssd1 vccd1 vccd1 _18464_/C
+ sky130_fd_sc_hd__a22o_1
X_11905_ _11905_/A _11905_/B _11900_/A vssd1 vssd1 vccd1 vccd1 _11905_/Y sky130_fd_sc_hd__nor3b_2
X_15673_ _15931_/A _15931_/B _16414_/B _16391_/B vssd1 vssd1 vccd1 vccd1 _15802_/A
+ sky130_fd_sc_hd__and4_1
XTAP_3285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14405__A1 _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_230 hold290/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ _12884_/B _12884_/C _12884_/A vssd1 vssd1 vccd1 vccd1 _12887_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14405__B2 _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_241 hold309/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17412_ _17520_/B _20774_/A _20774_/B _17619_/A vssd1 vssd1 vccd1 vccd1 _17413_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA_252 v0z[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_263 hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14624_ _14624_/A _14624_/B vssd1 vssd1 vccd1 vccd1 _14625_/B sky130_fd_sc_hd__nor2_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18392_ hold136/A fanout8/X _18390_/Y _11550_/A _18391_/Y vssd1 vssd1 vccd1 vccd1
+ _18392_/X sky130_fd_sc_hd__a221o_1
X_11836_ _11836_/A _11836_/B _11836_/C vssd1 vssd1 vccd1 vccd1 _11836_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_56_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_274 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_285 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18147__A2 _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_296 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17343_ _17343_/A _17343_/B _17343_/C vssd1 vssd1 vccd1 vccd1 _17345_/B sky130_fd_sc_hd__nand3_1
X_14555_ _14848_/A _14557_/D _14413_/X _14242_/X _14250_/B vssd1 vssd1 vccd1 vccd1
+ _14560_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_126_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _11767_/A _11767_/B _11767_/C vssd1 vssd1 vccd1 vccd1 _11772_/A sky130_fd_sc_hd__nand3_4
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11332__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22092__RESET_B _11089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13506_ _13248_/Y _13251_/Y _13503_/Y _13505_/X vssd1 vssd1 vccd1 vccd1 _13508_/A
+ sky130_fd_sc_hd__a211o_1
X_17274_ hold223/X _17273_/X fanout3/X vssd1 vssd1 vccd1 vccd1 _21887_/D sky130_fd_sc_hd__mux2_1
X_14486_ _14331_/B _14333_/B _14647_/A _14485_/Y vssd1 vssd1 vccd1 vccd1 _14647_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_83_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11698_ _12330_/B _11697_/B _11697_/C vssd1 vssd1 vccd1 vccd1 _11699_/C sky130_fd_sc_hd__a21o_1
X_19013_ _19493_/D _19337_/D _19013_/C vssd1 vssd1 vccd1 vccd1 _19013_/X sky130_fd_sc_hd__and3_1
XFILLER_0_153_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16225_ _16226_/A _16226_/B _16226_/C vssd1 vssd1 vccd1 vccd1 _16225_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_113_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13437_ _14024_/B _14537_/A _13437_/C _13437_/D vssd1 vssd1 vccd1 vccd1 _13439_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_10_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19438__C _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17658__A1 _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16156_ _16418_/A _16377_/A _16157_/C _16157_/D vssd1 vssd1 vccd1 vccd1 _16158_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__17658__B2 _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13368_ _13518_/C _13368_/B vssd1 vssd1 vccd1 vccd1 _13369_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_24_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15107_ _15108_/A _15108_/B _15254_/B _15108_/D vssd1 vssd1 vccd1 vccd1 _15107_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_122_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11568__A _12229_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12319_ _13554_/B _14621_/D _12319_/C _12420_/D vssd1 vssd1 vccd1 vccd1 _12401_/A
+ sky130_fd_sc_hd__and4_1
X_16087_ _16087_/A _21787_/Q _16087_/C _16087_/D vssd1 vssd1 vccd1 vccd1 _16201_/B
+ sky130_fd_sc_hd__and4_1
X_13299_ _13300_/B _13300_/A vssd1 vssd1 vccd1 vccd1 _13299_/X sky130_fd_sc_hd__and2b_2
X_15038_ _15037_/B _15037_/C _15037_/A vssd1 vssd1 vccd1 vccd1 _15040_/B sky130_fd_sc_hd__a21o_1
X_19915_ _19917_/B vssd1 vssd1 vccd1 vccd1 _19915_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_43_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19846_ _19847_/A _19847_/B vssd1 vssd1 vccd1 vccd1 _20381_/A sky130_fd_sc_hd__nor2_2
XANTENNA__20965__A1 _21293_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20965__B2 _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16989_ _16990_/A _16988_/Y _16989_/C _17146_/D vssd1 vssd1 vccd1 vccd1 _17033_/A
+ sky130_fd_sc_hd__and4bb_1
X_19777_ _19777_/A _19777_/B vssd1 vssd1 vccd1 vccd1 _19779_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11458__A1 _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_927 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18728_ _18847_/B _18726_/X _18610_/Y _18613_/Y vssd1 vssd1 vccd1 vccd1 _18728_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18659_ _18658_/B _18658_/C _18658_/A vssd1 vssd1 vccd1 vccd1 _18661_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_8_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15503__A _15907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21670_ _21939_/CLK _21670_/D vssd1 vssd1 vccd1 vccd1 hold70/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__14947__A2 _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18138__A2 _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20621_ _20621_/A _20621_/B _20621_/C vssd1 vssd1 vccd1 vccd1 _20621_/Y sky130_fd_sc_hd__nor3_2
XANTENNA_fanout141_A _20249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout239_A _17915_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12565__C _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20552_ _20552_/A _20552_/B vssd1 vssd1 vccd1 vccd1 _20554_/B sky130_fd_sc_hd__or2_1
XFILLER_0_144_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20483_ _20483_/A _20483_/B vssd1 vssd1 vccd1 vccd1 _20484_/B sky130_fd_sc_hd__or2_1
XANTENNA_fanout406_A _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21104_ _21105_/B _21105_/A vssd1 vssd1 vccd1 vccd1 _21222_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_22_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15892__B _15892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_22084_ _22096_/CLK _22084_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[20] sky130_fd_sc_hd__dfrtp_4
XANTENNA__20006__D _21286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout100 _20419_/A vssd1 vssd1 vccd1 vccd1 _19060_/B sky130_fd_sc_hd__buf_4
XFILLER_0_100_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout111 _21267_/A vssd1 vssd1 vccd1 vccd1 _19692_/C sky130_fd_sc_hd__clkbuf_4
Xfanout122 _21056_/A vssd1 vssd1 vccd1 vccd1 _17739_/C sky130_fd_sc_hd__buf_4
X_21035_ _21035_/A _21035_/B vssd1 vssd1 vccd1 vccd1 _21075_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_10_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout133 _19087_/B vssd1 vssd1 vccd1 vccd1 _18616_/D sky130_fd_sc_hd__clkbuf_8
Xfanout144 _21833_/Q vssd1 vssd1 vccd1 vccd1 _18624_/A sky130_fd_sc_hd__clkbuf_8
Xfanout155 _21830_/Q vssd1 vssd1 vccd1 vccd1 _16989_/C sky130_fd_sc_hd__clkbuf_8
Xfanout166 _21828_/Q vssd1 vssd1 vccd1 vccd1 _16813_/A sky130_fd_sc_hd__clkbuf_4
Xfanout177 _21826_/Q vssd1 vssd1 vccd1 vccd1 _16734_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__16500__C _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout188 _17146_/B vssd1 vssd1 vccd1 vccd1 _17141_/B sky130_fd_sc_hd__buf_4
XFILLER_0_57_1207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout199 _21256_/B vssd1 vssd1 vccd1 vccd1 _20242_/D sky130_fd_sc_hd__buf_4
XANTENNA__13438__A2 _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11449__A1 _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout54_A _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21415__A _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21937_ _21942_/CLK _21937_/D vssd1 vssd1 vccd1 vccd1 hold174/A sky130_fd_sc_hd__dfxtp_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14399__B1 _14398_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18427__C _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ _12668_/Y _12669_/X _13155_/A _12781_/D vssd1 vssd1 vccd1 vccd1 _12672_/A
+ sky130_fd_sc_hd__and4bb_1
X_21868_ _21942_/CLK hold141/X vssd1 vssd1 vccd1 vccd1 hold140/A sky130_fd_sc_hd__dfxtp_1
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14674__D _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _12316_/A _11621_/B vssd1 vssd1 vccd1 vccd1 _11623_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20819_ _20819_/A _20819_/B vssd1 vssd1 vccd1 vccd1 _20820_/B sky130_fd_sc_hd__or2_1
XANTENNA__18146__D _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21799_ _21803_/CLK _21799_/D vssd1 vssd1 vccd1 vccd1 _21799_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__13610__A2 _14218_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14340_ _14340_/A _14340_/B vssd1 vssd1 vccd1 vccd1 _14341_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_53_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11552_ _21412_/A _11551_/Y _21329_/B1 vssd1 vssd1 vccd1 vccd1 fanout4/A sky130_fd_sc_hd__o21a_4
XFILLER_0_135_542 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14271_ _14107_/X _14109_/X _14268_/X _14269_/Y vssd1 vssd1 vccd1 vccd1 _14273_/B
+ sky130_fd_sc_hd__a211o_1
X_11483_ _11498_/A1 t1y[11] t0x[11] _11501_/B2 vssd1 vssd1 vccd1 vccd1 _11483_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_52_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16010_ _16010_/A _16010_/B vssd1 vssd1 vccd1 vccd1 _16014_/A sky130_fd_sc_hd__xnor2_1
X_13222_ _13361_/A _13222_/B vssd1 vssd1 vccd1 vccd1 _13365_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_61_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13153_ _13153_/A _13153_/B vssd1 vssd1 vccd1 vccd1 _13154_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12104_ _12104_/A _12104_/B vssd1 vssd1 vccd1 vccd1 _12106_/B sky130_fd_sc_hd__xnor2_1
X_13084_ _13083_/B _13083_/C _13083_/A vssd1 vssd1 vccd1 vccd1 _13085_/B sky130_fd_sc_hd__o21a_1
X_17961_ _17958_/X _17959_/Y _17819_/B _17821_/A vssd1 vssd1 vccd1 vccd1 _17962_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16912_ _16912_/A _16912_/B vssd1 vssd1 vccd1 vccd1 _16912_/Y sky130_fd_sc_hd__nand2_1
X_12035_ _12035_/A _12035_/B vssd1 vssd1 vccd1 vccd1 _12289_/A sky130_fd_sc_hd__xnor2_4
X_19700_ _19700_/A _19700_/B vssd1 vssd1 vccd1 vccd1 _19708_/A sky130_fd_sc_hd__nand2_1
X_17892_ _17785_/A _17784_/B _17782_/X vssd1 vssd1 vccd1 vccd1 _17908_/A sky130_fd_sc_hd__a21o_1
XANTENNA__19801__A2 _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16843_ _16844_/A _16844_/B _16849_/C _16844_/D vssd1 vssd1 vccd1 vccd1 _16843_/Y
+ sky130_fd_sc_hd__nor4_1
X_19631_ _19631_/A _19631_/B vssd1 vssd1 vccd1 vccd1 _19634_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_137_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19562_ _19562_/A _19562_/B vssd1 vssd1 vccd1 vccd1 _19617_/A sky130_fd_sc_hd__nor2_1
X_16774_ _16764_/X _16770_/X _16783_/A _16773_/Y vssd1 vssd1 vccd1 vccd1 _16783_/B
+ sky130_fd_sc_hd__o211ai_2
X_13986_ _13986_/A _13986_/B vssd1 vssd1 vccd1 vccd1 _13987_/A sky130_fd_sc_hd__or2_1
XFILLER_0_137_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18513_ _18363_/B _18363_/Y _18510_/X _18512_/Y vssd1 vssd1 vccd1 vccd1 _18516_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_38_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19565__A1 _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15725_ _15727_/A _15727_/B _15727_/C vssd1 vssd1 vccd1 vccd1 _15725_/Y sky130_fd_sc_hd__a21oi_1
XTAP_3060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19565__B2 _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17522__B _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19493_ _18849_/B _20178_/B _20721_/C _19493_/D vssd1 vssd1 vccd1 vccd1 _19496_/A
+ sky130_fd_sc_hd__and4b_2
X_12937_ _12934_/X _12935_/Y _12807_/C _12808_/X vssd1 vssd1 vccd1 vccd1 _12938_/C
+ sky130_fd_sc_hd__o211ai_4
XTAP_3071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18444_ _19529_/B _19531_/A _19068_/C _19238_/C vssd1 vssd1 vccd1 vccd1 _18594_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_75_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15656_ _15656_/A _15849_/B vssd1 vssd1 vccd1 vccd1 _15667_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14929__A2 _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12868_ _12868_/A _12868_/B _12868_/C vssd1 vssd1 vccd1 vccd1 _12869_/C sky130_fd_sc_hd__nand3_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14607_ hold216/X _14606_/X fanout4/X vssd1 vssd1 vccd1 vccd1 _21871_/D sky130_fd_sc_hd__mux2_1
X_18375_ _18225_/B _18224_/Y _18373_/X _18374_/Y vssd1 vssd1 vccd1 vccd1 _18377_/C
+ sky130_fd_sc_hd__o211ai_4
X_11819_ _11819_/A _11819_/B _11819_/C vssd1 vssd1 vccd1 vccd1 _11823_/A sky130_fd_sc_hd__nand3_4
X_15587_ _15587_/A _15587_/B vssd1 vssd1 vccd1 vccd1 _15598_/A sky130_fd_sc_hd__or2_1
XFILLER_0_84_952 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11062__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12799_ _12798_/B _12798_/C _12798_/A vssd1 vssd1 vccd1 vccd1 _12799_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_56_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17326_ _17324_/X _17326_/B vssd1 vssd1 vccd1 vccd1 _17327_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_56_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14538_ _14538_/A _14538_/B vssd1 vssd1 vccd1 vccd1 _14546_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21060__A _21171_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13778__A _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17257_ _17256_/A _17256_/B _17256_/C _17256_/D vssd1 vssd1 vccd1 vccd1 _17257_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_109_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14469_ _14469_/A _14469_/B vssd1 vssd1 vccd1 vccd1 _14471_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16154__A _16391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16208_ _16207_/A _16207_/B _16207_/C vssd1 vssd1 vccd1 vccd1 _16209_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17188_ _17188_/A _17188_/B vssd1 vssd1 vccd1 vccd1 _17191_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16139_ _16007_/A _16009_/X _16251_/B _16138_/X vssd1 vssd1 vccd1 vccd1 _16142_/A
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11729__C _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14314__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12340__A2 _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19829_ _19828_/B _19828_/C _19828_/A vssd1 vssd1 vccd1 vccd1 _19830_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_120_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13018__A _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout189_A _21823_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11300__A0 _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14774__A_N _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout356_A _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17031__A2 _17145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21722_ _21722_/CLK _21722_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[114]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__11851__A1 _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11851__B2 _12242_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21653_ _21888_/CLK _21653_/D vssd1 vssd1 vccd1 vccd1 hold72/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout523_A _13877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11911__D _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11603__A1 _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20604_ _20863_/C _21283_/B _21305_/B _21261_/A vssd1 vssd1 vccd1 vccd1 _20608_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11603__B2 _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21584_ _22106_/CLK _21584_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[47] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_90_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20535_ _20918_/A _20535_/B vssd1 vssd1 vccd1 vccd1 _20665_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_90_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16542__A1 _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20466_ _20466_/A _20466_/B _20466_/C vssd1 vssd1 vccd1 vccd1 _20468_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_120_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19375__A _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11639__C _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20397_ _20397_/A _20397_/B vssd1 vssd1 vccd1 vccd1 _20398_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14305__B1 _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17730__A1_N _18851_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11119__A0 _10978_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14856__A1 _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14856__B2 _12771_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16511__B _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22067_ _22069_/CLK _22067_/D fanout639/X vssd1 vssd1 vccd1 vccd1 mstream_o[3] sky130_fd_sc_hd__dfrtp_4
XANTENNA__20929__A1 _21842_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21018_ _21129_/A _21016_/Y _20880_/X _20882_/Y vssd1 vssd1 vccd1 vccd1 _21018_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13573__D _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11147__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13840_ _13707_/D _13708_/B _13838_/Y _13839_/X vssd1 vssd1 vccd1 vccd1 _13842_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_134_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19547__A1 _21839_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15455__A2_N _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13771_ _14848_/A _14077_/B vssd1 vssd1 vccd1 vccd1 _13775_/A sky130_fd_sc_hd__nand2_1
X_10983_ _10978_/A _10977_/A _10977_/B vssd1 vssd1 vccd1 vccd1 _10984_/B sky130_fd_sc_hd__a21bo_2
XANTENNA__17558__B1 _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_908 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15510_ _16027_/A _15510_/B _15510_/C _15670_/A vssd1 vssd1 vccd1 vccd1 _15670_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12722_ _13975_/B _13682_/C _13258_/C _13258_/D vssd1 vssd1 vccd1 vccd1 _12851_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_97_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16490_ _17636_/B _17387_/A _16489_/C _16489_/D vssd1 vssd1 vccd1 vccd1 _16491_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__15033__A1 _15933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15441_ _15439_/D _16406_/B _16374_/B _21735_/Q vssd1 vssd1 vccd1 vccd1 _15442_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_12653_ _12653_/A _12653_/B _12653_/C vssd1 vssd1 vccd1 vccd1 _12653_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_84_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18160_ _18157_/Y _18158_/X _18044_/B _18046_/A vssd1 vssd1 vccd1 vccd1 _18160_/Y
+ sky130_fd_sc_hd__o211ai_1
X_11604_ _12319_/C _12420_/D _12268_/B _12302_/A vssd1 vssd1 vccd1 vccd1 _11612_/A
+ sky130_fd_sc_hd__and4_1
X_15372_ _15373_/B _16286_/B _16027_/B _15373_/A vssd1 vssd1 vccd1 vccd1 _15374_/A
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_108_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12584_ _12583_/A _12583_/B _12583_/C _12583_/D vssd1 vssd1 vccd1 vccd1 _12584_/Y
+ sky130_fd_sc_hd__o22ai_4
XFILLER_0_37_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17111_ _17156_/C _17110_/X _17156_/A _17156_/B vssd1 vssd1 vccd1 vccd1 _17111_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_25_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14323_ _15159_/D _14936_/D _14155_/C _14155_/D _14157_/X vssd1 vssd1 vccd1 vccd1
+ _14331_/A sky130_fd_sc_hd__a41o_1
XFILLER_0_52_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18091_ _18091_/A _18091_/B _18091_/C vssd1 vssd1 vccd1 vccd1 _18091_/Y sky130_fd_sc_hd__nand3_4
X_11535_ _11544_/A1 t2x[28] v1z[28] fanout20/X _11534_/X vssd1 vssd1 vccd1 vccd1 _11535_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_151_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17042_ _17058_/A _17036_/B _17034_/Y vssd1 vssd1 vccd1 vccd1 _17044_/B sky130_fd_sc_hd__o21a_1
X_14254_ _14254_/A _14418_/A _14254_/C vssd1 vssd1 vccd1 vccd1 _14255_/C sky130_fd_sc_hd__or3_1
XFILLER_0_123_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11466_ _21718_/D t2x[5] v1z[5] fanout17/X _11465_/X vssd1 vssd1 vccd1 vccd1 _11466_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_68_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13748__D _14212_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18901__B _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13205_ _13204_/B _13204_/C _13204_/A vssd1 vssd1 vccd1 vccd1 _13205_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_0_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14185_ _14659_/A _15022_/B _14185_/C _14185_/D vssd1 vssd1 vccd1 vccd1 _14185_/Y
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_110_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11397_ hold304/X fanout28/X _11396_/X vssd1 vssd1 vccd1 vccd1 _11397_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_104_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13136_ _13136_/A _13136_/B _13136_/C vssd1 vssd1 vccd1 vccd1 _13140_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_104_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18993_ _18830_/B _18833_/B _19155_/B _18992_/Y vssd1 vssd1 vccd1 vccd1 _18995_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14847__A1 _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ _13067_/A _13067_/B _13067_/C vssd1 vssd1 vccd1 vccd1 _13067_/X sky130_fd_sc_hd__or3_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17944_ _17943_/B _17943_/C _17943_/A vssd1 vssd1 vccd1 vccd1 _17944_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__13764__C _14873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12018_ _12426_/B _12312_/A _11952_/C _11952_/D vssd1 vssd1 vccd1 vccd1 _12019_/B
+ sky130_fd_sc_hd__a22oi_1
X_17875_ _17874_/A _17741_/B _18006_/A _17874_/D vssd1 vssd1 vccd1 vccd1 _17876_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19732__B _19732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15580__A1_N _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19614_ _19453_/A _19453_/B _19451_/X vssd1 vssd1 vccd1 vccd1 _19616_/B sky130_fd_sc_hd__a21oi_2
X_16826_ _16844_/A vssd1 vssd1 vccd1 vccd1 _16826_/Y sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_41_clk_i_A _21822_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14876__B _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16757_ _16704_/X _16755_/Y _16754_/Y _16754_/A vssd1 vssd1 vccd1 vccd1 _16757_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16794__D _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19545_ _20146_/B _18773_/B _19546_/D _19906_/A vssd1 vssd1 vccd1 vccd1 _19548_/C
+ sky130_fd_sc_hd__a22o_1
X_13969_ _12291_/B _13967_/X _13968_/X vssd1 vssd1 vccd1 vccd1 _13969_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_49_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11581__A _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15708_ _15709_/A _15709_/B vssd1 vssd1 vccd1 vccd1 _15708_/Y sky130_fd_sc_hd__nand2_1
X_16688_ _17141_/A _17141_/B _17433_/A _17526_/B vssd1 vssd1 vccd1 vccd1 _16691_/A
+ sky130_fd_sc_hd__nand4_2
X_19476_ _19476_/A _19476_/B vssd1 vssd1 vccd1 vccd1 _19476_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_119_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15639_ _15763_/A _15638_/X _15770_/A vssd1 vssd1 vccd1 vccd1 _15641_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__13035__B1 _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18427_ _19487_/B _18873_/A _18732_/C _19221_/C vssd1 vssd1 vccd1 vccd1 _18429_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_150_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_963 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18358_ _18357_/B _18357_/C _18357_/A vssd1 vssd1 vccd1 vccd1 _18360_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_51_1181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19179__B _19493_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17309_ _17307_/X _17309_/B vssd1 vssd1 vccd1 vccd1 _17310_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16524__A1 _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18289_ _18290_/B _18290_/A vssd1 vssd1 vccd1 vccd1 _18414_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__16524__B2 _16743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17721__B1 _18894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20320_ _20321_/B _20321_/C _20321_/A vssd1 vssd1 vccd1 vccd1 _20322_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_82_1119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20251_ _20251_/A _20251_/B vssd1 vssd1 vccd1 vccd1 _20253_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_101_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout104_A _19691_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20084__A1 _19636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20084__B2 _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12561__A2 _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20182_ _20029_/X _20035_/A _20035_/B _20031_/B vssd1 vssd1 vccd1 vccd1 _20184_/B
+ sky130_fd_sc_hd__o31ai_2
XFILLER_0_0_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18029__A1 _19823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11756__A _12268_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20432__A2_N _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18029__B2 _18030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17146__C _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20387__A2 _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17443__A _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16059__A _16173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1019 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_1271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21705_ _22096_/CLK _21705_/D vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__16763__A1 _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21636_ _21722_/CLK hold257/X fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[99] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19089__B _19089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20309__A _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout17_A fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19701__A1 _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20847__B1 _10798_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19701__B2 _19868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15410__B _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16515__A1 _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16515__B2 _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21567_ mstream_o[30] hold53/X _21568_/S vssd1 vssd1 vccd1 vccd1 _22094_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_35_679 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11320_ hold241/X _11319_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21781_/D sky130_fd_sc_hd__mux2_1
X_20518_ _20391_/A _20559_/B _20399_/B _20398_/B _20398_/A vssd1 vssd1 vccd1 vccd1
+ _20533_/A sky130_fd_sc_hd__a32o_1
XFILLER_0_133_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21498_ hold261/X sstream_i[75] _21510_/S vssd1 vssd1 vccd1 vccd1 _22025_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14026__B _14663_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11251_ fanout59/X v0z[6] fanout19/X _11250_/X vssd1 vssd1 vccd1 vccd1 _11251_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20449_ _20449_/A _20449_/B _20449_/C vssd1 vssd1 vccd1 vccd1 _20450_/C sky130_fd_sc_hd__and3_1
XFILLER_0_132_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12552__A2 _12897_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11182_ hold162/X fanout22/X _11181_/X vssd1 vssd1 vccd1 vccd1 _11182_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17337__B _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14829__A1 _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15990_ _15987_/X _15988_/Y _15861_/Y _15863_/Y vssd1 vssd1 vccd1 vccd1 _15991_/C
+ sky130_fd_sc_hd__a211oi_1
X_14941_ _14778_/A _14777_/A _14777_/B _14773_/B _14773_/A vssd1 vssd1 vccd1 vccd1
+ _14942_/B sky130_fd_sc_hd__o32ai_4
XANTENNA__20378__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17779__B1 _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21575__A1 _11057_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17660_ _19892_/A _19432_/A _17777_/A _17659_/D vssd1 vssd1 vccd1 vccd1 _17660_/X
+ sky130_fd_sc_hd__a22o_1
X_14872_ _15093_/B _14871_/X _14870_/X vssd1 vssd1 vccd1 vccd1 _14874_/A sky130_fd_sc_hd__a21bo_1
X_16611_ _21824_/Q _18166_/A vssd1 vssd1 vccd1 vccd1 _16613_/B sky130_fd_sc_hd__and2_1
X_13823_ _13983_/B _16404_/B _13821_/Y _13979_/A vssd1 vssd1 vccd1 vccd1 _13827_/A
+ sky130_fd_sc_hd__o2bb2a_1
X_17591_ _17590_/A _17593_/A _17705_/A vssd1 vssd1 vccd1 vccd1 _17592_/B sky130_fd_sc_hd__a21boi_2
XFILLER_0_58_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_16542_ _17282_/A _17739_/C _17739_/D _17277_/A vssd1 vssd1 vccd1 vccd1 _16543_/B
+ sky130_fd_sc_hd__a22o_1
X_19330_ _19810_/D _20838_/C _20838_/D _19650_/D vssd1 vssd1 vccd1 vccd1 _19330_/X
+ sky130_fd_sc_hd__a22o_1
X_13754_ _13754_/A _13754_/B vssd1 vssd1 vccd1 vccd1 _13756_/B sky130_fd_sc_hd__xor2_1
X_10966_ mstream_o[59] _10965_/Y _11005_/S vssd1 vssd1 vccd1 vccd1 _21596_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_70_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_930 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_19261_ _20394_/B _19262_/C _19414_/C _19972_/A vssd1 vssd1 vccd1 vccd1 _19264_/C
+ sky130_fd_sc_hd__a22o_1
X_12705_ _12947_/A _12831_/C vssd1 vssd1 vccd1 vccd1 _12825_/C sky130_fd_sc_hd__nand2b_2
XFILLER_0_70_1056 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16473_ _17636_/B _17493_/A _16472_/C _16472_/D vssd1 vssd1 vccd1 vccd1 _16474_/B
+ sky130_fd_sc_hd__a22oi_1
X_13685_ _13685_/A _13685_/B vssd1 vssd1 vccd1 vccd1 _13687_/B sky130_fd_sc_hd__and2_1
XFILLER_0_85_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10897_ _10897_/A _10897_/B vssd1 vssd1 vccd1 vccd1 _10902_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18212_ _18212_/A _18212_/B _18212_/C vssd1 vssd1 vccd1 vccd1 _18215_/B sky130_fd_sc_hd__nand3_4
X_15424_ _15283_/Y _15285_/Y _15422_/X _15423_/Y vssd1 vssd1 vccd1 vccd1 _15426_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_26_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17622__A1_N _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19192_ _19192_/A _19192_/B vssd1 vssd1 vccd1 vccd1 _19194_/B sky130_fd_sc_hd__or2_1
X_12636_ _12716_/A _12634_/Y _12522_/B _12522_/Y vssd1 vssd1 vccd1 vccd1 _12697_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_26_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18143_ _18143_/A _18143_/B vssd1 vssd1 vccd1 vccd1 _18143_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15355_ _15492_/A _15209_/B _15204_/A vssd1 vssd1 vccd1 vccd1 _15356_/B sky130_fd_sc_hd__o21ba_1
XFILLER_0_54_966 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12567_ _12567_/A _12567_/B _12567_/C vssd1 vssd1 vccd1 vccd1 _12570_/A sky130_fd_sc_hd__nand3_1
XANTENNA__14217__A _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11340__S _11348_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14306_ _14306_/A _14621_/D _16084_/D vssd1 vssd1 vccd1 vccd1 _14306_/X sky130_fd_sc_hd__and3_1
XFILLER_0_81_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11518_ _11517_/X _19221_/C _11521_/S vssd1 vssd1 vccd1 vccd1 _21844_/D sky130_fd_sc_hd__mux2_1
X_18074_ _18074_/A _18074_/B _18074_/C vssd1 vssd1 vccd1 vccd1 _18077_/B sky130_fd_sc_hd__nand3_4
X_15286_ _15286_/A _15286_/B vssd1 vssd1 vccd1 vccd1 _15288_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_0_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12498_ _12496_/B _12388_/Y _12497_/B _12496_/X vssd1 vssd1 vccd1 vccd1 _12498_/Y
+ sky130_fd_sc_hd__o31ai_1
Xhold208 hold208/A vssd1 vssd1 vccd1 vccd1 hold208/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold219 hold219/A vssd1 vssd1 vccd1 vccd1 hold219/X sky130_fd_sc_hd__dlygate4sd3_1
X_17025_ _17025_/A _17025_/B _17025_/C vssd1 vssd1 vccd1 vccd1 _17073_/A sky130_fd_sc_hd__nand3_1
X_14237_ _14237_/A _14237_/B _14403_/B vssd1 vssd1 vccd1 vccd1 _14237_/X sky130_fd_sc_hd__and3_1
XFILLER_0_40_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11449_ _11448_/X _21056_/B _11470_/S vssd1 vssd1 vccd1 vccd1 _21821_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18350__C _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14168_ _14301_/B _14168_/B _14303_/A _14168_/D vssd1 vssd1 vccd1 vccd1 _14303_/B
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_81_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15977__A2_N _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ _14936_/D _14306_/A _21776_/Q _21777_/Q vssd1 vssd1 vccd1 vccd1 _13121_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14099_ _14098_/A _14098_/B _14098_/C vssd1 vssd1 vccd1 vccd1 _14101_/C sky130_fd_sc_hd__a21o_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18976_ _18975_/B _18975_/C _18975_/A vssd1 vssd1 vccd1 vccd1 _18976_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__15493__A1 _14916_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16690__B1 _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17927_ _17927_/A _17927_/B vssd1 vssd1 vccd1 vccd1 _17928_/B sky130_fd_sc_hd__nor2_1
XANTENNA__18431__A1 _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17858_ _18857_/B _19223_/B _17857_/C _17857_/D vssd1 vssd1 vccd1 vccd1 _17859_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__18431__B2 _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16442__B1 _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16809_ _16810_/A _16810_/B _16810_/C vssd1 vssd1 vccd1 vccd1 _16809_/X sky130_fd_sc_hd__and3_1
XFILLER_0_117_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17789_ _17670_/B _17788_/X _17787_/X vssd1 vssd1 vccd1 vccd1 _17790_/B sky130_fd_sc_hd__a21bo_1
XANTENNA__11515__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19528_ _19686_/B _21278_/A _20265_/D _20721_/D vssd1 vssd1 vccd1 vccd1 _19528_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_113_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16745__A1 _16813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19459_ _19460_/A _19460_/B vssd1 vssd1 vccd1 vccd1 _19459_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20541__A2 _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16745__B2 _16743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16326__B _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21421_ hold187/X _21420_/X _21421_/S vssd1 vssd1 vccd1 vccd1 _21949_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_56_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout221_A _21311_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout319_A _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16045__C _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21352_ _21412_/A _21352_/B vssd1 vssd1 vccd1 vccd1 _21352_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11990__B1 _12530_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20303_ _20302_/A _20302_/B _20302_/C vssd1 vssd1 vccd1 vccd1 _20303_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_13_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout2 fanout4/A vssd1 vssd1 vccd1 vccd1 fanout2/X sky130_fd_sc_hd__buf_4
X_21283_ _21283_/A _21283_/B vssd1 vssd1 vccd1 vccd1 _21285_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_97_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20234_ _20235_/A _20235_/B vssd1 vssd1 vccd1 vccd1 _20386_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_12_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout590_A _11224_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20165_ _20166_/A _20166_/B vssd1 vssd1 vccd1 vccd1 _20165_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_0_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12298__A1 _12402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20096_ _20097_/A _20097_/B vssd1 vssd1 vccd1 vccd1 _20096_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_23_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17173__A _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17225__A2 _19430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_1192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15787__A2 _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11425__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10820_ hold203/A hold215/A vssd1 vssd1 vccd1 vccd1 _10821_/B sky130_fd_sc_hd__or2_1
XTAP_2958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20998_ _20999_/A _20999_/B _20999_/C vssd1 vssd1 vccd1 vccd1 _20998_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_156_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13470_ _13468_/X _13470_/B vssd1 vssd1 vccd1 vccd1 _13471_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_82_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14211__A2 _14212_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12421_ _12510_/A vssd1 vssd1 vccd1 vccd1 _12421_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_118_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21619_ _21939_/CLK _21619_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[82] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_118_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14037__A _21741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18732__A _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15140_ _15140_/A _15253_/A _15140_/C vssd1 vssd1 vccd1 vccd1 _15253_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_106_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_9_clk_i_A _21806_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12352_ _13155_/B _12780_/A _12780_/B _13157_/A vssd1 vssd1 vccd1 vccd1 _12354_/A
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_105_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11303_ fanout58/X v0z[19] fanout18/X _11302_/X vssd1 vssd1 vccd1 vccd1 _11303_/X
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_50_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15071_ _21720_/Q hold87/X _10919_/X fanout6/A _15070_/Y vssd1 vssd1 vccd1 vccd1
+ _15071_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_65_1158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12780__A _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12283_ _12174_/X _12175_/Y _12282_/X _12173_/X vssd1 vssd1 vccd1 vccd1 _12283_/X
+ sky130_fd_sc_hd__a31o_1
X_14022_ _14508_/A _15808_/C _14354_/C _14024_/B vssd1 vssd1 vccd1 vccd1 _14027_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19989__A1 fanout96/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ _21718_/D t1x[2] v2z[2] _21724_/D _11233_/X vssd1 vssd1 vccd1 vccd1 _11234_/X
+ sky130_fd_sc_hd__a221o_2
X_18830_ _18830_/A _18830_/B _18830_/C vssd1 vssd1 vccd1 vccd1 _18833_/B sky130_fd_sc_hd__nor3_2
X_11165_ _12444_/B _11164_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21738_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15973_ _15973_/A _15973_/B vssd1 vssd1 vccd1 vccd1 _15981_/A sky130_fd_sc_hd__nand2_1
X_18761_ _18758_/Y _18759_/X _18631_/X _18669_/A vssd1 vssd1 vccd1 vccd1 _18761_/X
+ sky130_fd_sc_hd__a211o_1
X_11096_ _11057_/Y hold16/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21690_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12004__B _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14924_ _14924_/A _14924_/B vssd1 vssd1 vccd1 vccd1 _15060_/A sky130_fd_sc_hd__or2_1
XFILLER_0_101_1089 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17712_ hold229/X _17711_/X fanout3/X vssd1 vssd1 vccd1 vccd1 _21891_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_117_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18692_ _18683_/A _18683_/B _18682_/A vssd1 vssd1 vccd1 vccd1 _18834_/A sky130_fd_sc_hd__a21oi_4
Xhold80 hold80/A vssd1 vssd1 vccd1 vccd1 hold80/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 hold91/A vssd1 vssd1 vccd1 vccd1 hold91/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14857__D _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14855_ _14716_/A _16380_/B _14848_/C _14712_/X vssd1 vssd1 vccd1 vccd1 _14860_/A
+ sky130_fd_sc_hd__a31o_1
X_17643_ _19823_/A _18319_/B _18622_/B _18030_/B vssd1 vssd1 vccd1 vccd1 _17643_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11843__B _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20771__A2 _15888_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13806_ _13652_/C _13652_/Y _13804_/X _13805_/X vssd1 vssd1 vccd1 vccd1 _13806_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__13116__A _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17574_ _17575_/A _17575_/B _17575_/C _17575_/D vssd1 vssd1 vccd1 vccd1 _17574_/Y
+ sky130_fd_sc_hd__nor4_2
X_14786_ _15702_/D _15788_/B _14656_/X _14657_/X _15653_/C vssd1 vssd1 vccd1 vccd1
+ _14791_/A sky130_fd_sc_hd__a32o_1
XANTENNA__20648__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12020__A _12020_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11998_ _11924_/A _11924_/B _11924_/C vssd1 vssd1 vccd1 vccd1 _11999_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_133_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16525_ _16525_/A _16525_/B _16525_/C vssd1 vssd1 vccd1 vccd1 _16532_/A sky130_fd_sc_hd__nand3_2
X_19313_ _19313_/A _19313_/B vssd1 vssd1 vccd1 vccd1 _19316_/A sky130_fd_sc_hd__xnor2_1
X_13737_ _13734_/Y _13735_/X _13603_/X _13643_/A vssd1 vssd1 vccd1 vccd1 _13737_/X
+ sky130_fd_sc_hd__a211o_2
X_10949_ hold263/A hold273/A _10946_/A vssd1 vssd1 vccd1 vccd1 _10950_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16456_ _16456_/A _16456_/B vssd1 vssd1 vccd1 vccd1 _16703_/B sky130_fd_sc_hd__xnor2_2
X_19244_ _19243_/B _19243_/C _19243_/A vssd1 vssd1 vccd1 vccd1 _19246_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_144_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13668_ _13668_/A _13668_/B vssd1 vssd1 vccd1 vccd1 _13814_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_128_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12674__B _12785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15407_ _15407_/A _15407_/B vssd1 vssd1 vccd1 vccd1 _15415_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_112_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18064__D _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19175_ _19046_/A _19176_/B _19045_/B _19047_/Y vssd1 vssd1 vccd1 vccd1 _19313_/A
+ sky130_fd_sc_hd__o31ai_2
X_12619_ _12619_/A _13556_/A _13269_/C _12991_/D vssd1 vssd1 vccd1 vccd1 _12732_/A
+ sky130_fd_sc_hd__and4_1
X_16387_ _16387_/A _16387_/B vssd1 vssd1 vccd1 vccd1 _16393_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_115_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13599_ _13600_/A _13600_/B vssd1 vssd1 vccd1 vccd1 _13599_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_27_988 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18126_ _18126_/A _18126_/B vssd1 vssd1 vccd1 vccd1 _18129_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_42_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15338_ _15338_/A _15338_/B _15338_/C vssd1 vssd1 vccd1 vccd1 _15340_/A sky130_fd_sc_hd__nor3_2
XFILLER_0_124_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18057_ _18057_/A _18057_/B vssd1 vssd1 vccd1 vccd1 _18077_/A sky130_fd_sc_hd__xor2_2
X_15269_ _15270_/A _15270_/B vssd1 vssd1 vccd1 vccd1 _15464_/B sky130_fd_sc_hd__or2_1
XFILLER_0_77_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17008_ _17005_/B _17005_/C _17005_/A vssd1 vssd1 vccd1 vccd1 _17008_/X sky130_fd_sc_hd__o21a_1
XFILLER_0_22_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1080 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout507 _14367_/A vssd1 vssd1 vccd1 vccd1 _13155_/A sky130_fd_sc_hd__buf_4
Xfanout518 _21740_/Q vssd1 vssd1 vccd1 vccd1 _15961_/D sky130_fd_sc_hd__clkbuf_4
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout529 _21738_/Q vssd1 vssd1 vccd1 vccd1 _14659_/A sky130_fd_sc_hd__clkbuf_4
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18959_ _20242_/D _18958_/X _18957_/X vssd1 vssd1 vccd1 vccd1 _18960_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_77_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21970_ _21974_/CLK _21970_/D vssd1 vssd1 vccd1 vccd1 hold267/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__16415__B1 _15907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20921_ _21301_/A _21305_/A _21153_/B _21151_/A vssd1 vssd1 vccd1 vccd1 _20924_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout171_A _16870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout269_A _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20852_ _20852_/A _20852_/B vssd1 vssd1 vccd1 vccd1 _20853_/A sky130_fd_sc_hd__xnor2_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19904__A1 _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19904__B2 _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20783_ _20913_/A _20783_/B vssd1 vssd1 vccd1 vccd1 _20784_/B sky130_fd_sc_hd__or2_1
XFILLER_0_18_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout436_A _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19380__A2 _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_1125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13401__B1 _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout603_A _11459_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21404_ _21412_/A _21404_/B vssd1 vssd1 vccd1 vccd1 _21404_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15895__B _16380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17143__A1 _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18271__B _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18891__A1 _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21335_ _21349_/A _12392_/B _21381_/B vssd1 vssd1 vccd1 vccd1 _21335_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18891__B2 _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13704__A1 _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13704__B2 _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21266_ _21266_/A _21266_/B vssd1 vssd1 vccd1 vccd1 _21323_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20217_ _20218_/A _20218_/B vssd1 vssd1 vccd1 vccd1 _20217_/Y sky130_fd_sc_hd__nor2_1
X_21197_ _21197_/A _21197_/B vssd1 vssd1 vccd1 vccd1 _21201_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_25_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11647__C _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_1055 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15807__A2_N _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout84_A _21846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14023__C _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20148_ _20145_/Y _20281_/A _20148_/C _20924_/A vssd1 vssd1 vccd1 vccd1 _20281_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_95_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12970_ _12971_/A _12971_/B _12971_/C vssd1 vssd1 vccd1 vccd1 _13218_/A sky130_fd_sc_hd__a21oi_2
X_20079_ _20079_/A _20079_/B vssd1 vssd1 vccd1 vccd1 _20372_/A sky130_fd_sc_hd__nand2_1
XTAP_3401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17334__C _17666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11921_ _12094_/A _12094_/B _12637_/B _12639_/A vssd1 vssd1 vccd1 vccd1 _11922_/B
+ sky130_fd_sc_hd__and4_1
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14640_ _14640_/A _14640_/B _14640_/C vssd1 vssd1 vccd1 vccd1 _14642_/B sky130_fd_sc_hd__nand3_2
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ _12637_/B _11556_/X _11851_/X vssd1 vssd1 vccd1 vccd1 _11853_/B sky130_fd_sc_hd__a21bo_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21153__A _21264_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10803_ hold51/A hold151/A vssd1 vssd1 vccd1 vccd1 _10859_/A sky130_fd_sc_hd__nand2_1
X_14571_ _14571_/A _14571_/B vssd1 vssd1 vccd1 vccd1 _14575_/A sky130_fd_sc_hd__nor2_2
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11783_ _11758_/A _11758_/C _11758_/B vssd1 vssd1 vccd1 vccd1 _11784_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16310_ _16311_/B _16310_/B vssd1 vssd1 vccd1 vccd1 _16312_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_71_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14693__C _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15151__A _15151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13522_ _14294_/D _13366_/Y _13517_/Y _14293_/A vssd1 vssd1 vccd1 vccd1 _13664_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_32_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12994__A2 _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17290_ _17290_/A _17290_/B vssd1 vssd1 vccd1 vccd1 _17293_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_1168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16241_ _16347_/A _16240_/B _16348_/B _16240_/D vssd1 vssd1 vccd1 vccd1 _16241_/X
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_82_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13453_ _13299_/X _13301_/X _13450_/X _13451_/Y vssd1 vssd1 vccd1 vccd1 _13453_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_36_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18462__A _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20269__A1 _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20269__B2 _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12404_ _12403_/A _12858_/C _12991_/D _12403_/B vssd1 vssd1 vccd1 vccd1 _12405_/B
+ sky130_fd_sc_hd__a22o_1
X_16172_ _15894_/B _16028_/B _15894_/A vssd1 vssd1 vccd1 vccd1 _16287_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_91_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13384_ _13384_/A _13384_/B vssd1 vssd1 vccd1 vccd1 _13386_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_24_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15123_ _15122_/A _15266_/B _15122_/C vssd1 vssd1 vccd1 vccd1 _15124_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_23_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12335_ _12336_/A _12336_/B _12336_/C vssd1 vssd1 vccd1 vccd1 _12416_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_133_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15054_ _15055_/A _15055_/B vssd1 vssd1 vccd1 vccd1 _15054_/Y sky130_fd_sc_hd__nand2_1
X_19931_ _19932_/B _19932_/A vssd1 vssd1 vccd1 vccd1 _20072_/A sky130_fd_sc_hd__nand2b_1
X_12266_ _12267_/A _12269_/D _12267_/C _12267_/D vssd1 vssd1 vccd1 vccd1 _12271_/A
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__15932__A1_N _15933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14214__B _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14005_ _14004_/B _14004_/C _13993_/Y vssd1 vssd1 vccd1 vccd1 _14005_/Y sky130_fd_sc_hd__a21boi_2
XANTENNA__13171__A2 _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11217_ hold120/X fanout51/X fanout48/X hold237/A vssd1 vssd1 vccd1 vccd1 _11217_/X
+ sky130_fd_sc_hd__a22o_1
X_19862_ _19863_/A _19863_/B _19863_/C vssd1 vssd1 vccd1 vccd1 _19885_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12197_ _12197_/A _12197_/B vssd1 vssd1 vccd1 vccd1 _12199_/C sky130_fd_sc_hd__nor2_1
XANTENNA__11557__C _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18813_ _18813_/A _18813_/B _18813_/C vssd1 vssd1 vccd1 vccd1 _18813_/Y sky130_fd_sc_hd__nand3_2
X_11148_ hold260/X _11126_/A _11126_/B hold149/X vssd1 vssd1 vccd1 vccd1 _11148_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_128_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19793_ _20770_/B _21387_/B vssd1 vssd1 vccd1 vccd1 _19793_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__17525__B _20249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18744_ _18742_/X _18744_/B vssd1 vssd1 vccd1 vccd1 _18745_/B sky130_fd_sc_hd__nand2b_1
X_15956_ _16092_/D _21787_/Q _15957_/C _15957_/D vssd1 vssd1 vccd1 vccd1 _15958_/A
+ sky130_fd_sc_hd__a22oi_1
X_11079_ _10934_/Y hold18/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21674_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12669__B _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14907_ _14755_/A _14755_/B _14753_/Y vssd1 vssd1 vccd1 vccd1 _14909_/B sky130_fd_sc_hd__a21oi_1
X_15887_ _16016_/A _15758_/B _15756_/A vssd1 vssd1 vccd1 vccd1 _15888_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_608 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18675_ _18674_/A _18674_/B _18674_/C _18674_/D vssd1 vssd1 vccd1 vccd1 _18675_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_37_1024 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17626_ _17627_/A _17627_/B vssd1 vssd1 vccd1 vccd1 _17749_/B sky130_fd_sc_hd__nand2_1
X_14838_ _14836_/A _14836_/B _14836_/C vssd1 vssd1 vccd1 vccd1 _14840_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_114_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14769_ _14769_/A _14769_/B vssd1 vssd1 vccd1 vccd1 _14771_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_86_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17557_ _17557_/A _17557_/B _17670_/B _20270_/C vssd1 vssd1 vccd1 vccd1 _17559_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__16157__A _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16508_ _17144_/A _17526_/B _17223_/A _17129_/B vssd1 vssd1 vccd1 vccd1 _16508_/Y
+ sky130_fd_sc_hd__a22oi_1
X_17488_ _17488_/A _17488_/B _17489_/B vssd1 vssd1 vccd1 vccd1 _17704_/A sky130_fd_sc_hd__or3_4
XFILLER_0_74_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_1022 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19227_ _19379_/B _19382_/A _19227_/C _19227_/D vssd1 vssd1 vccd1 vccd1 _19230_/D
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_143_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16439_ _10988_/Y fanout5/X _16438_/X vssd1 vssd1 vccd1 vccd1 _16439_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_147_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17125__A1 _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19158_ _19159_/A _19159_/B vssd1 vssd1 vccd1 vccd1 _19320_/B sky130_fd_sc_hd__and2_1
XFILLER_0_147_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17125__B2 _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18109_ _19008_/D _19223_/B _17993_/B _17991_/X vssd1 vssd1 vccd1 vccd1 _18114_/A
+ sky130_fd_sc_hd__a31oi_1
XFILLER_0_147_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19089_ _20103_/A _19089_/B vssd1 vssd1 vccd1 vccd1 _19090_/B sky130_fd_sc_hd__and2_1
XFILLER_0_44_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21120_ _21003_/Y _21005_/X _21236_/A _21119_/X vssd1 vssd1 vccd1 vccd1 _21236_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__16884__B1 _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21051_ _21052_/A _21052_/B vssd1 vssd1 vccd1 vccd1 _21207_/B sky130_fd_sc_hd__or2_1
XFILLER_0_121_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout304 _17504_/C vssd1 vssd1 vccd1 vccd1 _17086_/C sky130_fd_sc_hd__clkbuf_4
XANTENNA__19822__B1 _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout315 _21792_/Q vssd1 vssd1 vccd1 vccd1 _17282_/A sky130_fd_sc_hd__buf_4
XANTENNA__16620__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout326 hold319/A vssd1 vssd1 vccd1 vccd1 _16314_/D sky130_fd_sc_hd__clkbuf_8
X_20002_ _19867_/A _19869_/B _19867_/B vssd1 vssd1 vccd1 vccd1 _20007_/A sky130_fd_sc_hd__a21boi_1
Xfanout337 _21784_/Q vssd1 vssd1 vccd1 vccd1 _16328_/B sky130_fd_sc_hd__buf_4
Xfanout348 hold241/A vssd1 vssd1 vccd1 vccd1 _13997_/C sky130_fd_sc_hd__clkbuf_8
XANTENNA__16977__D _17124_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout359 _14176_/C vssd1 vssd1 vccd1 vccd1 _16391_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__10920__A1 _10919_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout386_A _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13682__C _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14140__A _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__18928__A2 _18773_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19050__A1 _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21953_ _21963_/CLK _21953_/D vssd1 vssd1 vccd1 vccd1 hold317/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__19050__B2 _20026_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19650__B _20178_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout553_A _13554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18547__A _18703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20904_ _20904_/A _20904_/B _20904_/C _20904_/D vssd1 vssd1 vccd1 vccd1 _20906_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_90_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17600__A2 _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21884_ _21948_/CLK hold93/X vssd1 vssd1 vccd1 vccd1 hold92/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20835_ _20747_/B _20835_/B vssd1 vssd1 vccd1 vccd1 _20883_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__19889__B1 _20265_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11930__C _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20766_ _20634_/Y _20638_/A _20896_/B _20764_/X vssd1 vssd1 vccd1 vccd1 _20904_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_147_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20697_ _20698_/A _20698_/B _20698_/C vssd1 vssd1 vccd1 vccd1 _20699_/B sky130_fd_sc_hd__a21o_1
XANTENNA__14018__C _14018_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18432__D _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12120_ _12120_/A _12120_/B _12120_/C vssd1 vssd1 vccd1 vccd1 _12121_/B sky130_fd_sc_hd__or3_1
X_21318_ _21318_/A _21318_/B vssd1 vssd1 vccd1 vccd1 _21319_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__11658__B _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19825__B _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12051_ _12050_/B _12050_/C _12050_/A vssd1 vssd1 vccd1 vccd1 _12053_/B sky130_fd_sc_hd__a21bo_1
X_21249_ _11550_/B _16362_/Y fanout8/X vssd1 vssd1 vccd1 vccd1 _21249_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_102_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_1040 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11002_ mstream_o[76] hold55/X _11012_/S vssd1 vssd1 vccd1 vccd1 _21613_/D sky130_fd_sc_hd__mux2_1
XANTENNA__12900__A2 _12899_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11674__A _12223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15810_ _15811_/A _15811_/B vssd1 vssd1 vccd1 vccd1 _15940_/A sky130_fd_sc_hd__or2_1
X_16790_ _16790_/A _17165_/A vssd1 vssd1 vccd1 vccd1 _16792_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_99_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15741_ _15741_/A _15741_/B _15741_/C _15741_/D vssd1 vssd1 vccd1 vccd1 _15741_/X
+ sky130_fd_sc_hd__or4_2
XTAP_3220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12953_ fanout9/X _17834_/B vssd1 vssd1 vccd1 vccd1 _12953_/Y sky130_fd_sc_hd__nor2_1
XTAP_3231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11904_ _11836_/Y _11902_/X _11901_/X _11894_/X vssd1 vssd1 vccd1 vccd1 _11905_/B
+ sky130_fd_sc_hd__a211oi_2
X_15672_ _15675_/D vssd1 vssd1 vccd1 vccd1 _15672_/Y sky130_fd_sc_hd__inv_2
XTAP_3264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18460_ _18456_/X _18457_/Y _18305_/A _18305_/Y vssd1 vssd1 vccd1 vccd1 _18521_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA_220 hold277/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12884_ _12884_/A _12884_/B _12884_/C vssd1 vssd1 vccd1 vccd1 _12887_/A sky130_fd_sc_hd__nand3_1
XTAP_3286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_231 hold290/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14623_ _14621_/D _15838_/B _16374_/B _14463_/D vssd1 vssd1 vccd1 vccd1 _14624_/B
+ sky130_fd_sc_hd__o2bb2a_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17411_ _17520_/B _17619_/A _20774_/A _20774_/B vssd1 vssd1 vccd1 vccd1 _17413_/C
+ sky130_fd_sc_hd__nand4_2
XANTENNA_242 _11347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18391_ _21142_/A _21361_/B vssd1 vssd1 vccd1 vccd1 _18391_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_253 v0z[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11835_ _11801_/X _11831_/Y _11829_/X _11826_/Y vssd1 vssd1 vccd1 vccd1 _11836_/C
+ sky130_fd_sc_hd__a211o_1
XANTENNA_264 hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_275 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_286 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17342_ _17240_/A _17240_/C _17240_/B vssd1 vssd1 vccd1 vccd1 _17343_/C sky130_fd_sc_hd__a21bo_1
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14554_ _14554_/A _14554_/B vssd1 vssd1 vccd1 vccd1 _14563_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_135_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_297 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11766_ _11748_/A _11748_/B _11748_/C vssd1 vssd1 vccd1 vccd1 _11767_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_67_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13505_ _13500_/X _13502_/Y _13353_/B _13353_/Y vssd1 vssd1 vccd1 vccd1 _13505_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_126_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13113__B _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17273_ hold132/X fanout7/X _17272_/X vssd1 vssd1 vccd1 vccd1 _17273_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_71_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14485_ _14484_/B _14484_/C _14473_/Y vssd1 vssd1 vccd1 vccd1 _14485_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_0_83_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11697_ _12330_/B _11697_/B _11697_/C vssd1 vssd1 vccd1 vccd1 _12318_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_36_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16224_ _16337_/B _16224_/B vssd1 vssd1 vccd1 vccd1 _16226_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_126_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19012_ _19493_/D _19013_/C _19179_/C _19337_/D vssd1 vssd1 vccd1 vccd1 _19012_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13436_ _14195_/A _13875_/B _14384_/A _14212_/B vssd1 vssd1 vccd1 vccd1 _13437_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_70_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16424__B _21784_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19438__D _21056_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16155_ _16324_/A vssd1 vssd1 vccd1 vccd1 _16157_/D sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_31_clk_i clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _22106_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_144_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13367_ _14294_/D _13366_/Y _13365_/X vssd1 vssd1 vccd1 vccd1 _13368_/B sky130_fd_sc_hd__a21boi_4
XANTENNA__17658__A2 _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15106_ _15254_/A _15104_/Y _15004_/B _15006_/B vssd1 vssd1 vccd1 vccd1 _15108_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_11_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12318_ _12318_/A _12318_/B vssd1 vssd1 vccd1 vccd1 _12338_/A sky130_fd_sc_hd__nand2_1
X_16086_ _16087_/A _16404_/B _16087_/C _16087_/D vssd1 vssd1 vccd1 vccd1 _16088_/A
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__11568__B _12155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13298_ _13298_/A _13298_/B vssd1 vssd1 vccd1 vccd1 _13300_/B sky130_fd_sc_hd__and2_1
XFILLER_0_107_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15037_ _15037_/A _15037_/B _15037_/C vssd1 vssd1 vccd1 vccd1 _15040_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_20_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19914_ _19914_/A _19914_/B _19914_/C vssd1 vssd1 vccd1 vccd1 _19917_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_121_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12249_ _12268_/A _21727_/Q _12249_/C _12249_/D vssd1 vssd1 vccd1 vccd1 _12264_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1095 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12352__B1 _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21058__A _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19280__A1 _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19845_ _19961_/A vssd1 vssd1 vccd1 vccd1 _20380_/A sky130_fd_sc_hd__inv_2
XFILLER_0_78_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19751__A _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19776_ _19776_/A _19776_/B vssd1 vssd1 vccd1 vccd1 _19777_/B sky130_fd_sc_hd__xnor2_1
X_16988_ _17029_/A _17145_/B _17146_/C _17029_/B vssd1 vssd1 vccd1 vccd1 _16988_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_39_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18727_ _18610_/Y _18613_/Y _18847_/B _18726_/X vssd1 vssd1 vccd1 vccd1 _18846_/A
+ sky130_fd_sc_hd__a211oi_2
X_15939_ _15940_/A _15940_/B _15940_/C vssd1 vssd1 vccd1 vccd1 _16078_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_64_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18658_ _18658_/A _18658_/B _18658_/C vssd1 vssd1 vccd1 vccd1 _18661_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_59_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17609_ _17732_/A vssd1 vssd1 vccd1 vccd1 _17611_/C sky130_fd_sc_hd__inv_2
XFILLER_0_93_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18589_ _18590_/A _18590_/B vssd1 vssd1 vccd1 vccd1 _18720_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1010 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20620_ _20617_/X _20618_/Y _20485_/Y _20487_/Y vssd1 vssd1 vccd1 vccd1 _20621_/C
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_80_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11091__A0 _11045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12565__D _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15357__B1 _10934_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20551_ _20551_/A _20679_/B vssd1 vssd1 vccd1 vccd1 _20554_/A sky130_fd_sc_hd__or2_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout134_A _19087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20482_ _20483_/A _20483_/B vssd1 vssd1 vccd1 vccd1 _20484_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_36_clk_i_A clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout301_A _21795_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14465__A1_N _14463_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21103_ _21103_/A _21208_/B vssd1 vssd1 vccd1 vccd1 _21105_/B sky130_fd_sc_hd__or2_1
XFILLER_0_26_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22083_ _22096_/CLK _22083_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[19] sky130_fd_sc_hd__dfrtp_4
Xfanout101 _21842_/Q vssd1 vssd1 vccd1 vccd1 _20419_/A sky130_fd_sc_hd__clkbuf_8
Xfanout112 _21840_/Q vssd1 vssd1 vccd1 vccd1 _21267_/A sky130_fd_sc_hd__buf_4
X_21034_ _21034_/A _21034_/B vssd1 vssd1 vccd1 vccd1 _21035_/B sky130_fd_sc_hd__xnor2_1
Xfanout123 _20689_/A vssd1 vssd1 vccd1 vccd1 _21056_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_96_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout134 _19087_/B vssd1 vssd1 vccd1 vccd1 _20101_/B sky130_fd_sc_hd__buf_4
Xfanout145 _17417_/D vssd1 vssd1 vccd1 vccd1 _16899_/B sky130_fd_sc_hd__buf_4
Xfanout156 _20088_/A vssd1 vssd1 vccd1 vccd1 _19432_/A sky130_fd_sc_hd__clkbuf_8
Xfanout167 _19732_/A vssd1 vssd1 vccd1 vccd1 _19951_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__16500__D _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 _17443_/D vssd1 vssd1 vccd1 vccd1 _19587_/B sky130_fd_sc_hd__buf_4
Xfanout189 _21823_/Q vssd1 vssd1 vccd1 vccd1 _17146_/B sky130_fd_sc_hd__buf_4
XANTENNA__20169__B1 _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17181__A _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21936_ _21938_/CLK _21936_/D vssd1 vssd1 vccd1 vccd1 hold169/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout47_A fanout49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21867_ _21942_/CLK _21867_/D vssd1 vssd1 vccd1 vccd1 hold133/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__18427__D _19221_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_93_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12756__C _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _11615_/X _11617_/Y _11588_/A _11591_/A vssd1 vssd1 vccd1 vccd1 _11621_/B
+ sky130_fd_sc_hd__a211o_1
X_20818_ _20819_/A _20819_/B vssd1 vssd1 vccd1 vccd1 _20951_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15132__C _15933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21798_ _21803_/CLK _21798_/D vssd1 vssd1 vccd1 vccd1 _21798_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_132_1199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11082__A0 _10950_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_975 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11551_ _20770_/B _21142_/A vssd1 vssd1 vccd1 vccd1 _11551_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_25_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20749_ _20574_/X _20578_/B _20835_/B _20748_/Y vssd1 vssd1 vccd1 vccd1 _20750_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_108_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14270_ _14107_/X _14109_/X _14268_/X _14269_/Y vssd1 vssd1 vccd1 vccd1 _14270_/Y
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_18_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11482_ _11481_/X _18622_/B _11521_/S vssd1 vssd1 vccd1 vccd1 _21832_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_150_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13221_ _13217_/X _13219_/Y _13080_/Y _13083_/X vssd1 vssd1 vccd1 vccd1 _13222_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_21_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18740__A _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13152_ _14024_/B _14027_/A _13152_/C _13152_/D vssd1 vssd1 vccd1 vccd1 _13153_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_33_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12103_ _12223_/A _12246_/C _12096_/B _12094_/X vssd1 vssd1 vccd1 vccd1 _12106_/A
+ sky130_fd_sc_hd__a31oi_2
XANTENNA__14323__A1 _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13083_ _13083_/A _13083_/B _13083_/C vssd1 vssd1 vccd1 vccd1 _13083_/X sky130_fd_sc_hd__or3_1
XFILLER_0_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17960_ _17819_/B _17821_/A _17958_/X _17959_/Y vssd1 vssd1 vccd1 vccd1 _17962_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_1257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16911_ _17165_/A _17165_/B _17165_/C _17168_/A vssd1 vssd1 vccd1 vccd1 _16912_/B
+ sky130_fd_sc_hd__a211o_1
X_12034_ _11980_/B _12294_/C _12294_/D _12388_/B vssd1 vssd1 vccd1 vccd1 _12035_/B
+ sky130_fd_sc_hd__a31o_1
XANTENNA__18065__A2 _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17891_ _17891_/A _17891_/B vssd1 vssd1 vccd1 vccd1 _17910_/A sky130_fd_sc_hd__nand2_1
XANTENNA__13095__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19630_ _19628_/Y _19630_/B vssd1 vssd1 vccd1 vccd1 _19631_/B sky130_fd_sc_hd__and2b_1
XANTENNA__19571__A _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16842_ _16849_/B _16840_/X _16834_/Y _16837_/Y vssd1 vssd1 vccd1 vccd1 _16844_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_18_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19014__A1 _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19561_ _19560_/B _19560_/C _19560_/A vssd1 vssd1 vccd1 vccd1 _19562_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13985_ _13985_/A _16374_/B _13985_/C _13985_/D vssd1 vssd1 vccd1 vccd1 _13986_/B
+ sky130_fd_sc_hd__nor4_2
X_16773_ _16773_/A _16773_/B _16773_/C vssd1 vssd1 vccd1 vccd1 _16773_/Y sky130_fd_sc_hd__nand3_1
X_18512_ _18511_/B _18511_/C _18511_/A vssd1 vssd1 vccd1 vccd1 _18512_/Y sky130_fd_sc_hd__a21oi_2
X_15724_ _15724_/A _15724_/B vssd1 vssd1 vccd1 vccd1 _15727_/C sky130_fd_sc_hd__xnor2_1
XTAP_3050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12936_ _12807_/C _12808_/X _12934_/X _12935_/Y vssd1 vssd1 vccd1 vccd1 _12938_/B
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_137_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19492_ _19492_/A _19492_/B vssd1 vssd1 vccd1 vccd1 _19497_/A sky130_fd_sc_hd__xnor2_2
XTAP_3072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__21372__A2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18443_ _19529_/B _19068_/C _19238_/C _19373_/B vssd1 vssd1 vccd1 vccd1 _18443_/Y
+ sky130_fd_sc_hd__a22oi_1
X_15655_ _16404_/A _15913_/B _15655_/C _15849_/A vssd1 vssd1 vccd1 vccd1 _15849_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12867_ _12868_/A _12868_/B _12868_/C vssd1 vssd1 vccd1 vccd1 _12869_/B sky130_fd_sc_hd__a21o_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1098 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14606_ _21725_/D hold111/X _10892_/Y fanout6/X _14605_/Y vssd1 vssd1 vccd1 vccd1
+ _14606_/X sky130_fd_sc_hd__a221o_1
X_11818_ _11788_/A _11788_/B _11788_/C vssd1 vssd1 vccd1 vccd1 _11819_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_145_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15586_ _15586_/A _15586_/B vssd1 vssd1 vccd1 vccd1 _15605_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_111_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18374_ _18373_/A _18373_/B _18373_/C _18373_/D vssd1 vssd1 vccd1 vccd1 _18374_/Y
+ sky130_fd_sc_hd__o22ai_4
X_12798_ _12798_/A _12798_/B _12798_/C vssd1 vssd1 vccd1 vccd1 _12798_/Y sky130_fd_sc_hd__nand3_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11073__A0 _10886_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14537_ _14537_/A _16409_/A vssd1 vssd1 vccd1 vccd1 _14538_/B sky130_fd_sc_hd__nand2_1
X_17325_ _17434_/B _19430_/A _17324_/D _17433_/A vssd1 vssd1 vccd1 vccd1 _17326_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11749_ _11748_/B _11748_/C _11748_/A vssd1 vssd1 vccd1 vccd1 _11750_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_71_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13778__B _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14468_ _14316_/A _14315_/A _14315_/B _14311_/B _14311_/A vssd1 vssd1 vccd1 vccd1
+ _14469_/B sky130_fd_sc_hd__o32ai_4
XFILLER_0_4_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17256_ _17256_/A _17256_/B _17256_/C _17256_/D vssd1 vssd1 vccd1 vccd1 _17256_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_126_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16154__B _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1060 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16207_ _16207_/A _16207_/B _16207_/C vssd1 vssd1 vccd1 vccd1 _16209_/A sky130_fd_sc_hd__nor3_1
X_13419_ _13867_/A _13573_/D _13417_/Y _13569_/A vssd1 vssd1 vccd1 vccd1 _13419_/X
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17187_ _17187_/A _17187_/B vssd1 vssd1 vccd1 vccd1 _17188_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__19746__A _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14399_ _14532_/B _14398_/C _14398_/A vssd1 vssd1 vccd1 vccd1 _14399_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18650__A _19445_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16138_ _16251_/A _16136_/X _15968_/B _15970_/Y vssd1 vssd1 vccd1 vccd1 _16138_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11729__D _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16069_ _16069_/A _16069_/B _16069_/C vssd1 vssd1 vccd1 vccd1 _16070_/C sky130_fd_sc_hd__nand3_1
XANTENNA__14314__B2 _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11518__S _11521_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19828_ _19828_/A _19828_/B _19828_/C vssd1 vssd1 vccd1 vccd1 _19830_/B sky130_fd_sc_hd__nand3_2
XANTENNA__13018__B _13018_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19759_ _19759_/A vssd1 vssd1 vccd1 vccd1 _19759_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_155_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15514__A _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11300__A1 _11299_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21363__A2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21721_ _21974_/CLK _21721_/D _21422_/A vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout251_A _17334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11851__A2 _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout349_A _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_1072 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13034__A _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21652_ _21888_/CLK _21652_/D vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11064__A0 _11063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20603_ _20603_/A _20603_/B vssd1 vssd1 vccd1 vccd1 _20611_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11603__A2 _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21583_ _22106_/CLK _21583_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[46] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_74_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout516_A _13875_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20534_ _20918_/A _20535_/B vssd1 vssd1 vccd1 vccd1 _20536_/A sky130_fd_sc_hd__and2_1
XFILLER_0_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16542__A2 _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_1224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20047__A2_N _20193_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20465_ _20465_/A _20465_/B vssd1 vssd1 vccd1 vccd1 _20466_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19375__B _20671_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_980 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20396_ _20650_/B _20396_/B vssd1 vssd1 vccd1 vccd1 _20397_/B sky130_fd_sc_hd__and2b_1
XANTENNA__11639__D _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14305__A1 _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_1218 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14305__B2 _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14856__A2 _21755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16511__C _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22066_ _22069_/CLK _22066_/D fanout639/X vssd1 vssd1 vccd1 vccd1 mstream_o[2] sky130_fd_sc_hd__dfrtp_4
XANTENNA__16058__A1 _16284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14312__B _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20929__A2 _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16058__B2 _16173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11428__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21017_ _20880_/X _20882_/Y _21129_/A _21016_/Y vssd1 vssd1 vccd1 vccd1 _21129_/B
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__13816__B1 _10860_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__A _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ _13770_/A _13770_/B vssd1 vssd1 vccd1 vccd1 _13790_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_134_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10982_ _10982_/A _10982_/B vssd1 vssd1 vccd1 vccd1 _10984_/A sky130_fd_sc_hd__nand2_2
XANTENNA__17558__A1 _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12095__A2 _12512_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21354__A2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12721_ _12721_/A _12834_/A vssd1 vssd1 vccd1 vccd1 _12731_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_97_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21919_ _22106_/CLK _21919_/D vssd1 vssd1 vccd1 vccd1 hold132/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_57_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15033__A2 _16409_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15440_ _15442_/A vssd1 vssd1 vccd1 vccd1 _15586_/A sky130_fd_sc_hd__inv_2
XFILLER_0_66_931 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12652_ _12653_/A _12653_/B _12653_/C vssd1 vssd1 vccd1 vccd1 _12652_/X sky130_fd_sc_hd__a21o_4
XFILLER_0_139_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14241__B1 _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11603_ _12319_/C _12402_/A _12302_/A _12420_/D vssd1 vssd1 vccd1 vccd1 _11606_/C
+ sky130_fd_sc_hd__a22o_1
X_15371_ _15371_/A _15548_/B vssd1 vssd1 vccd1 vccd1 _15380_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_108_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12583_ _12583_/A _12583_/B _12583_/C _12583_/D vssd1 vssd1 vccd1 vccd1 _12583_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_80_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14322_ _14189_/A _14188_/B _14186_/X vssd1 vssd1 vccd1 vccd1 _14322_/Y sky130_fd_sc_hd__a21oi_1
X_17110_ _17110_/A _17110_/B _17110_/C vssd1 vssd1 vccd1 vccd1 _17110_/X sky130_fd_sc_hd__and3_1
XFILLER_0_37_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18090_ _18087_/X _18088_/Y _17953_/B _17952_/Y vssd1 vssd1 vccd1 vccd1 _18091_/C
+ sky130_fd_sc_hd__a211o_1
X_11534_ _11089_/B t1y[28] t0x[28] _11223_/A vssd1 vssd1 vccd1 vccd1 _11534_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_135_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_576 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_1107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17041_ _17041_/A _17146_/D vssd1 vssd1 vccd1 vccd1 _17044_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14253_ _14418_/A _14254_/C _14254_/A vssd1 vssd1 vccd1 vccd1 _14255_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11465_ _11123_/A t1y[5] t0x[5] _21724_/D vssd1 vssd1 vccd1 vccd1 _11465_/X sky130_fd_sc_hd__a22o_1
XANTENNA__19566__A _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13204_ _13204_/A _13204_/B _13204_/C vssd1 vssd1 vccd1 vccd1 _13204_/X sky130_fd_sc_hd__or3_2
XFILLER_0_21_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14184_ _14659_/A _15022_/B _14185_/C _14185_/D vssd1 vssd1 vccd1 vccd1 _14184_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_110_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11396_ _21718_/D hold266/X fanout49/X hold198/X vssd1 vssd1 vccd1 vccd1 _11396_/X
+ sky130_fd_sc_hd__a22o_1
X_13135_ _13267_/B _13134_/C _13134_/A vssd1 vssd1 vccd1 vccd1 _13136_/C sky130_fd_sc_hd__a21o_1
XANTENNA__17086__A _17146_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1021 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18992_ _18991_/B _18991_/C _18991_/A vssd1 vssd1 vccd1 vccd1 _18992_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__14847__A2 _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13066_ _13067_/A _13067_/B _13067_/C vssd1 vssd1 vccd1 vccd1 _13066_/Y sky130_fd_sc_hd__nor3_2
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17943_ _17943_/A _17943_/B _17943_/C vssd1 vssd1 vccd1 vccd1 _17943_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__13764__D _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21042__A1 _21841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13119__A _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12017_ _12017_/A _12017_/B vssd1 vssd1 vccd1 vccd1 _12023_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__21042__B2 _21267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17874_ _17874_/A _20148_/C _18006_/A _17874_/D vssd1 vssd1 vccd1 vccd1 _18006_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__11530__A1 _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19732__C _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19613_ _19613_/A _19613_/B vssd1 vssd1 vccd1 vccd1 _19616_/A sky130_fd_sc_hd__xor2_4
X_16825_ _16809_/X _16823_/X _16824_/X _16754_/Y vssd1 vssd1 vccd1 vccd1 _16844_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14876__C _16414_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19544_ _20103_/A _19546_/D _19408_/X _19409_/X _19906_/D vssd1 vssd1 vccd1 vccd1
+ _19549_/A sky130_fd_sc_hd__a32o_1
X_16756_ _16754_/A _16754_/Y _16755_/Y _16704_/X vssd1 vssd1 vccd1 vccd1 _16756_/Y
+ sky130_fd_sc_hd__a211oi_4
X_13968_ _16363_/A hold47/X _10867_/X fanout5/X vssd1 vssd1 vccd1 vccd1 _13968_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21345__A2 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15707_ _15582_/A _15712_/A _15581_/B _15578_/B _15578_/A vssd1 vssd1 vccd1 vccd1
+ _15709_/B sky130_fd_sc_hd__o32ai_4
XANTENNA__11581__B _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12919_ _12918_/B _12918_/C _12918_/A vssd1 vssd1 vccd1 vccd1 _12921_/B sky130_fd_sc_hd__a21o_1
X_19475_ _19475_/A _19475_/B vssd1 vssd1 vccd1 vccd1 _19476_/B sky130_fd_sc_hd__and2_1
X_13899_ _15763_/A _14212_/C vssd1 vssd1 vccd1 vccd1 _13901_/C sky130_fd_sc_hd__and2_1
XFILLER_0_5_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16687_ _16686_/B _16686_/C _16686_/A vssd1 vssd1 vccd1 vccd1 _16687_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18426_ _19487_/B _18732_/C _19221_/C _18873_/A vssd1 vssd1 vccd1 vccd1 _18429_/C
+ sky130_fd_sc_hd__a22o_1
X_15638_ _15517_/A _15516_/B _15763_/B vssd1 vssd1 vccd1 vccd1 _15638_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_146_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13035__A1 _13173_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13035__B2 _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11046__A0 _11045_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18357_ _18357_/A _18357_/B _18357_/C vssd1 vssd1 vccd1 vccd1 _18360_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_145_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15569_ _15426_/B _15426_/Y _15567_/X _15568_/Y vssd1 vssd1 vccd1 vccd1 _15612_/A
+ sky130_fd_sc_hd__o211a_2
XFILLER_0_127_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19179__C _19179_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17308_ _17525_/A _17417_/C _17417_/D _17520_/A vssd1 vssd1 vccd1 vccd1 _17309_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18288_ _18288_/A _18288_/B vssd1 vssd1 vccd1 vccd1 _18290_/B sky130_fd_sc_hd__and2_1
XANTENNA__16524__A2 _17504_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17721__A1 _17854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_1256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17721__B2 _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17239_ _17915_/A _17557_/B _17915_/D _17557_/A vssd1 vssd1 vccd1 vccd1 _17240_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11349__B2 _11089_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_371 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20250_ _20250_/A _20250_/B vssd1 vssd1 vccd1 vccd1 _20253_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20084__A2 _15210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17485__B1 _17484_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20181_ _20181_/A _20181_/B vssd1 vssd1 vccd1 vccd1 _20184_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__18029__A2 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11756__B _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_994 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17146__D _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11248__S _11260_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout299_A _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11521__A1 _19223_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17443__B _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout466_A _14698_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15263__A2 _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18258__C _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21336__A2 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16059__B _16284_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout633_A _21776_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21704_ _22096_/CLK _21704_/D vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21635_ _21682_/CLK hold240/X fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[98] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_997 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20309__B _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19701__A2 _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20847__B2 _20721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21566_ mstream_o[29] hold61/X _21579_/S vssd1 vssd1 vccd1 vccd1 _22093_/D sky130_fd_sc_hd__mux2_1
XANTENNA_hold309_A hold309/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16515__A2 _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20028__C _20178_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20517_ hold273/X _20516_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _21910_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21497_ hold316/X sstream_i[74] _21507_/S vssd1 vssd1 vccd1 vccd1 _22024_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_132_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11250_ _11502_/A1 t1x[6] v2z[6] _21724_/D _11249_/X vssd1 vssd1 vccd1 vccd1 _11250_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_127_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20448_ _20450_/B vssd1 vssd1 vccd1 vccd1 _20448_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_1031 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11181_ hold295/X fanout51/X fanout47/X hold281/A vssd1 vssd1 vccd1 vccd1 _11181_/X
+ sky130_fd_sc_hd__a22o_1
X_20379_ hold101/X _20378_/X fanout4/X vssd1 vssd1 vccd1 vccd1 _21909_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14829__A2 _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22049_ _22049_/CLK _22049_/D vssd1 vssd1 vccd1 vccd1 hold256/A sky130_fd_sc_hd__dfxtp_4
X_14940_ _14940_/A _14940_/B vssd1 vssd1 vccd1 vccd1 _14942_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__11512__A1 _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17779__A1 _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17779__B2 _17657_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21156__A _21267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14871_ _14993_/A _15632_/B _16418_/A vssd1 vssd1 vccd1 vccd1 _14871_/X sky130_fd_sc_hd__and3_1
XFILLER_0_89_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_5_clk_i_A _21806_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16610_ _21822_/Q _21823_/Q _17657_/A _17334_/B vssd1 vssd1 vccd1 vccd1 _16613_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_138_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13822_ _14312_/D _13822_/B _16399_/B _16409_/B vssd1 vssd1 vccd1 vccd1 _13979_/A
+ sky130_fd_sc_hd__and4_1
X_17590_ _17590_/A _17593_/A vssd1 vssd1 vccd1 vccd1 _17590_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11276__A0 _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_1160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13753_ _13754_/A _13754_/B vssd1 vssd1 vccd1 vccd1 _13753_/Y sky130_fd_sc_hd__nand2b_1
X_16541_ _17282_/A _17277_/A _17739_/C _17739_/D vssd1 vssd1 vccd1 vccd1 _16541_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_70_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10965_ _10965_/A _10965_/B vssd1 vssd1 vccd1 vccd1 _10965_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_0_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12704_ _12701_/Y _12702_/X _12589_/X _12591_/Y vssd1 vssd1 vccd1 vccd1 _12831_/C
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_85_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_1166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19260_ _19260_/A _19260_/B vssd1 vssd1 vccd1 vccd1 _19268_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13684_ _13681_/X _13835_/B _13556_/D _13557_/B vssd1 vssd1 vccd1 vccd1 _13685_/B
+ sky130_fd_sc_hd__o211ai_1
X_16472_ _17636_/B _17277_/A _16472_/C _16472_/D vssd1 vssd1 vccd1 vccd1 _16474_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_35_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10896_ _10897_/B vssd1 vssd1 vccd1 vccd1 _10911_/A sky130_fd_sc_hd__inv_2
XFILLER_0_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_964 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18211_ _18071_/A _18071_/C _18071_/B vssd1 vssd1 vccd1 vccd1 _18212_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_54_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15423_ _15420_/Y _15421_/X _15243_/X _15246_/Y vssd1 vssd1 vccd1 vccd1 _15423_/Y
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_109_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12635_ _12522_/B _12522_/Y _12716_/A _12634_/Y vssd1 vssd1 vccd1 vccd1 _12716_/B
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19191_ _19190_/A _19190_/B _19190_/C vssd1 vssd1 vccd1 vccd1 _19192_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13402__A _13554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15354_ _15354_/A _15354_/B vssd1 vssd1 vccd1 vccd1 _15492_/B sky130_fd_sc_hd__xor2_4
X_18142_ _18142_/A _18142_/B vssd1 vssd1 vccd1 vccd1 _18143_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_25_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12566_ _12785_/B _14386_/B _14384_/C _14248_/A vssd1 vssd1 vccd1 vccd1 _12567_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14217__B _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14517__A1 _14365_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14305_ _14306_/A _16084_/C _16084_/D _14621_/D vssd1 vssd1 vccd1 vccd1 _14305_/X
+ sky130_fd_sc_hd__a22o_1
X_11517_ _11224_/A t2x[22] v1z[22] fanout21/X _11516_/X vssd1 vssd1 vccd1 vccd1 _11517_/X
+ sky130_fd_sc_hd__a221o_1
X_15285_ _15286_/A _15286_/B vssd1 vssd1 vccd1 vccd1 _15285_/Y sky130_fd_sc_hd__nand2_1
X_18073_ _17937_/A _17937_/C _17937_/B vssd1 vssd1 vccd1 vccd1 _18074_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_145_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12497_ _12497_/A _12497_/B vssd1 vssd1 vccd1 vccd1 _12497_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14236_ _14859_/A _15093_/B _14236_/C _14403_/A vssd1 vssd1 vccd1 vccd1 _14403_/B
+ sky130_fd_sc_hd__nand4_2
X_17024_ _17018_/A _17018_/B _17018_/C vssd1 vssd1 vccd1 vccd1 _17025_/C sky130_fd_sc_hd__a21o_1
Xhold209 hold209/A vssd1 vssd1 vccd1 vccd1 hold209/X sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ hold251/A _11124_/Y _11447_/X vssd1 vssd1 vccd1 vccd1 _11448_/X sky130_fd_sc_hd__a21o_2
XFILLER_0_40_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14167_ _14338_/B _14165_/Y _14004_/X _14007_/A vssd1 vssd1 vccd1 vccd1 _14168_/D
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_22_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ hold298/X fanout29/X _11378_/X vssd1 vssd1 vccd1 vccd1 _11379_/X sky130_fd_sc_hd__a21o_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ _14138_/A _14018_/C vssd1 vssd1 vccd1 vccd1 _13121_/A sky130_fd_sc_hd__and2_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14098_ _14098_/A _14098_/B _14098_/C vssd1 vssd1 vccd1 vccd1 _14101_/B sky130_fd_sc_hd__nand3_4
X_18975_ _18975_/A _18975_/B _18975_/C vssd1 vssd1 vccd1 vccd1 _18975_/Y sky130_fd_sc_hd__nand3_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ _14089_/A _14087_/A _13913_/C _14077_/B vssd1 vssd1 vccd1 vccd1 _13051_/B
+ sky130_fd_sc_hd__nand4_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17926_ _19438_/B _19703_/C _18640_/B _19438_/A vssd1 vssd1 vccd1 vccd1 _17927_/B
+ sky130_fd_sc_hd__a22oi_2
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11503__A1 _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16427__D1 _16286_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17857_ _18857_/B _19223_/B _17857_/C _17857_/D vssd1 vssd1 vccd1 vccd1 _17980_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__18431__A2 _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_156_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16442__B2 _16734_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16808_ _16738_/A _16738_/B _16738_/C vssd1 vssd1 vccd1 vccd1 _16810_/C sky130_fd_sc_hd__a21o_1
X_17788_ _19438_/A _19438_/B _17924_/B vssd1 vssd1 vccd1 vccd1 _17788_/X sky130_fd_sc_hd__and3_1
XFILLER_0_49_706 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11267__B1 _11266_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19187__A2_N _19185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19527_ _19398_/A _19398_/B _19398_/C _19400_/X vssd1 vssd1 vccd1 vccd1 _19560_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_152_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16739_ _16738_/B _16738_/C _16738_/A vssd1 vssd1 vccd1 vccd1 _16741_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_89_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19458_ _19304_/A _19304_/B _19302_/X vssd1 vssd1 vccd1 vccd1 _19460_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_48_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16745__A2 _16743_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18409_ _18409_/A _18409_/B vssd1 vssd1 vccd1 vccd1 _18411_/B sky130_fd_sc_hd__and2_1
XANTENNA__15953__B1 _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19389_ _20146_/B _19692_/B _19705_/B _19906_/A vssd1 vssd1 vccd1 vccd1 _19392_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14408__A _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16326__C _16396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21420_ _16437_/Y _21324_/Y _21420_/S vssd1 vssd1 vccd1 vccd1 _21420_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_29_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16045__D _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21351_ hold96/X _21403_/S _21349_/Y _21350_/Y vssd1 vssd1 vccd1 vccd1 _21924_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_115_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20302_ _20302_/A _20302_/B _20302_/C vssd1 vssd1 vccd1 vccd1 _20302_/Y sky130_fd_sc_hd__nor3_4
XFILLER_0_114_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21282_ _21201_/A _21200_/A _21287_/A _21197_/B vssd1 vssd1 vccd1 vccd1 _21321_/A
+ sky130_fd_sc_hd__a31o_1
Xfanout3 fanout4/A vssd1 vssd1 vccd1 vccd1 fanout3/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_40_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20233_ _20089_/A _20089_/B _20087_/A vssd1 vssd1 vccd1 vccd1 _20235_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_130_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20164_ _20164_/A _20164_/B vssd1 vssd1 vccd1 vccd1 _20166_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_0_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout583_A _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12298__A2 _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20095_ _20380_/A _20095_/B vssd1 vssd1 vccd1 vccd1 _20097_/B sky130_fd_sc_hd__nand2_1
XANTENNA__14692__B1 _16418_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17173__B _17173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20997_ _20997_/A _20997_/B vssd1 vssd1 vccd1 vccd1 _20999_/C sky130_fd_sc_hd__nand2_1
XANTENNA__18285__A _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12420_ _12639_/A _12530_/A _13152_/C _12420_/D vssd1 vssd1 vccd1 vccd1 _12510_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_75_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21618_ _21906_/CLK _21618_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[81] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_36_956 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14037__B _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18732__B _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ _13017_/A _12781_/D vssd1 vssd1 vccd1 vccd1 _12355_/A sky130_fd_sc_hd__nand2_1
X_21549_ mstream_o[12] hold152/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22076_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_106_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11302_ _11224_/A t1x[19] v2z[19] _11507_/B2 _11301_/X vssd1 vssd1 vccd1 vccd1 _11302_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_22_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15070_ fanout9/X _15070_/B vssd1 vssd1 vccd1 vccd1 _15070_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_120_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12282_ _12209_/X _12281_/X _12208_/X vssd1 vssd1 vccd1 vccd1 _12282_/X sky130_fd_sc_hd__a21o_1
XANTENNA__12780__B _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14021_ _14021_/A _14021_/B vssd1 vssd1 vccd1 vccd1 _14031_/A sky130_fd_sc_hd__and2_1
X_11233_ _11122_/A t2y[2] t0y[2] _11123_/A vssd1 vssd1 vccd1 vccd1 _11233_/X sky130_fd_sc_hd__a22o_1
XANTENNA__17449__B1 _17670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14053__A _14212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16121__B1 _16119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11164_ hold123/X fanout23/X _11163_/X vssd1 vssd1 vccd1 vccd1 _11164_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_140_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18760_ _18631_/X _18669_/A _18758_/Y _18759_/X vssd1 vssd1 vccd1 vccd1 _18760_/Y
+ sky130_fd_sc_hd__o211ai_4
X_15972_ _15972_/A _15972_/B vssd1 vssd1 vccd1 vccd1 _15983_/A sky130_fd_sc_hd__or2_1
X_11095_ _11055_/Y hold15/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21689_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_101_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12004__C _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17711_ hold163/X fanout7/X _21346_/B _11547_/X _17599_/Y vssd1 vssd1 vccd1 vccd1
+ _17711_/X sky130_fd_sc_hd__a221o_1
X_14923_ _14780_/A _14780_/B _14783_/A vssd1 vssd1 vccd1 vccd1 _15065_/A sky130_fd_sc_hd__a21o_1
X_18691_ hold22/X _18690_/X fanout1/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__mux2_1
XFILLER_0_26_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold70 hold70/A vssd1 vssd1 vccd1 vccd1 hold70/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 hold81/A vssd1 vssd1 vccd1 vccd1 hold81/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 hold92/A vssd1 vssd1 vccd1 vccd1 hold92/X sky130_fd_sc_hd__dlygate4sd3_1
X_17642_ _19823_/A _18030_/B _18622_/B vssd1 vssd1 vccd1 vccd1 _17642_/X sky130_fd_sc_hd__and3_1
X_14854_ _14854_/A _14854_/B vssd1 vssd1 vccd1 vccd1 _14862_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13805_ _13819_/B _13804_/B _13802_/Y _13803_/X vssd1 vssd1 vccd1 vccd1 _13805_/X
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13116__B _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17573_ _17569_/X _17571_/Y _17461_/B _17461_/Y vssd1 vssd1 vccd1 vccd1 _17575_/D
+ sky130_fd_sc_hd__o211a_1
X_14785_ _14785_/A _14785_/B vssd1 vssd1 vccd1 vccd1 _14793_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12020__B _12326_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11997_ _11996_/B _11996_/C _11996_/A vssd1 vssd1 vccd1 vccd1 _11999_/B sky130_fd_sc_hd__a21bo_1
X_19312_ _19313_/A _19313_/B vssd1 vssd1 vccd1 vccd1 _19467_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_97_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16524_ _17206_/B _17504_/C _16459_/X _16460_/X _16743_/C vssd1 vssd1 vccd1 vccd1
+ _16525_/C sky130_fd_sc_hd__a32o_1
X_10948_ hold78/A hold276/A vssd1 vssd1 vccd1 vccd1 _10950_/A sky130_fd_sc_hd__xnor2_4
X_13736_ _13603_/X _13643_/A _13734_/Y _13735_/X vssd1 vssd1 vccd1 vccd1 _13736_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_133_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19243_ _19243_/A _19243_/B _19243_/C vssd1 vssd1 vccd1 vccd1 _19246_/A sky130_fd_sc_hd__nand3_1
X_16455_ _16989_/C _17063_/C _16454_/B _16451_/X vssd1 vssd1 vccd1 vccd1 _16703_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18345__D _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10879_ _10880_/A _10880_/B _10878_/Y vssd1 vssd1 vccd1 vccd1 _10885_/B sky130_fd_sc_hd__o21bai_2
X_13667_ hold51/X _13666_/X fanout1/X vssd1 vssd1 vccd1 vccd1 _21865_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_144_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13132__A _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12674__C _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15406_ _15406_/A _15406_/B vssd1 vssd1 vccd1 vccd1 _15417_/A sky130_fd_sc_hd__or2_1
XFILLER_0_143_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19174_ _19174_/A _19174_/B vssd1 vssd1 vccd1 vccd1 _19318_/A sky130_fd_sc_hd__or2_1
X_12618_ _13682_/C _13573_/D _12514_/B _12512_/X vssd1 vssd1 vccd1 vccd1 _12627_/A
+ sky130_fd_sc_hd__a31o_1
X_16386_ _16273_/A _16391_/B _16270_/X _16271_/X _16177_/B vssd1 vssd1 vccd1 vccd1
+ _16387_/B sky130_fd_sc_hd__a32o_1
XANTENNA__15050__C _15050_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13598_ _13444_/A _13444_/B _13443_/B vssd1 vssd1 vccd1 vccd1 _13600_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18125_ _18126_/A _18126_/B vssd1 vssd1 vccd1 vccd1 _18125_/Y sky130_fd_sc_hd__nand2_1
X_15337_ _15430_/B _15336_/C _15336_/A vssd1 vssd1 vccd1 vccd1 _15338_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12549_ _12456_/A _12455_/A _12455_/B vssd1 vssd1 vccd1 vccd1 _12556_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_14_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_937 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18056_ _18057_/A _18057_/B vssd1 vssd1 vccd1 vccd1 _18181_/B sky130_fd_sc_hd__nand2_1
XANTENNA_1 _21721_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19429__A1 _17324_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15268_ _15268_/A _15268_/B vssd1 vssd1 vccd1 vccd1 _15270_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_41_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19429__B2 _19430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17973__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17007_ _16961_/Y _16963_/X _17005_/B _17005_/Y vssd1 vssd1 vccd1 vccd1 _17007_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__11587__A _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14219_ _14220_/A _14220_/B _14220_/C vssd1 vssd1 vccd1 vccd1 _14222_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_112_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15199_ _15199_/A _15199_/B vssd1 vssd1 vccd1 vccd1 _15200_/B sky130_fd_sc_hd__and2_1
Xfanout508 _21742_/Q vssd1 vssd1 vccd1 vccd1 _14367_/A sky130_fd_sc_hd__clkbuf_8
Xfanout519 _21740_/Q vssd1 vssd1 vccd1 vccd1 _14508_/A sky130_fd_sc_hd__buf_4
XFILLER_0_6_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18958_ _19445_/A _19587_/A _20249_/B vssd1 vssd1 vccd1 vccd1 _18958_/X sky130_fd_sc_hd__and3_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17909_ _18026_/B _17908_/C _17908_/A vssd1 vssd1 vccd1 vccd1 _17910_/C sky130_fd_sc_hd__a21o_1
X_18889_ _18889_/A _18889_/B _18889_/C vssd1 vssd1 vccd1 vccd1 _18987_/A sky130_fd_sc_hd__and3_1
X_20920_ _20920_/A _20920_/B vssd1 vssd1 vccd1 vccd1 _20960_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__14977__A1 _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20851_ _20852_/A _20852_/B vssd1 vssd1 vccd1 vccd1 _20851_/Y sky130_fd_sc_hd__nand2_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18168__A1 _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout164_A _21829_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20782_ _20913_/A _20783_/B vssd1 vssd1 vccd1 vccd1 _20784_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11255__A3 fanout19/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11660__B1 _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout331_A _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14138__A _14138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout429_A _21763_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13401__A1 _13554_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13401__B2 _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21403_ hold185/X _21402_/X _21403_/S vssd1 vssd1 vccd1 vccd1 _21942_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_32_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17143__A2 _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21334_ _21407_/S _21334_/B vssd1 vssd1 vccd1 vccd1 _21334_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_142_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18891__A2 _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13704__A2 _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21265_ _21265_/A _21265_/B vssd1 vssd1 vccd1 vccd1 _21266_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19664__A _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12912__B1 _13913_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_1143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1034 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20216_ _20216_/A _20216_/B vssd1 vssd1 vccd1 vccd1 _20218_/B sky130_fd_sc_hd__nor2_1
XANTENNA__16103__B1 _16418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21196_ _21195_/B _21196_/B vssd1 vssd1 vccd1 vccd1 _21197_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_99_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11647__D _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20147_ _20148_/C _20924_/A _20145_/Y _20281_/A vssd1 vssd1 vccd1 vccd1 _20149_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_95_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout77_A _21848_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20078_ _20078_/A _20078_/B vssd1 vssd1 vccd1 vccd1 _20079_/B sky130_fd_sc_hd__nand2_1
XTAP_3402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17334__D _17443_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11920_ _12094_/A _12637_/B _12639_/A _12094_/B vssd1 vssd1 vccd1 vccd1 _11922_/A
+ sky130_fd_sc_hd__a22oi_2
XTAP_3435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11851_ _12267_/A _12751_/B _12637_/B _12242_/B vssd1 vssd1 vccd1 vccd1 _11851_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_3479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ hold51/A hold151/A vssd1 vssd1 vccd1 vccd1 _10802_/X sky130_fd_sc_hd__or2_1
X_14570_ _14567_/X _14568_/Y _14418_/A _14418_/B vssd1 vssd1 vccd1 vccd1 _14571_/B
+ sky130_fd_sc_hd__a211oi_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18446__C _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_1261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21153__B _21153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11782_ _11781_/B _11781_/C _11781_/A vssd1 vssd1 vccd1 vccd1 _11784_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_138_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13521_ _13518_/C _13365_/X _13518_/D _13520_/Y vssd1 vssd1 vccd1 vccd1 _14293_/A
+ sky130_fd_sc_hd__o31ai_4
XFILLER_0_27_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19108__B1 _19751_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11171__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16240_ _16347_/A _16240_/B _16348_/B _16240_/D vssd1 vssd1 vccd1 vccd1 _16347_/B
+ sky130_fd_sc_hd__nor4_2
X_13452_ _13299_/X _13301_/X _13450_/X _13451_/Y vssd1 vssd1 vccd1 vccd1 _13491_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_137_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18462__B _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12403_ _12403_/A _12403_/B _12858_/C _12991_/D vssd1 vssd1 vccd1 vccd1 _12403_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_141_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20269__A2 _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16171_ _16171_/A _16171_/B vssd1 vssd1 vccd1 vccd1 _16181_/A sky130_fd_sc_hd__or2_1
X_13383_ _13384_/A _13384_/B vssd1 vssd1 vccd1 vccd1 _13383_/X sky130_fd_sc_hd__or2_1
XFILLER_0_36_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_959 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15122_ _15122_/A _15266_/B _15122_/C vssd1 vssd1 vccd1 vccd1 _15328_/A sky130_fd_sc_hd__nand3_2
X_12334_ _12334_/A _12334_/B vssd1 vssd1 vccd1 vccd1 _12336_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13156__B1 _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15053_ _14893_/A _14893_/B _14891_/X vssd1 vssd1 vccd1 vccd1 _15055_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_121_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19930_ _19773_/A _19773_/B _19771_/Y vssd1 vssd1 vccd1 vccd1 _19932_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_32_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12265_ _12264_/A _12264_/B _12264_/C vssd1 vssd1 vccd1 vccd1 _12267_/D sky130_fd_sc_hd__a21o_1
XANTENNA__19574__A _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14004_ _13993_/Y _14004_/B _14004_/C vssd1 vssd1 vccd1 vccd1 _14004_/X sky130_fd_sc_hd__and3b_2
X_11216_ _15234_/C _11215_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21755_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_103_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19861_ _19740_/B _19740_/C _19740_/D _19726_/X vssd1 vssd1 vccd1 vccd1 _19863_/C
+ sky130_fd_sc_hd__a31o_1
X_12196_ _12229_/A _12269_/C _12269_/D _12155_/B vssd1 vssd1 vccd1 vccd1 _12197_/B
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__11557__D _12751_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18812_ _18813_/A _18813_/B _18813_/C vssd1 vssd1 vccd1 vccd1 _18812_/X sky130_fd_sc_hd__and3_1
X_11147_ _12530_/A _11146_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21732_/D sky130_fd_sc_hd__mux2_1
X_19792_ _20081_/A _19792_/B vssd1 vssd1 vccd1 vccd1 _21387_/B sky130_fd_sc_hd__xor2_2
XANTENNA__14656__B1 _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18743_ _18739_/X _18741_/Y _18584_/X _18587_/B vssd1 vssd1 vccd1 vccd1 _18744_/B
+ sky130_fd_sc_hd__a211o_1
X_15955_ _16089_/A vssd1 vssd1 vccd1 vccd1 _15957_/D sky130_fd_sc_hd__inv_2
X_11078_ _10926_/X hold52/X _11087_/S vssd1 vssd1 vccd1 vccd1 _21673_/D sky130_fd_sc_hd__mux2_1
X_14906_ _14906_/A _14906_/B vssd1 vssd1 vccd1 vccd1 _14909_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__12669__C _12780_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18674_ _18674_/A _18674_/B _18674_/C _18674_/D vssd1 vssd1 vccd1 vccd1 _18674_/X
+ sky130_fd_sc_hd__or4_1
X_15886_ _16016_/B _16016_/C vssd1 vssd1 vccd1 vccd1 _15888_/A sky130_fd_sc_hd__or2_1
XFILLER_0_76_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17625_ _17749_/A _17625_/B vssd1 vssd1 vccd1 vccd1 _17627_/B sky130_fd_sc_hd__and2_1
XFILLER_0_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14837_ _14840_/B vssd1 vssd1 vccd1 vccd1 _14837_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_148_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17556_ _19445_/A _17924_/B vssd1 vssd1 vccd1 vccd1 _17559_/A sky130_fd_sc_hd__and2_1
XFILLER_0_59_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14768_ _15155_/C _15159_/D _15829_/C _15954_/D vssd1 vssd1 vccd1 vccd1 _14769_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__16157__B _16377_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16507_ _17144_/A _16734_/B _17526_/B _17223_/A vssd1 vssd1 vccd1 vccd1 _16507_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_74_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13719_ _13846_/B _13719_/B vssd1 vssd1 vccd1 vccd1 _13734_/A sky130_fd_sc_hd__and2_1
X_17487_ _17487_/A _17487_/B vssd1 vssd1 vccd1 vccd1 _17489_/B sky130_fd_sc_hd__nor2_1
X_14699_ _14702_/D vssd1 vssd1 vccd1 vccd1 _14699_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_39_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19226_ _19686_/A _19382_/A _19227_/C _19227_/D vssd1 vssd1 vccd1 vccd1 _19226_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_116_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16438_ _16363_/A hold187/X _12291_/B _16437_/Y vssd1 vssd1 vccd1 vccd1 _16438_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15308__A_N _21734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_1067 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19157_ _19157_/A _19157_/B vssd1 vssd1 vccd1 vccd1 _19159_/B sky130_fd_sc_hd__xor2_2
X_16369_ _16369_/A _16369_/B vssd1 vssd1 vccd1 vccd1 _16370_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_54_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16173__A _16173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17125__A2 _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18108_ _18005_/A _18004_/B _18004_/A vssd1 vssd1 vccd1 vccd1 _18119_/A sky130_fd_sc_hd__o21ba_1
X_19088_ _19088_/A _19088_/B vssd1 vssd1 vccd1 vccd1 _19090_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_124_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16884__A1 _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18039_ _18175_/B _18038_/B _18038_/C vssd1 vssd1 vccd1 vccd1 _18040_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_112_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__16884__B2 _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21050_ _21050_/A _21050_/B vssd1 vssd1 vccd1 vccd1 _21052_/B sky130_fd_sc_hd__xor2_1
XANTENNA__19822__A1 _19823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout305 _21794_/Q vssd1 vssd1 vccd1 vccd1 _17504_/C sky130_fd_sc_hd__clkbuf_8
Xfanout316 _17854_/B vssd1 vssd1 vccd1 vccd1 _19008_/D sky130_fd_sc_hd__buf_4
XANTENNA__16620__B _17434_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19822__B2 _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11173__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20001_ _20001_/A _20001_/B vssd1 vssd1 vccd1 vccd1 _20009_/A sky130_fd_sc_hd__nand2_1
Xfanout327 _16406_/B vssd1 vssd1 vccd1 vccd1 _15838_/B sky130_fd_sc_hd__clkbuf_4
Xfanout338 _15174_/D vssd1 vssd1 vccd1 vccd1 _15978_/B sky130_fd_sc_hd__buf_4
Xfanout349 _16377_/A vssd1 vssd1 vccd1 vccd1 _15788_/B sky130_fd_sc_hd__buf_4
XANTENNA__13682__D _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14140__B _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout281_A _18008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout379_A _14828_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11256__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21952_ _21963_/CLK _21952_/D vssd1 vssd1 vccd1 vccd1 hold222/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__19050__A2 _19051_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19650__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_32_clk_i_A clkbuf_2_2__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17597__C1 _11553_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20903_ _20903_/A _20903_/B _20641_/B vssd1 vssd1 vccd1 vccd1 _20904_/D sky130_fd_sc_hd__or3b_2
XANTENNA__18547__B _19181_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21883_ _21949_/CLK hold129/X vssd1 vssd1 vccd1 vccd1 hold128/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12876__A _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout546_A _21734_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20834_ _21016_/A _20834_/B vssd1 vssd1 vccd1 vccd1 _20885_/A sky130_fd_sc_hd__nor2_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__19889__A1 _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19889__B2 _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20765_ _20896_/B _20764_/X _20634_/Y _20638_/A vssd1 vssd1 vccd1 vccd1 _20903_/A
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11930__D _12621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19378__B _19379_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20696_ _20696_/A _20696_/B vssd1 vssd1 vccd1 vccd1 _20698_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14018__D _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__20317__B _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21317_ _21317_/A _21317_/B vssd1 vssd1 vccd1 vccd1 _21318_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_60_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12050_ _12050_/A _12050_/B _12050_/C vssd1 vssd1 vccd1 vccd1 _12102_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_130_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21248_ _21248_/A _21248_/B vssd1 vssd1 vccd1 vccd1 _21248_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__20333__A _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11001_ mstream_o[75] hold27/X _11012_/S vssd1 vssd1 vccd1 vccd1 _21612_/D sky130_fd_sc_hd__mux2_1
XANTENNA__11164__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11955__A _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21179_ _21179_/A _21179_/B vssd1 vssd1 vccd1 vccd1 _21180_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11674__B _12877_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1096 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18738__A _19531_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13310__B1 _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15740_ _15741_/A _15741_/B _15741_/C _15741_/D vssd1 vssd1 vccd1 vccd1 _15740_/Y
+ sky130_fd_sc_hd__nor4_1
XANTENNA__15850__A2 _16396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__17642__A _19823_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12952_ _12952_/A _12952_/B vssd1 vssd1 vccd1 vccd1 _17834_/B sky130_fd_sc_hd__xor2_4
XTAP_3232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20463__A1_N _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11903_ _11894_/X _11901_/X _11902_/X _11836_/Y vssd1 vssd1 vccd1 vccd1 _11905_/A
+ sky130_fd_sc_hd__o211a_1
X_15671_ _15931_/B _14698_/D _16391_/B _15931_/A vssd1 vssd1 vccd1 vccd1 _15675_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_3265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_210 hold275/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ _13157_/A _13155_/C _13155_/D _14024_/B vssd1 vssd1 vccd1 vccd1 _12884_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA_221 hold277/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_232 hold299/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17410_ _17487_/A _17409_/C _17409_/A vssd1 vssd1 vccd1 vccd1 _17470_/B sky130_fd_sc_hd__o21a_1
XTAP_3298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14622_ _14624_/A vssd1 vssd1 vccd1 vccd1 _14782_/A sky130_fd_sc_hd__inv_2
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_243 _11347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18390_ _18390_/A _18394_/C vssd1 vssd1 vccd1 vccd1 _18390_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA_254 v2z[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11834_ _11834_/A _11834_/B vssd1 vssd1 vccd1 vccd1 _11836_/B sky130_fd_sc_hd__nor2_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14810__B1 _15112_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_265 hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_276 v0z[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_1080 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_287 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17341_ _17340_/B _17340_/C _17340_/A vssd1 vssd1 vccd1 vccd1 _17343_/B sky130_fd_sc_hd__a21o_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_298 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14553_ _14553_/A _14553_/B vssd1 vssd1 vccd1 vccd1 _14580_/A sky130_fd_sc_hd__nor2_2
X_11765_ _11764_/B _11764_/C _11764_/A vssd1 vssd1 vccd1 vccd1 _11767_/B sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13504_ _13353_/B _13353_/Y _13500_/X _13502_/Y vssd1 vssd1 vccd1 vccd1 _13504_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_153_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17272_ _21142_/A _12392_/B _21334_/B _20770_/B vssd1 vssd1 vccd1 vccd1 _17272_/X
+ sky130_fd_sc_hd__o22a_1
X_14484_ _14473_/Y _14484_/B _14484_/C vssd1 vssd1 vccd1 vccd1 _14647_/A sky130_fd_sc_hd__and3b_1
XANTENNA__13113__C _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11696_ _11640_/A _11640_/B _11640_/C vssd1 vssd1 vccd1 vccd1 _11697_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19011_ _19011_/A vssd1 vssd1 vccd1 vccd1 _19021_/A sky130_fd_sc_hd__inv_2
XFILLER_0_67_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16223_ _16223_/A _16223_/B vssd1 vssd1 vccd1 vccd1 _16224_/B sky130_fd_sc_hd__or2_1
X_13435_ _14195_/A _14384_/A _14212_/B _13875_/B vssd1 vssd1 vccd1 vccd1 _13437_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16154_ _16391_/A _16414_/A _16268_/B _16266_/C vssd1 vssd1 vccd1 vccd1 _16324_/A
+ sky130_fd_sc_hd__and4_1
X_13366_ _13518_/A _13518_/B vssd1 vssd1 vccd1 vccd1 _13366_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15105_ _15004_/B _15006_/B _15254_/A _15104_/Y vssd1 vssd1 vccd1 vccd1 _15254_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_11_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12317_ _12317_/A _12317_/B vssd1 vssd1 vccd1 vccd1 _12379_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__15853__A2_N _15978_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16085_ _16201_/A vssd1 vssd1 vccd1 vccd1 _16087_/D sky130_fd_sc_hd__inv_2
X_13297_ _13445_/B _13297_/B vssd1 vssd1 vccd1 vccd1 _13300_/A sky130_fd_sc_hd__nor2_1
XANTENNA__11568__C _12528_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15036_ _15035_/B _15127_/B _15035_/A vssd1 vssd1 vccd1 vccd1 _15037_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_48_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19913_ _19708_/A _19708_/C _19708_/B vssd1 vssd1 vccd1 vccd1 _19914_/C sky130_fd_sc_hd__a21bo_1
X_12248_ _12784_/A _21727_/Q _12249_/C _12249_/D vssd1 vssd1 vccd1 vccd1 _12248_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_20_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11155__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12352__A1 _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12352__B2 _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19844_ _19847_/A _19847_/B _19844_/C vssd1 vssd1 vccd1 vccd1 _19961_/A sky130_fd_sc_hd__and3_2
XFILLER_0_120_1230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__21058__B _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12179_ _12139_/A _12139_/C _12139_/B vssd1 vssd1 vccd1 vccd1 _12185_/B sky130_fd_sc_hd__a21o_1
XANTENNA__19280__A2 _19753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19775_ _19776_/B _19776_/A vssd1 vssd1 vccd1 vccd1 _19775_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__19751__B _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16987_ _17029_/A _17029_/B _17145_/B _17146_/C vssd1 vssd1 vccd1 vccd1 _16990_/A
+ sky130_fd_sc_hd__and4_1
X_18726_ _18847_/A _18725_/C _18725_/A vssd1 vssd1 vccd1 vccd1 _18726_/X sky130_fd_sc_hd__o21a_1
XANTENNA__17552__A _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15938_ _15938_/A _15938_/B vssd1 vssd1 vccd1 vccd1 _15940_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18657_ _18656_/A _18656_/B _18656_/C vssd1 vssd1 vccd1 vccd1 _18658_/C sky130_fd_sc_hd__a21o_1
X_15869_ _15687_/B _15689_/B _15952_/B _15868_/Y vssd1 vssd1 vccd1 vccd1 _15870_/A
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_78_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17608_ _19337_/D _18851_/C _20797_/A _21258_/A vssd1 vssd1 vccd1 vccd1 _17732_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18588_ _18588_/A _18588_/B vssd1 vssd1 vccd1 vccd1 _18590_/B sky130_fd_sc_hd__or2_1
XFILLER_0_47_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17539_ _17535_/X _17536_/Y _17422_/X _17424_/X vssd1 vssd1 vccd1 vccd1 _17575_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_4_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11615__B1 _12991_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_156_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20550_ _21256_/A _20924_/A _20550_/C _20550_/D vssd1 vssd1 vccd1 vccd1 _20679_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__15357__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_818 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1099 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19209_ _19363_/A _19207_/Y _19035_/B _19037_/B vssd1 vssd1 vccd1 vccd1 _19210_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_105_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20481_ _20481_/A _20481_/B vssd1 vssd1 vccd1 vccd1 _20483_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout127_A _20910_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13320__A _14712_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20102__A1 _20103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21102_ _21296_/A _21311_/B _21102_/C _21102_/D vssd1 vssd1 vccd1 vccd1 _21208_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_11_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22082_ _22096_/CLK _22082_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[18] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_11_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11146__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout496_A _16404_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout102 _21841_/Q vssd1 vssd1 vccd1 vccd1 _21258_/A sky130_fd_sc_hd__buf_6
X_21033_ _21033_/A _21033_/B vssd1 vssd1 vccd1 vccd1 _21034_/B sky130_fd_sc_hd__xor2_2
Xfanout113 _17741_/B vssd1 vssd1 vccd1 vccd1 _21171_/A sky130_fd_sc_hd__buf_4
Xfanout124 _19906_/A vssd1 vssd1 vccd1 vccd1 _19068_/C sky130_fd_sc_hd__buf_4
Xfanout135 _21835_/Q vssd1 vssd1 vccd1 vccd1 _19087_/B sky130_fd_sc_hd__buf_4
Xfanout146 _21832_/Q vssd1 vssd1 vccd1 vccd1 _17417_/D sky130_fd_sc_hd__buf_2
Xfanout157 _20088_/A vssd1 vssd1 vccd1 vccd1 _18789_/A sky130_fd_sc_hd__clkbuf_8
Xfanout168 _19732_/A vssd1 vssd1 vccd1 vccd1 _19430_/A sky130_fd_sc_hd__clkbuf_4
Xfanout179 _17443_/D vssd1 vssd1 vccd1 vccd1 _19438_/B sky130_fd_sc_hd__buf_4
XANTENNA__20169__A1 _20590_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20169__B2 _20462_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17181__B _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21935_ _21938_/CLK _21935_/D vssd1 vssd1 vccd1 vccd1 hold111/A sky130_fd_sc_hd__dfxtp_1
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16509__C _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold241_A hold241/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21866_ _21948_/CLK hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_78_962 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20817_ _20817_/A _20817_/B vssd1 vssd1 vccd1 vccd1 _20819_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21797_ _21803_/CLK _21797_/D vssd1 vssd1 vccd1 vccd1 _21797_/Q sky130_fd_sc_hd__dfxtp_1
XANTENNA__15132__D _16328_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_1189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19731__B1 _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11550_ _11550_/A _11550_/B vssd1 vssd1 vccd1 vccd1 fanout8/A sky130_fd_sc_hd__nor2_1
XFILLER_0_9_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20748_ _20747_/B _20747_/C _20747_/A vssd1 vssd1 vccd1 vccd1 _20748_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout6_A fanout6/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_615 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11481_ _11502_/A1 t2x[10] v1z[10] fanout20/X _11480_/X vssd1 vssd1 vccd1 vccd1 _11481_/X
+ sky130_fd_sc_hd__a221o_1
X_20679_ _20679_/A _20679_/B vssd1 vssd1 vccd1 vccd1 _20681_/B sky130_fd_sc_hd__or2_1
XANTENNA__14326__A _15155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13220_ _13080_/Y _13083_/X _13217_/X _13219_/Y vssd1 vssd1 vccd1 vccd1 _13361_/A
+ sky130_fd_sc_hd__a211o_2
XANTENNA__18740__B _19382_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11385__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ _14024_/B _13152_/C _12420_/D _14027_/A vssd1 vssd1 vccd1 vccd1 _13153_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17637__A _18008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16541__A _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12102_ _12102_/A _12102_/B _12102_/C vssd1 vssd1 vccd1 vccd1 _12115_/A sky130_fd_sc_hd__and3_2
XANTENNA__14323__A2 _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13082_ _13083_/A _13083_/B _13083_/C vssd1 vssd1 vccd1 vccd1 _13085_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_27_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11137__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16910_ _17168_/A _17168_/B _17167_/A _17167_/B vssd1 vssd1 vccd1 vccd1 _16912_/A
+ sky130_fd_sc_hd__and4bb_1
X_12033_ _11905_/Y _11910_/X _11976_/A _11977_/X vssd1 vssd1 vccd1 vccd1 _12294_/D
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__19852__A _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17890_ _17975_/B _17890_/B vssd1 vssd1 vccd1 vccd1 _17953_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16841_ _16834_/Y _16837_/Y _16849_/B _16840_/X vssd1 vssd1 vccd1 vccd1 _16849_/C
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__19571__B _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_19560_ _19560_/A _19560_/B _19560_/C vssd1 vssd1 vccd1 vccd1 _19562_/A sky130_fd_sc_hd__and3_1
X_16772_ _16773_/A _16773_/B _16773_/C vssd1 vssd1 vccd1 vccd1 _16783_/A sky130_fd_sc_hd__a21o_1
X_13984_ _13985_/A _16374_/B _13985_/C _13985_/D vssd1 vssd1 vccd1 vccd1 _13986_/A
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_88_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18511_ _18511_/A _18511_/B _18511_/C vssd1 vssd1 vccd1 vccd1 _18511_/Y sky130_fd_sc_hd__nand3_2
X_15723_ _15724_/A _15724_/B vssd1 vssd1 vccd1 vccd1 _15723_/Y sky130_fd_sc_hd__nand2_1
XTAP_3040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1191 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19491_ _20838_/C _19331_/X _19334_/A _19334_/B vssd1 vssd1 vccd1 vccd1 _19492_/B
+ sky130_fd_sc_hd__o2bb2a_2
X_12935_ _12971_/B _12934_/B _12934_/C _12934_/D vssd1 vssd1 vccd1 vccd1 _12935_/Y
+ sky130_fd_sc_hd__a22oi_4
XFILLER_0_88_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1033 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18442_ _18442_/A _18442_/B vssd1 vssd1 vccd1 vccd1 _18451_/A sky130_fd_sc_hd__or2_1
X_15654_ _16404_/A _15913_/B _15655_/C _15849_/A vssd1 vssd1 vccd1 vccd1 _15656_/A
+ sky130_fd_sc_hd__a22o_1
XTAP_3095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ _12868_/A _12868_/B _12868_/C vssd1 vssd1 vccd1 vccd1 _12866_/Y sky130_fd_sc_hd__a21oi_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_984 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14605_ fanout9/X _14605_/B vssd1 vssd1 vccd1 vccd1 _14605_/Y sky130_fd_sc_hd__nor2_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18373_ _18373_/A _18373_/B _18373_/C _18373_/D vssd1 vssd1 vccd1 vccd1 _18373_/X
+ sky130_fd_sc_hd__or4_2
XFILLER_0_8_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11817_ _11816_/B _11816_/C _11816_/A vssd1 vssd1 vccd1 vccd1 _11819_/B sky130_fd_sc_hd__a21bo_1
X_15585_ _15585_/A _15585_/B vssd1 vssd1 vccd1 vccd1 _15586_/B sky130_fd_sc_hd__xnor2_2
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ _12798_/A _12798_/B _12798_/C vssd1 vssd1 vccd1 vccd1 _12797_/X sky130_fd_sc_hd__and3_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17324_ _17434_/B _17433_/A _19430_/A _17324_/D vssd1 vssd1 vccd1 vccd1 _17324_/X
+ sky130_fd_sc_hd__and4_1
X_14536_ _16326_/A _14535_/X _14534_/X vssd1 vssd1 vccd1 vccd1 _14538_/A sky130_fd_sc_hd__a21bo_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11748_ _11748_/A _11748_/B _11748_/C vssd1 vssd1 vccd1 vccd1 _11767_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_55_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17255_ _17256_/A _17256_/B _17256_/C _17256_/D vssd1 vssd1 vccd1 vccd1 _17255_/Y
+ sky130_fd_sc_hd__nor4_1
X_14467_ _14467_/A _14467_/B vssd1 vssd1 vccd1 vccd1 _14469_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_148_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14236__A _14859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13778__C _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ _12229_/A _12155_/B _12642_/A _12751_/B vssd1 vssd1 vccd1 vccd1 _11705_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_153_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16206_ _16206_/A _16206_/B vssd1 vssd1 vccd1 vccd1 _16207_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_141_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13418_ _14027_/A _13864_/B _14516_/A _14365_/C vssd1 vssd1 vccd1 vccd1 _13569_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_10_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17186_ _17187_/A _17186_/B _17185_/B vssd1 vssd1 vccd1 vccd1 _17186_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_148_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14398_ _14398_/A _14532_/B _14398_/C vssd1 vssd1 vccd1 vccd1 _14398_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_3_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19746__B _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11376__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16137_ _15968_/B _15970_/Y _16251_/A _16136_/X vssd1 vssd1 vccd1 vccd1 _16251_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13349_ _13348_/B _13348_/C _13348_/A vssd1 vssd1 vccd1 vccd1 _13349_/Y sky130_fd_sc_hd__o21ai_2
XFILLER_0_51_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16451__A _17029_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16068_ _16069_/A _16069_/B _16069_/C vssd1 vssd1 vccd1 vccd1 _16070_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_121_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11128__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15019_ _15019_/A _15019_/B vssd1 vssd1 vccd1 vccd1 _15028_/A sky130_fd_sc_hd__xnor2_2
XANTENNA__10887__A1 _10886_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18461__B1 _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19827_ _19826_/B _20043_/B _19826_/A vssd1 vssd1 vccd1 vccd1 _19828_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_120_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17282__A _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13018__C _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19758_ _19758_/A _19758_/B _19758_/C vssd1 vssd1 vccd1 vccd1 _19759_/A sky130_fd_sc_hd__and3_1
XFILLER_0_155_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18709_ _18709_/A _18709_/B vssd1 vssd1 vccd1 vccd1 _18718_/A sky130_fd_sc_hd__or2_1
XANTENNA__15514__B _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19689_ _19689_/A _19689_/B vssd1 vssd1 vccd1 vccd1 _19699_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_151_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_1129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21720_ _21934_/CLK _21720_/D _11041_/A vssd1 vssd1 vccd1 vccd1 _21720_/Q sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_921 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21651_ _22063_/CLK _21651_/D _21422_/A vssd1 vssd1 vccd1 vccd1 mstream_o[115] sky130_fd_sc_hd__dfrtp_4
XANTENNA__13034__B _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout244_A _21807_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20602_ _20602_/A _20602_/B vssd1 vssd1 vccd1 vccd1 _20613_/A sky130_fd_sc_hd__or2_1
XFILLER_0_75_965 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19002__A _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21520__A0 hold258/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21582_ _22106_/CLK _21582_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[45] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_1073 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20533_ _20533_/A _20533_/B vssd1 vssd1 vccd1 vccd1 _20535_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout411_A _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout509_A _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20464_ _20600_/A _20464_/B vssd1 vssd1 vccd1 vccd1 _20465_/B sky130_fd_sc_hd__nor2_1
XANTENNA__11367__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13985__A _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_1213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20395_ _19972_/A _20394_/B _20247_/D vssd1 vssd1 vccd1 vccd1 _20396_/B sky130_fd_sc_hd__o21a_1
XANTENNA__14305__A2 _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22065_ _22069_/CLK _22065_/D fanout639/X vssd1 vssd1 vccd1 vccd1 mstream_o[1] sky130_fd_sc_hd__dfrtp_4
XANTENNA__16511__D _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14312__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21016_ _21016_/A _21016_/B _21016_/C vssd1 vssd1 vccd1 vccd1 _21016_/Y sky130_fd_sc_hd__nor3_1
XANTENNA__17192__A _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1017 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13816__A1 _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13816__B2 fanout5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11952__B _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10981_ hold92/A hold171/A vssd1 vssd1 vccd1 vccd1 _10982_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_30_clk_i clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 _21948_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA__17558__A2 _17670_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19952__B1 _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13225__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12720_ _13983_/B _13394_/A _14176_/C _13402_/D vssd1 vssd1 vccd1 vccd1 _12834_/A
+ sky130_fd_sc_hd__and4_2
XANTENNA__15569__A1 _15426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21918_ _21926_/CLK _21918_/D vssd1 vssd1 vccd1 vccd1 hold156/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_139_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16766__B1 _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12651_ _12651_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _12653_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__14241__A1 _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21849_ _21853_/CLK _21849_/D vssd1 vssd1 vccd1 vccd1 _21849_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_155_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14241__B2 _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11602_ _11602_/A _11602_/B vssd1 vssd1 vccd1 vccd1 _11887_/A sky130_fd_sc_hd__xor2_1
X_15370_ _16027_/A _15370_/B _15370_/C _15548_/A vssd1 vssd1 vccd1 vccd1 _15548_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_26_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12582_ _12583_/A _12583_/B _12583_/C _12583_/D vssd1 vssd1 vccd1 vccd1 _12582_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19180__A1 _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14321_ _14321_/A _14321_/B vssd1 vssd1 vccd1 vccd1 _14341_/A sky130_fd_sc_hd__xor2_4
XFILLER_0_93_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11533_ _11532_/X _19013_/C _11545_/S vssd1 vssd1 vccd1 vccd1 _21849_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_81_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18751__A _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13595__A2_N _15763_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_1_clk_i_A _21822_/CLK vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17040_ _17028_/Y _17038_/X _16994_/Y _17010_/X vssd1 vssd1 vccd1 vccd1 _17040_/X
+ sky130_fd_sc_hd__a211o_1
X_14252_ _14251_/A _14251_/B _14251_/C vssd1 vssd1 vccd1 vccd1 _14254_/C sky130_fd_sc_hd__a21oi_1
X_11464_ _11463_/X _17443_/D _11470_/S vssd1 vssd1 vccd1 vccd1 _21826_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_40_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19566__B _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11358__A2 fanout29/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13895__A _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13203_ _13204_/A _13204_/B _13204_/C vssd1 vssd1 vccd1 vccd1 _13203_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_150_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14183_ _14659_/A _15022_/B _14185_/C _14185_/D vssd1 vssd1 vccd1 vccd1 _14183_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11395_ _11394_/X _17434_/B _11401_/S vssd1 vssd1 vccd1 vccd1 _21803_/D sky130_fd_sc_hd__mux2_1
XANTENNA__16271__A _16380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17494__A1 _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13134_ _13134_/A _13267_/B _13134_/C vssd1 vssd1 vccd1 vccd1 _13136_/B sky130_fd_sc_hd__nand3_1
X_18991_ _18991_/A _18991_/B _18991_/C vssd1 vssd1 vccd1 vccd1 _19155_/B sky130_fd_sc_hd__or3_1
XANTENNA__17086__B _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ _13061_/X _13063_/Y _12924_/B _12924_/Y vssd1 vssd1 vccd1 vccd1 _13067_/C
+ sky130_fd_sc_hd__o211a_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17942_ _17943_/A _17943_/B _17943_/C vssd1 vssd1 vccd1 vccd1 _17942_/X sky130_fd_sc_hd__and3_1
X_12016_ _12017_/A _12017_/B vssd1 vssd1 vccd1 vccd1 _12036_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__21042__A2 _21278_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18443__B1 _19238_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13119__B _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17873_ _18008_/B _19906_/A _20146_/B _18010_/A vssd1 vssd1 vccd1 vccd1 _17874_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19732__D _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16824_ _16754_/A _16754_/B _16754_/C vssd1 vssd1 vccd1 vccd1 _16824_/X sky130_fd_sc_hd__a21o_1
X_19612_ _19612_/A _19612_/B vssd1 vssd1 vccd1 vccd1 _19613_/B sky130_fd_sc_hd__xor2_4
XFILLER_0_136_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20722__A2_N _21293_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19543_ _19543_/A _19543_/B vssd1 vssd1 vccd1 vccd1 _19551_/A sky130_fd_sc_hd__nand2_1
XANTENNA__14876__D _16391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16755_ _16705_/A _16705_/B _16705_/C vssd1 vssd1 vccd1 vccd1 _16755_/Y sky130_fd_sc_hd__a21oi_2
X_13967_ _14291_/A _13967_/B vssd1 vssd1 vccd1 vccd1 _13967_/X sky130_fd_sc_hd__xor2_4
XANTENNA__18746__A1 _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15706_ _15706_/A _15706_/B vssd1 vssd1 vccd1 vccd1 _15709_/A sky130_fd_sc_hd__xnor2_2
X_12918_ _12918_/A _12918_/B _12918_/C vssd1 vssd1 vccd1 vccd1 _12921_/A sky130_fd_sc_hd__nand3_2
X_19474_ _19788_/A _19788_/B _19169_/B vssd1 vssd1 vccd1 vccd1 _19475_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_0_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16686_ _16686_/A _16686_/B _16686_/C vssd1 vssd1 vccd1 vccd1 _16686_/X sky130_fd_sc_hd__and3_2
X_13898_ _15514_/A _15514_/B _14212_/D _14218_/B vssd1 vssd1 vccd1 vccd1 _13901_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__21352__A _21412_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18425_ _18542_/A _18423_/X _18269_/Y _18272_/X vssd1 vssd1 vccd1 vccd1 _18525_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_5_1213 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18645__B _19414_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15637_ _15763_/A _16027_/B _15516_/B vssd1 vssd1 vccd1 vccd1 _15770_/A sky130_fd_sc_hd__a21oi_2
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_932 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13035__A2 _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12849_ _13682_/C _14018_/C _12984_/A _12847_/Y vssd1 vssd1 vccd1 vccd1 _12850_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_69_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14232__A1 _14713_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14232__B2 _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_1257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_18356_ _18355_/A _18355_/B _18355_/C vssd1 vssd1 vccd1 vccd1 _18357_/C sky130_fd_sc_hd__a21o_1
X_15568_ _15567_/B _15567_/C _15567_/A vssd1 vssd1 vccd1 vccd1 _15568_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_84_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19171__A1 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17307_ _17525_/A _17520_/A _17417_/C _17417_/D vssd1 vssd1 vccd1 vccd1 _17307_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_154_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14519_ _14519_/A _14519_/B _14671_/B vssd1 vssd1 vccd1 vccd1 _14521_/B sky130_fd_sc_hd__nand3_1
X_18287_ _18287_/A _18287_/B vssd1 vssd1 vccd1 vccd1 _18290_/A sky130_fd_sc_hd__xor2_2
X_15499_ _12291_/B _21399_/B _15498_/X vssd1 vssd1 vccd1 vccd1 _15499_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_86_1235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17182__B1 _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_1246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17721__A2 _19051_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17238_ _17557_/A _17915_/A _17557_/B _17915_/D vssd1 vssd1 vccd1 vccd1 _17240_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_47_1219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_102_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17169_ _17169_/A _17169_/B _17169_/C vssd1 vssd1 vccd1 vccd1 _17169_/X sky130_fd_sc_hd__or3_1
XFILLER_0_24_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_1090 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17485__B2 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20180_ _20328_/A _20180_/B vssd1 vssd1 vccd1 vccd1 _20181_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20431__A _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15525__A _16036_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16996__B1 _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17443__C _17666_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18258__D _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout361_A _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11264__S _11284_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout459_A _21755_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20862__A1_N _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11285__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21703_ _22096_/CLK _21703_/D vssd1 vssd1 vccd1 vccd1 hold144/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_137_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_954 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout626_A _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11037__A1 hold268/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21634_ _21682_/CLK hold259/X fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[97] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13982__B1 _16406_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21565_ mstream_o[28] hold5/X _21579_/S vssd1 vssd1 vccd1 vccd1 _22092_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_145_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15410__D _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20516_ _11550_/A _20514_/Y _20515_/X vssd1 vssd1 vccd1 vccd1 _20516_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_90_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20028__D _20841_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21496_ hold308/X sstream_i[73] _21510_/S vssd1 vssd1 vccd1 vccd1 _22023_/D sky130_fd_sc_hd__mux2_1
XANTENNA__20606__A _21261_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20447_ _20449_/A _20449_/B _20449_/C vssd1 vssd1 vccd1 vccd1 _20450_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_127_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11180_ _13173_/C _11179_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21743_/D sky130_fd_sc_hd__mux2_1
X_20378_ hold95/X fanout7/X _21399_/B _11550_/B _20377_/Y vssd1 vssd1 vccd1 vccd1
+ _20378_/X sky130_fd_sc_hd__a221o_1
XANTENNA__17915__A _17915_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_1139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22048_ _22049_/CLK _22048_/D vssd1 vssd1 vccd1 vccd1 hold239/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__17779__A2 _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15435__A _15435_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14870_ _15632_/B _14217_/D _16268_/B _14993_/A vssd1 vssd1 vccd1 vccd1 _14870_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21156__B _21841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13821_ _13824_/D vssd1 vssd1 vccd1 vccd1 _13821_/Y sky130_fd_sc_hd__inv_2
XANTENNA__15961__A_N _14813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11174__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16540_ _17741_/B _17387_/A vssd1 vssd1 vccd1 vccd1 _16544_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_134_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13752_ _13752_/A _13752_/B vssd1 vssd1 vccd1 vccd1 _13754_/B sky130_fd_sc_hd__or2_1
X_10964_ _10959_/A _10958_/Y _10957_/A vssd1 vssd1 vccd1 vccd1 _10965_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_97_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14993__B _15892_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12703_ _12589_/X _12591_/Y _12701_/Y _12702_/X vssd1 vssd1 vccd1 vccd1 _12947_/A
+ sky130_fd_sc_hd__o211a_1
X_16471_ _16471_/A vssd1 vssd1 vccd1 vccd1 _16472_/D sky130_fd_sc_hd__inv_2
X_13683_ _13556_/D _13557_/B _13681_/X _13835_/B vssd1 vssd1 vccd1 vccd1 _13685_/A
+ sky130_fd_sc_hd__a211o_1
XANTENNA__16266__A _16391_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10895_ hold83/A hold137/A vssd1 vssd1 vccd1 vccd1 _10897_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19495__A1_N _18849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18210_ _18209_/B _18209_/C _18209_/A vssd1 vssd1 vccd1 vccd1 _18212_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_35_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15422_ _15243_/X _15246_/Y _15420_/Y _15421_/X vssd1 vssd1 vccd1 vccd1 _15422_/X
+ sky130_fd_sc_hd__o211a_2
XANTENNA__11028__A1 hold275/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19190_ _19190_/A _19190_/B _19190_/C vssd1 vssd1 vccd1 vccd1 _19192_/A sky130_fd_sc_hd__nor3_1
X_12634_ _12631_/A _12632_/Y _12543_/X _12546_/Y vssd1 vssd1 vccd1 vccd1 _12634_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_155_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18141_ _18288_/B _18140_/B _18140_/C vssd1 vssd1 vccd1 vccd1 _18142_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15353_ _15354_/B _15354_/A vssd1 vssd1 vccd1 vccd1 _15353_/X sky130_fd_sc_hd__and2b_1
XANTENNA__13402__B _13556_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_946 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_1121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12565_ _14248_/A _12785_/B _14386_/B _14384_/C vssd1 vssd1 vccd1 vccd1 _12567_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_0_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14217__C _14873_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14304_ _14208_/A _14208_/B _14207_/A vssd1 vssd1 vccd1 vccd1 _14343_/A sky130_fd_sc_hd__o21ai_4
XFILLER_0_53_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14517__A2 _15808_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11516_ _21723_/D t1y[22] t0x[22] _11223_/A vssd1 vssd1 vccd1 vccd1 _11516_/X sky130_fd_sc_hd__a22o_1
X_18072_ _18071_/B _18071_/C _18071_/A vssd1 vssd1 vccd1 vccd1 _18074_/B sky130_fd_sc_hd__a21o_1
X_15284_ _15284_/A _15284_/B vssd1 vssd1 vccd1 vccd1 _15286_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12496_ _12496_/A _12496_/B _12708_/B vssd1 vssd1 vccd1 vccd1 _12496_/X sky130_fd_sc_hd__or3_1
XFILLER_0_124_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17023_ _17023_/A _17023_/B vssd1 vssd1 vccd1 vccd1 _17025_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_34_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14235_ _14859_/A _15093_/B _14236_/C _14403_/A vssd1 vssd1 vccd1 vccd1 _14237_/B
+ sky130_fd_sc_hd__a22o_1
X_11447_ _11447_/A1 hold148/A fanout48/X hold202/A vssd1 vssd1 vccd1 vccd1 _11447_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_1117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14166_ _14004_/X _14007_/A _14338_/B _14165_/Y vssd1 vssd1 vccd1 vccd1 _14303_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11378_ _11124_/A hold248/X fanout45/X hold183/X vssd1 vssd1 vccd1 vccd1 _11378_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13117_ _13117_/A _13117_/B vssd1 vssd1 vccd1 vccd1 _13127_/A sky130_fd_sc_hd__xnor2_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14097_ _13933_/A _13933_/C _13933_/B vssd1 vssd1 vccd1 vccd1 _14098_/C sky130_fd_sc_hd__a21bo_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18974_ _18975_/A _18975_/B _18975_/C vssd1 vssd1 vccd1 vccd1 _18974_/X sky130_fd_sc_hd__and3_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ _14572_/A _14391_/B vssd1 vssd1 vccd1 vccd1 _13051_/A sky130_fd_sc_hd__and2_1
XANTENNA__16690__A2 _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17925_ _19438_/A _19438_/B _19703_/C _18640_/B vssd1 vssd1 vccd1 vccd1 _17927_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_147_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17856_ _18851_/C _19051_/C _19221_/C _17854_/B vssd1 vssd1 vccd1 vccd1 _17857_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16442__A2 _17223_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16807_ _16806_/B _16806_/C _16806_/A vssd1 vssd1 vccd1 vccd1 _16810_/B sky130_fd_sc_hd__a21bo_1
X_17787_ _19438_/B _17924_/B _17670_/B _19438_/A vssd1 vssd1 vccd1 vccd1 _17787_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_156_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14999_ _15373_/A _15373_/B _15098_/B _15368_/D vssd1 vssd1 vccd1 vccd1 _15001_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_89_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16738_ _16738_/A _16738_/B _16738_/C vssd1 vssd1 vccd1 vccd1 _16810_/A sky130_fd_sc_hd__nand3_1
X_19526_ _19526_/A _19526_/B vssd1 vssd1 vccd1 vccd1 _19621_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19457_ _19457_/A _19457_/B vssd1 vssd1 vccd1 vccd1 _19460_/A sky130_fd_sc_hd__xnor2_2
X_16669_ _16669_/A _16669_/B _16669_/C vssd1 vssd1 vccd1 vccd1 _16701_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_14_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_431 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18408_ _18405_/X _18552_/B _18281_/D _18282_/B vssd1 vssd1 vccd1 vccd1 _18409_/B
+ sky130_fd_sc_hd__o211ai_1
XANTENNA__12216__B1 _12246_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19388_ _19258_/A _19260_/B _19258_/B vssd1 vssd1 vccd1 vccd1 _19393_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_57_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__15953__B2 _16203_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_924 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14408__B _15091_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18339_ _18339_/A _18481_/B vssd1 vssd1 vccd1 vccd1 _18341_/B sky130_fd_sc_hd__or2_1
XFILLER_0_56_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16326__D _16418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19487__A _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18391__A _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21350_ _21407_/S _17834_/B _21403_/S vssd1 vssd1 vccd1 vccd1 _21350_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20301_ _20301_/A _20301_/B vssd1 vssd1 vccd1 vccd1 _20302_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__11990__A2 _12639_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21281_ _21281_/A _21281_/B vssd1 vssd1 vccd1 vccd1 _21322_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_12_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout4 fanout4/A vssd1 vssd1 vccd1 vccd1 fanout4/X sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout207_A _21816_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20232_ _20237_/A _20094_/B _19961_/A vssd1 vssd1 vccd1 vccd1 _20239_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_60_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_1238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20163_ _20163_/A _20163_/B vssd1 vssd1 vccd1 vccd1 _20166_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_110_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20094_ _20237_/A _20094_/B vssd1 vssd1 vccd1 vccd1 _20097_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_23_1071 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14692__A1 _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout576_A _21727_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14692__B2 _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1036 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11258__A1 _11502_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11258__B2 _11501_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20996_ _20996_/A _20996_/B vssd1 vssd1 vccd1 vccd1 _20997_/B sky130_fd_sc_hd__or2_1
XFILLER_0_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18285__B _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15702__B _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_937 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_902 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout22_A fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_935 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12758__A1 _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21617_ _21906_/CLK _21617_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[80] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_146_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_968 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18732__C _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12350_ _12350_/A _12350_/B vssd1 vssd1 vccd1 vccd1 _12370_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_21548_ mstream_o[11] hold49/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22075_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_117_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11301_ _11325_/A1 t2y[19] t0y[19] _11507_/A1 vssd1 vssd1 vccd1 vccd1 _11301_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_22_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_27_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12281_ _12279_/Y _12280_/X _12239_/X vssd1 vssd1 vccd1 vccd1 _12281_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_65_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21479_ hold130/X sstream_i[56] _21481_/S vssd1 vssd1 vccd1 vccd1 _22006_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12780__C _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14020_ _15155_/C _15112_/D _14020_/C _14020_/D vssd1 vssd1 vccd1 vccd1 _14021_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__17449__A1 _17557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11232_ _12245_/B _11231_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21759_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18646__B1 _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17449__B2 _17557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14053__B _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11163_ hold250/X _11126_/A fanout45/X hold303/A vssd1 vssd1 vccd1 vccd1 _11163_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15971_ _15971_/A _15971_/B vssd1 vssd1 vccd1 vccd1 _15991_/A sky130_fd_sc_hd__xor2_2
X_11094_ _11053_/X hold4/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21688_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_140_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17710_ _17837_/A _17710_/B vssd1 vssd1 vccd1 vccd1 _21346_/B sky130_fd_sc_hd__xor2_4
X_14922_ _14910_/A _14922_/B vssd1 vssd1 vccd1 vccd1 _15069_/A sky130_fd_sc_hd__nand2b_2
XANTENNA__11497__A1 _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12004__D _12403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18690_ hold150/A fanout8/X _21367_/B _11550_/A _18689_/Y vssd1 vssd1 vccd1 vccd1
+ _18690_/X sky130_fd_sc_hd__a221o_1
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold71 hold71/A vssd1 vssd1 vccd1 vccd1 hold71/X sky130_fd_sc_hd__dlygate4sd3_1
X_17641_ _19664_/B _18624_/A vssd1 vssd1 vccd1 vccd1 _17645_/A sky130_fd_sc_hd__nand2_1
Xhold82 hold82/A vssd1 vssd1 vccd1 vccd1 hold82/X sky130_fd_sc_hd__dlygate4sd3_1
X_14853_ _14974_/B _14971_/C _14974_/A _14718_/X vssd1 vssd1 vccd1 vccd1 _14865_/B
+ sky130_fd_sc_hd__a211o_1
Xhold93 hold93/A vssd1 vssd1 vccd1 vccd1 hold93/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13804_ _13819_/B _13804_/B _13802_/Y _13803_/X vssd1 vssd1 vccd1 vccd1 _13804_/X
+ sky130_fd_sc_hd__or4bb_4
XANTENNA__11249__A1 _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11249__B2 _11123_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17572_ _17461_/B _17461_/Y _17569_/X _17571_/Y vssd1 vssd1 vccd1 vccd1 _17575_/C
+ sky130_fd_sc_hd__a211oi_4
X_14784_ _14670_/A _14669_/B _14667_/X vssd1 vssd1 vccd1 vccd1 _14784_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11996_ _11996_/A _11996_/B _11996_/C vssd1 vssd1 vccd1 vccd1 _12053_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12020__C _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19311_ _19311_/A _19311_/B vssd1 vssd1 vccd1 vccd1 _19313_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__19374__A1 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16523_ _16522_/B _16522_/C _16522_/A vssd1 vssd1 vccd1 vccd1 _16525_/B sky130_fd_sc_hd__a21o_1
X_13735_ _13734_/B _13734_/C _13734_/A vssd1 vssd1 vccd1 vccd1 _13735_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_156_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10947_ mstream_o[56] _10946_/Y _21568_/S vssd1 vssd1 vccd1 vccd1 _21593_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17385__B1 _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19242_ _19241_/B _19387_/B _19241_/A vssd1 vssd1 vccd1 vccd1 _19243_/C sky130_fd_sc_hd__a21o_1
X_16454_ _16451_/X _16454_/B vssd1 vssd1 vccd1 vccd1 _16749_/B sky130_fd_sc_hd__and2b_1
X_13666_ _16363_/A hold94/X _10852_/X fanout5/X _13665_/Y vssd1 vssd1 vccd1 vccd1
+ _13666_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_2_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10878_ _10878_/A _10885_/A vssd1 vssd1 vccd1 vccd1 _10878_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15405_ _15600_/B _15405_/B vssd1 vssd1 vccd1 vccd1 _15420_/A sky130_fd_sc_hd__and2_1
XFILLER_0_94_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_650 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13132__B _13573_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12674__D _14384_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19173_ _19163_/B _19169_/B _19161_/Y vssd1 vssd1 vccd1 vccd1 _19322_/A sky130_fd_sc_hd__a21oi_1
X_12617_ _12617_/A _12617_/B vssd1 vssd1 vccd1 vccd1 _12630_/A sky130_fd_sc_hd__xnor2_1
X_16385_ _16356_/A _16356_/B _16353_/X vssd1 vssd1 vccd1 vccd1 _16387_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_54_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13597_ _13597_/A _13752_/B vssd1 vssd1 vccd1 vccd1 _13600_/A sky130_fd_sc_hd__or2_1
XFILLER_0_155_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18124_ _18277_/A _18124_/B vssd1 vssd1 vccd1 vccd1 _18126_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_54_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15336_ _15336_/A _15430_/B _15336_/C vssd1 vssd1 vccd1 vccd1 _15338_/B sky130_fd_sc_hd__and3_2
XFILLER_0_54_776 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12548_ _12443_/A _12899_/B _12446_/B _12444_/X vssd1 vssd1 vccd1 vccd1 _12558_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18055_ _18055_/A _18055_/B vssd1 vssd1 vccd1 vccd1 _18057_/B sky130_fd_sc_hd__xnor2_2
X_15267_ _15267_/A _15400_/B _15268_/B vssd1 vssd1 vccd1 vccd1 _15464_/A sky130_fd_sc_hd__or3b_2
XFILLER_0_123_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_2 _10792_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14244__A _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19429__A2 _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12479_ _12479_/A _12479_/B _12479_/C _12479_/D vssd1 vssd1 vccd1 vccd1 _12479_/Y
+ sky130_fd_sc_hd__nor4_2
XFILLER_0_1_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17006_ _17005_/B _17005_/Y _16961_/Y _16963_/X vssd1 vssd1 vccd1 vccd1 _17006_/Y
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_50_960 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14218_ _15375_/A _14218_/B vssd1 vssd1 vccd1 vccd1 _14220_/C sky130_fd_sc_hd__and2_1
XFILLER_0_10_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11587__B _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16148__B1_N _15907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15198_ _15199_/A _15199_/B vssd1 vssd1 vccd1 vccd1 _15200_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_1_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14149_ _14149_/A _14149_/B _14149_/C vssd1 vssd1 vccd1 vccd1 _14149_/Y sky130_fd_sc_hd__nand3_1
Xfanout509 _16203_/D vssd1 vssd1 vccd1 vccd1 _16087_/A sky130_fd_sc_hd__buf_4
XFILLER_0_1_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18957_ _19587_/A _20242_/D _20249_/B _19445_/A vssd1 vssd1 vccd1 vccd1 _18957_/X
+ sky130_fd_sc_hd__a22o_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11488__A1 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17908_ _17908_/A _18026_/B _17908_/C vssd1 vssd1 vccd1 vccd1 _17910_/B sky130_fd_sc_hd__nand3_2
X_18888_ _19006_/B _18886_/X _18760_/Y _18763_/Y vssd1 vssd1 vccd1 vccd1 _18889_/C
+ sky130_fd_sc_hd__o211ai_2
XANTENNA__17612__A1 _17854_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17839_ _17708_/X _17837_/X _17838_/X _17831_/B vssd1 vssd1 vccd1 vccd1 _17839_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_117_1021 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20850_ _20724_/A _20855_/A _20723_/B _20720_/B _20720_/A vssd1 vssd1 vccd1 vccd1
+ _20852_/B sky130_fd_sc_hd__o32ai_4
XFILLER_0_7_1105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_1116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18168__A2 _18769_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_1065 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19509_ _20178_/D _20193_/D _19509_/C _19661_/A vssd1 vssd1 vccd1 vccd1 _19661_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__15522__B _15523_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20781_ _20916_/B _20781_/B vssd1 vssd1 vccd1 vccd1 _20783_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_18_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11542__S _11545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout157_A _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11660__A1 _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11660__B2 _13525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14138__B _14463_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17128__B1 _17146_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13401__A2 _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout324_A _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_979 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21402_ _15626_/Y _20514_/Y _21407_/S vssd1 vssd1 vccd1 vccd1 _21402_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_17_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12881__B _13157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_804 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21333_ hold156/X _21421_/S _21331_/Y _21332_/Y vssd1 vssd1 vccd1 vccd1 _21918_/D
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21264_ _21264_/A _21264_/B vssd1 vssd1 vccd1 vccd1 _21265_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19664__B _19664_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12912__A1 _14087_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20215_ _20215_/A _20215_/B vssd1 vssd1 vccd1 vccd1 _20218_/A sky130_fd_sc_hd__xor2_1
XANTENNA__12912__B2 _14089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21195_ _21196_/B _21195_/B vssd1 vssd1 vccd1 vccd1 _21197_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_25_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20146_ _20689_/A _20146_/B _21305_/A _21153_/B vssd1 vssd1 vccd1 vccd1 _20281_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__11479__A1 _18319_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20077_ _20078_/A _20078_/B vssd1 vssd1 vccd1 vccd1 _20079_/A sky130_fd_sc_hd__or2_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12402__A _12402_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18800__B1 _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _12223_/A _12528_/B vssd1 vssd1 vccd1 vccd1 _11853_/A sky130_fd_sc_hd__nand2_1
XANTENNA__12428__B1 _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15090__A1 _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15090__B2 _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10801_ sstream_o sstream_i[114] vssd1 vssd1 vccd1 vccd1 _21721_/D sky130_fd_sc_hd__and2_2
XFILLER_0_131_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15432__B _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11100__A0 _11066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18446__D _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11781_ _11781_/A _11781_/B _11781_/C vssd1 vssd1 vccd1 vccd1 _11813_/A sky130_fd_sc_hd__nand3_1
X_20979_ _20979_/A _21091_/B vssd1 vssd1 vccd1 vccd1 _20981_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_36_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11452__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_1164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13520_ _13520_/A _13520_/B vssd1 vssd1 vccd1 vccd1 _13520_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_83_816 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_827 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19108__A1 _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19108__B2 _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13451_ _13451_/A _13451_/B _13451_/C vssd1 vssd1 vccd1 vccd1 _13451_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_94_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18462__C _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12402_ _12402_/A _12402_/B vssd1 vssd1 vccd1 vccd1 _12406_/A sky130_fd_sc_hd__nand2_1
X_16170_ _16322_/B _16170_/B vssd1 vssd1 vccd1 vccd1 _16185_/A sky130_fd_sc_hd__and2_1
X_13382_ _13382_/A _13527_/B vssd1 vssd1 vccd1 vccd1 _13384_/B sky130_fd_sc_hd__or2_1
XFILLER_0_63_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15121_ _15024_/A _15024_/C _15024_/B vssd1 vssd1 vccd1 vccd1 _15122_/C sky130_fd_sc_hd__a21bo_1
XANTENNA__11688__A _14621_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12333_ _12334_/A _12334_/B vssd1 vssd1 vccd1 vccd1 _12333_/X sky130_fd_sc_hd__and2_1
XFILLER_0_69_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13156__A1 _13155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15052_ _15050_/X _15052_/B vssd1 vssd1 vccd1 vccd1 _15055_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_105_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13156__B2 _13155_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12264_ _12264_/A _12264_/B _12264_/C vssd1 vssd1 vccd1 vccd1 _12267_/C sky130_fd_sc_hd__nand3_2
XANTENNA__19574__B _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14999__A _15373_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14003_ _14002_/B _14002_/C _14002_/A vssd1 vssd1 vccd1 vccd1 _14004_/C sky130_fd_sc_hd__a21o_1
X_11215_ hold180/X _11126_/Y _11214_/X vssd1 vssd1 vccd1 vccd1 _11215_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_120_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12195_ _12195_/A _12195_/B _12195_/C vssd1 vssd1 vccd1 vccd1 _12203_/A sky130_fd_sc_hd__and3_2
X_19860_ _19961_/A _20381_/A _19857_/Y _19858_/X vssd1 vssd1 vccd1 vccd1 _19863_/B
+ sky130_fd_sc_hd__or4bb_1
XFILLER_0_102_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18811_ _18810_/A _18810_/B _18810_/C vssd1 vssd1 vccd1 vccd1 _18813_/C sky130_fd_sc_hd__a21o_1
X_11146_ hold204/X fanout23/X _11145_/X vssd1 vssd1 vccd1 vccd1 _11146_/X sky130_fd_sc_hd__a21o_1
X_19791_ _19792_/B _20081_/A vssd1 vssd1 vccd1 vccd1 _19796_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__13408__A _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19590__A _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15954_ _16084_/A _16203_/D _16084_/C _15954_/D vssd1 vssd1 vccd1 vccd1 _16089_/A
+ sky130_fd_sc_hd__and4_1
X_11077_ _10919_/X hold14/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21672_/D sky130_fd_sc_hd__mux2_1
X_18742_ _18584_/X _18587_/B _18739_/X _18741_/Y vssd1 vssd1 vccd1 vccd1 _18742_/X
+ sky130_fd_sc_hd__o211a_1
XANTENNA__12312__A _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14905_ _14906_/A _14906_/B vssd1 vssd1 vccd1 vccd1 _15067_/B sky130_fd_sc_hd__nand2_1
X_18673_ _18674_/A _18674_/B _18674_/C _18674_/D vssd1 vssd1 vccd1 vccd1 _18673_/Y
+ sky130_fd_sc_hd__nor4_1
XANTENNA__12669__D _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15885_ _15749_/A _15751_/X _16011_/B _15883_/X vssd1 vssd1 vccd1 vccd1 _16016_/C
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14836_ _14836_/A _14836_/B _14836_/C vssd1 vssd1 vccd1 vccd1 _14840_/B sky130_fd_sc_hd__nand3_2
X_17624_ _17737_/B _17622_/X _17522_/C _17524_/A vssd1 vssd1 vccd1 vccd1 _17625_/B
+ sky130_fd_sc_hd__o211ai_1
XFILLER_0_53_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_1205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17555_ _17555_/A _17555_/B vssd1 vssd1 vccd1 vccd1 _17564_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_129_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14767_ _15155_/C _15829_/C _15954_/D _15159_/D vssd1 vssd1 vccd1 vccd1 _14769_/A
+ sky130_fd_sc_hd__a22o_1
X_11979_ _11979_/A _11979_/B vssd1 vssd1 vccd1 vccd1 _11980_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_1249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11362__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18934__A _20088_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16506_ _16715_/A _16715_/B _16715_/C vssd1 vssd1 vccd1 vccd1 _16721_/A sky130_fd_sc_hd__a21oi_2
X_13718_ _13718_/A _13718_/B vssd1 vssd1 vccd1 vccd1 _13719_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11642__A1 _12426_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15908__A1 _15907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17486_ hold90/X _17485_/X fanout3/X vssd1 vssd1 vccd1 vccd1 hold91/A sky130_fd_sc_hd__mux2_1
X_14698_ _14698_/A _15514_/B _16266_/C _14698_/D vssd1 vssd1 vccd1 vccd1 _14702_/D
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_128_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_1171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_1248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11642__B2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16437_ _16437_/A _16437_/B vssd1 vssd1 vccd1 vccd1 _16437_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_27_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19225_ _19379_/B _19227_/C _19227_/D _19382_/A vssd1 vssd1 vccd1 vccd1 _19230_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13649_ _13648_/A _13648_/B _13648_/C _13648_/D vssd1 vssd1 vccd1 vccd1 _13649_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_156_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19156_ _19157_/A _19157_/B vssd1 vssd1 vccd1 vccd1 _19320_/A sky130_fd_sc_hd__nor2_1
X_16368_ _16349_/A _16368_/B vssd1 vssd1 vccd1 vccd1 _16370_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_2_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_1100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16173__B _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18107_ _18107_/A _18107_/B vssd1 vssd1 vccd1 vccd1 _18126_/A sky130_fd_sc_hd__or2_2
X_15319_ _16092_/D _15961_/D _15717_/C _15976_/D vssd1 vssd1 vccd1 vccd1 _15450_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19087_ _20101_/A _19087_/B _19705_/B _19703_/C vssd1 vssd1 vccd1 vccd1 _19088_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_152_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16299_ _16300_/A _16300_/B vssd1 vssd1 vccd1 vccd1 _16301_/A sky130_fd_sc_hd__and2_1
XFILLER_0_124_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18038_ _18175_/B _18038_/B _18038_/C vssd1 vssd1 vccd1 vccd1 _18164_/A sky130_fd_sc_hd__nand3_1
XANTENNA__16884__A2 _17019_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14702__A _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20968__A1 _20838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19822__A2 _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout306 _19337_/D vssd1 vssd1 vccd1 vccd1 _18849_/B sky130_fd_sc_hd__buf_4
X_20000_ _20000_/A _20000_/B vssd1 vssd1 vccd1 vccd1 _20014_/A sky130_fd_sc_hd__xor2_1
Xfanout317 _21792_/Q vssd1 vssd1 vccd1 vccd1 _17854_/B sky130_fd_sc_hd__buf_4
Xfanout328 _21788_/Q vssd1 vssd1 vccd1 vccd1 _16406_/B sky130_fd_sc_hd__clkbuf_8
Xfanout339 _21784_/Q vssd1 vssd1 vccd1 vccd1 _15174_/D sky130_fd_sc_hd__clkbuf_4
X_19989_ fanout96/X _19988_/X _19987_/X vssd1 vssd1 vccd1 vccd1 _19991_/A sky130_fd_sc_hd__a21bo_1
XFILLER_0_94_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15236__C _15375_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21951_ _21963_/CLK _21951_/D vssd1 vssd1 vccd1 vccd1 hold224/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__17597__B1 _17595_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout274_A _21800_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19650__D _19650_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20902_ _20902_/A _20902_/B vssd1 vssd1 vccd1 vccd1 _20904_/C sky130_fd_sc_hd__or2_1
XFILLER_0_55_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21882_ _21949_/CLK _21882_/D vssd1 vssd1 vccd1 vccd1 hold76/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_94_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12876__B _13012_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20833_ _20830_/Y _20831_/X _20667_/B _20710_/A vssd1 vssd1 vccd1 vccd1 _20834_/B
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_49_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout441_A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11272__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19889__A2 _21278_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11633__A1 _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11633__B2 _12750_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20764_ _20896_/A _20762_/X _20596_/Y _20601_/A vssd1 vssd1 vccd1 vccd1 _20764_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20695_ _20696_/A _20696_/B vssd1 vssd1 vccd1 vccd1 _20823_/B sky130_fd_sc_hd__nand2_1
XANTENNA__19378__C _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__20317__C _20721_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17521__B1 _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_1228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21316_ _21316_/A _21316_/B vssd1 vssd1 vccd1 vccd1 _21317_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_131_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_993 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21247_ _21253_/B _21247_/B vssd1 vssd1 vccd1 vccd1 _21248_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_7_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20333__B _20975_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11000_ mstream_o[74] hold81/X _11005_/S vssd1 vssd1 vccd1 vccd1 _21611_/D sky130_fd_sc_hd__mux2_1
X_21178_ _21178_/A _21178_/B vssd1 vssd1 vccd1 vccd1 _21179_/B sky130_fd_sc_hd__and2_1
XANTENNA__11955__B _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_1153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20129_ _20838_/B _20671_/B _20130_/C _20330_/A vssd1 vssd1 vccd1 vccd1 _20131_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13310__A1 _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13310__B2 _15076_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18738__B _19051_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17642__B _18030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12951_ _12951_/A _12951_/B vssd1 vssd1 vccd1 vccd1 _12952_/B sky130_fd_sc_hd__nor2_2
XTAP_3211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_1204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11902_ _11836_/A _11836_/C _11836_/B vssd1 vssd1 vccd1 vccd1 _11902_/X sky130_fd_sc_hd__a21o_1
X_15670_ _15670_/A _15670_/B vssd1 vssd1 vccd1 vccd1 _15678_/A sky130_fd_sc_hd__nand2_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_200 hold268/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12882_ _13157_/A _14024_/B _13155_/C _13155_/D vssd1 vssd1 vccd1 vccd1 _12884_/B
+ sky130_fd_sc_hd__nand4_2
XTAP_3266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_211 hold275/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_222 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14621_ _14463_/D _15838_/B _16314_/D _14621_/D vssd1 vssd1 vccd1 vccd1 _14624_/A
+ sky130_fd_sc_hd__and4b_2
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_233 hold299/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ _11833_/A _11833_/B _11833_/C vssd1 vssd1 vccd1 vccd1 _11834_/B sky130_fd_sc_hd__and3_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_244 _11347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_255 v2z[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_266 hold286/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_974 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_277 hold283/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18001__A1 _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17340_ _17340_/A _17340_/B _17340_/C vssd1 vssd1 vccd1 vccd1 _17343_/A sky130_fd_sc_hd__nand3_1
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14552_ _14551_/B _14551_/C _14551_/A vssd1 vssd1 vccd1 vccd1 _14553_/B sky130_fd_sc_hd__a21oi_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_288 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11764_ _11764_/A _11764_/B _11764_/C vssd1 vssd1 vccd1 vccd1 _11791_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_55_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_299 hold306/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13503_ _13353_/B _13353_/Y _13500_/X _13502_/Y vssd1 vssd1 vccd1 vccd1 _13503_/Y
+ sky130_fd_sc_hd__a211oi_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13898__A _15514_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17271_ _17381_/A _17381_/B vssd1 vssd1 vccd1 vccd1 _21334_/B sky130_fd_sc_hd__xnor2_4
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14483_ _14482_/B _14482_/C _14482_/A vssd1 vssd1 vccd1 vccd1 _14484_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_128_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13113__D _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11695_ _12426_/B _12619_/A _12330_/A _11694_/D vssd1 vssd1 vccd1 vccd1 _11697_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__21629__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19010_ _19194_/A _19010_/B vssd1 vssd1 vccd1 vccd1 _19011_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_153_534 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_16222_ _16223_/A _16223_/B vssd1 vssd1 vccd1 vccd1 _16337_/B sky130_fd_sc_hd__nand2_1
XANTENNA__13377__A1 _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13377__B2 _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13434_ _13430_/X _13431_/Y _13280_/A _13280_/Y vssd1 vssd1 vccd1 vccd1 _13496_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_82_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16153_ _16414_/A _16268_/B _16266_/C _16391_/A vssd1 vssd1 vccd1 vccd1 _16157_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13365_ _13365_/A _13365_/B vssd1 vssd1 vccd1 vccd1 _13365_/X sky130_fd_sc_hd__or2_1
XFILLER_0_140_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13129__A1 _13867_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15104_ _15226_/B _15103_/C _15103_/A vssd1 vssd1 vccd1 vccd1 _15104_/Y sky130_fd_sc_hd__a21oi_2
XANTENNA__13129__B2 _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12316_ _12316_/A _12316_/B vssd1 vssd1 vccd1 vccd1 _12317_/B sky130_fd_sc_hd__or2_1
X_16084_ _16084_/A _16196_/A _16084_/C _16084_/D vssd1 vssd1 vccd1 vccd1 _16201_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_121_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13296_ _14195_/A _15763_/A _13293_/Y _13445_/A vssd1 vssd1 vccd1 vccd1 _13297_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_146_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14877__A1 _21769_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11568__D _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15035_ _15035_/A _15035_/B _15127_/B vssd1 vssd1 vccd1 vccd1 _15037_/B sky130_fd_sc_hd__nand3_1
X_19912_ _19911_/B _19911_/C _19911_/A vssd1 vssd1 vccd1 vccd1 _19914_/B sky130_fd_sc_hd__a21o_1
X_12247_ _12261_/A _12246_/C _12246_/D _12269_/B vssd1 vssd1 vccd1 vccd1 _12249_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12352__A2 _12780_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19843_ _19843_/A _19843_/B vssd1 vssd1 vccd1 vccd1 _19929_/A sky130_fd_sc_hd__xnor2_1
X_12178_ _12148_/A _12148_/C _12148_/B vssd1 vssd1 vccd1 vccd1 _12195_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_120_1242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18929__A _21833_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17833__A _20770_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ _12269_/D _11128_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21726_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19774_ _19621_/A _19621_/B _19619_/Y vssd1 vssd1 vccd1 vccd1 _19776_/B sky130_fd_sc_hd__a21oi_1
X_16986_ _16986_/A _16986_/B vssd1 vssd1 vccd1 vccd1 _16992_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__19751__C _19751_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21355__A _21720_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18725_ _18725_/A _18847_/A _18725_/C vssd1 vssd1 vccd1 vccd1 _18847_/B sky130_fd_sc_hd__nor3_1
X_15937_ _15938_/A _15938_/B vssd1 vssd1 vccd1 vccd1 _16069_/B sky130_fd_sc_hd__nand2_1
XANTENNA__11312__A0 _14176_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xwire16 wire16/A vssd1 vssd1 vccd1 vccd1 wire16/X sky130_fd_sc_hd__buf_4
X_15868_ _15867_/B _15867_/C _15867_/A vssd1 vssd1 vccd1 vccd1 _15868_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__22070__RESET_B fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18656_ _18656_/A _18656_/B _18656_/C vssd1 vssd1 vccd1 vccd1 _18658_/B sky130_fd_sc_hd__nand3_1
XANTENNA__11863__A1 _12109_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14819_ _16203_/D _15022_/B _14820_/C _14820_/D vssd1 vssd1 vccd1 vccd1 _14819_/X
+ sky130_fd_sc_hd__and4_1
X_17607_ _17607_/A _17715_/A vssd1 vssd1 vccd1 vccd1 _17617_/A sky130_fd_sc_hd__nor2_1
X_15799_ _15800_/A _15800_/B vssd1 vssd1 vccd1 vccd1 _15986_/B sky130_fd_sc_hd__or2_1
X_18587_ _18587_/A _18587_/B vssd1 vssd1 vccd1 vccd1 _18590_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_114_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_1108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11615__A1 _12302_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_1181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17538_ _17422_/X _17424_/X _17535_/X _17536_/Y vssd1 vssd1 vccd1 vccd1 _17538_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11615__B2 _13985_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17469_ _17466_/X _17467_/Y _17356_/C _17355_/Y vssd1 vssd1 vccd1 vccd1 _17469_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_74_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19208_ _19035_/B _19037_/B _19363_/A _19207_/Y vssd1 vssd1 vccd1 vccd1 _19363_/B
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20480_ _20481_/B _20481_/A vssd1 vssd1 vccd1 vccd1 _20480_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_6_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13320__B _14712_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19139_ _19139_/A _19139_/B _19139_/C vssd1 vssd1 vccd1 vccd1 _19139_/Y sky130_fd_sc_hd__nand3_2
XFILLER_0_131_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_921 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17503__B1 _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20102__A2 _21815_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_965 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21101_ _21296_/A _21311_/B _21102_/C _21102_/D vssd1 vssd1 vccd1 vccd1 _21103_/A
+ sky130_fd_sc_hd__a22oi_1
X_22081_ _22096_/CLK _22081_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[17] sky130_fd_sc_hd__dfrtp_4
XANTENNA__19256__B1 _18640_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21032_ _20912_/A _20912_/B _20651_/B vssd1 vssd1 vccd1 vccd1 _21033_/B sky130_fd_sc_hd__o21ai_4
Xfanout103 _19691_/D vssd1 vssd1 vccd1 vccd1 _19227_/D sky130_fd_sc_hd__buf_4
Xfanout114 _21839_/Q vssd1 vssd1 vccd1 vccd1 _17741_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_22_1125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout125 _20689_/A vssd1 vssd1 vccd1 vccd1 _19906_/A sky130_fd_sc_hd__buf_8
XANTENNA_fanout391_A _21771_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout136 _20774_/A vssd1 vssd1 vccd1 vccd1 _17300_/C sky130_fd_sc_hd__buf_4
XANTENNA_fanout489_A _21747_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout147 _19092_/B vssd1 vssd1 vccd1 vccd1 _18622_/B sky130_fd_sc_hd__clkbuf_8
XANTENNA__13048__A _14572_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout158 _21830_/Q vssd1 vssd1 vccd1 vccd1 _20088_/A sky130_fd_sc_hd__buf_6
Xfanout169 _19732_/A vssd1 vssd1 vccd1 vccd1 _18787_/A sky130_fd_sc_hd__buf_4
XFILLER_0_96_1259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11303__B1 _11302_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20169__A2 _20838_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16359__A _16359_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21934_ _21934_/CLK _21934_/D vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__17181__C _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_941 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_21865_ _21948_/CLK _21865_/D vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__16509__D _16860_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20816_ _20817_/B _20817_/A vssd1 vssd1 vccd1 vccd1 _20951_/A sky130_fd_sc_hd__nand2b_1
XANTENNA_hold234_A hold234/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21796_ _21803_/CLK _21796_/D vssd1 vssd1 vccd1 vccd1 _21796_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19731__A1 _19732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19731__B2 _19732_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20747_ _20747_/A _20747_/B _20747_/C vssd1 vssd1 vccd1 vccd1 _20835_/B sky130_fd_sc_hd__or3_1
XANTENNA__21722__RESET_B fanout644/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14556__B1 _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11480_ _11498_/A1 t1y[10] t0x[10] _11501_/B2 vssd1 vssd1 vccd1 vccd1 _11480_/X sky130_fd_sc_hd__a22o_1
X_20678_ _20678_/A _20801_/B vssd1 vssd1 vccd1 vccd1 _20681_/A sky130_fd_sc_hd__or2_1
XFILLER_0_33_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14326__B _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19495__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13150_ _13864_/B _14537_/A vssd1 vssd1 vccd1 vccd1 _13154_/A sky130_fd_sc_hd__and2_1
XFILLER_0_115_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_1025 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_1074 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17637__B _18008_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12101_ _12100_/B _12100_/C _12100_/A vssd1 vssd1 vccd1 vccd1 _12102_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_20_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13081_ _13077_/X _13078_/Y _12938_/B _12938_/Y vssd1 vssd1 vccd1 vccd1 _13083_/C
+ sky130_fd_sc_hd__o211a_1
XANTENNA__14323__A3 _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12032_ _12286_/B _12286_/C _12286_/A vssd1 vssd1 vccd1 vccd1 _12294_/C sky130_fd_sc_hd__o21a_1
Xhold190 hold190/A vssd1 vssd1 vccd1 vccd1 hold190/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19852__B _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18749__A _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11177__S _11195_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16840_ _16840_/A _16840_/B _16840_/C vssd1 vssd1 vccd1 vccd1 _16840_/X sky130_fd_sc_hd__and3_1
XANTENNA__17273__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19571__C _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16481__B1 _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16771_ _16771_/A _16771_/B vssd1 vssd1 vccd1 vccd1 _16773_/C sky130_fd_sc_hd__xnor2_1
X_13983_ _14133_/D _13983_/B _16404_/B _16406_/B vssd1 vssd1 vccd1 vccd1 _13985_/D
+ sky130_fd_sc_hd__and4_2
X_15722_ _15722_/A _15722_/B vssd1 vssd1 vccd1 vccd1 _15724_/B sky130_fd_sc_hd__xnor2_1
X_18510_ _18511_/A _18511_/B _18511_/C vssd1 vssd1 vccd1 vccd1 _18510_/X sky130_fd_sc_hd__and3_1
XFILLER_0_38_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_3030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12934_ _12971_/B _12934_/B _12934_/C _12934_/D vssd1 vssd1 vccd1 vccd1 _12934_/X
+ sky130_fd_sc_hd__and4_2
XFILLER_0_137_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_3041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_19490_ _19490_/A _19490_/B vssd1 vssd1 vccd1 vccd1 _19492_/A sky130_fd_sc_hd__xnor2_4
XTAP_3052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__16233__B1 _16232_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15653_ _16305_/B _16399_/A _15653_/C _15911_/C vssd1 vssd1 vccd1 vccd1 _15849_/A
+ sky130_fd_sc_hd__nand4_2
XTAP_3074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18441_ _18564_/B _18441_/B vssd1 vssd1 vccd1 vccd1 _18441_/X sky130_fd_sc_hd__and2_1
XTAP_3085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12865_ _12865_/A _12865_/B vssd1 vssd1 vccd1 vccd1 _12868_/C sky130_fd_sc_hd__xnor2_2
XTAP_3096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18484__A _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14604_ _14608_/B _14604_/B vssd1 vssd1 vccd1 vccd1 _14605_/B sky130_fd_sc_hd__or2_4
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15901__A _16031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18372_ _18373_/A _18373_/B _18373_/C _18373_/D vssd1 vssd1 vccd1 vccd1 _18372_/Y
+ sky130_fd_sc_hd__nor4_1
X_11816_ _11816_/A _11816_/B _11816_/C vssd1 vssd1 vccd1 vccd1 _11857_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_68_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15584_ _15585_/A _15585_/B vssd1 vssd1 vccd1 vccd1 _15584_/Y sky130_fd_sc_hd__nand2_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12796_ _12795_/A _12795_/B _12795_/C vssd1 vssd1 vccd1 vccd1 _12798_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_28_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17323_ _17417_/A _19432_/A vssd1 vssd1 vccd1 vccd1 _17327_/A sky130_fd_sc_hd__nand2_1
XANTENNA__19722__A1 _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14535_ _14993_/A _15892_/B _16328_/A vssd1 vssd1 vccd1 vccd1 _14535_/X sky130_fd_sc_hd__and3_1
XFILLER_0_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11747_ _11747_/A _11747_/B vssd1 vssd1 vccd1 vccd1 _11748_/C sky130_fd_sc_hd__nor2_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17254_ _17250_/X _17252_/Y _16634_/B _16634_/Y vssd1 vssd1 vccd1 vccd1 _17256_/D
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14466_ _14466_/A _14466_/B vssd1 vssd1 vccd1 vccd1 _14467_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_3_1185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11678_ _12229_/A _12642_/A _12637_/A _12155_/B vssd1 vssd1 vccd1 vccd1 _11680_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13778__D _15234_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14236__B _15093_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16205_ _16321_/A _16205_/B vssd1 vssd1 vccd1 vccd1 _16206_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_141_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13417_ _14027_/A _14516_/A _14365_/C _13864_/B vssd1 vssd1 vccd1 vccd1 _13417_/Y
+ sky130_fd_sc_hd__a22oi_1
XANTENNA__16154__D _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17185_ _17186_/B _17185_/B vssd1 vssd1 vccd1 vccd1 _17187_/B sky130_fd_sc_hd__and2b_1
XANTENNA__19486__B1 _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14397_ _14398_/A _14532_/B _14398_/C vssd1 vssd1 vccd1 vccd1 _14397_/X sky130_fd_sc_hd__and3_1
XFILLER_0_52_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16732__A _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_1084 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__19746__C _19868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16136_ _16133_/Y _16134_/X _16001_/X _16003_/Y vssd1 vssd1 vccd1 vccd1 _16136_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_141_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_1114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13348_ _13348_/A _13348_/B _13348_/C vssd1 vssd1 vccd1 vccd1 _13348_/X sky130_fd_sc_hd__or3_2
XFILLER_0_84_1174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_1027 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16451__B _17029_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16067_ _16067_/A _16067_/B vssd1 vssd1 vccd1 vccd1 _16069_/C sky130_fd_sc_hd__xnor2_1
X_13279_ _13427_/B _13278_/B _13278_/C vssd1 vssd1 vccd1 vccd1 _13280_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_59_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_957 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15018_ _15961_/D _15788_/B vssd1 vssd1 vccd1 vccd1 _15019_/B sky130_fd_sc_hd__and2_1
XANTENNA__11087__S _11087_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18461__A1 _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19826_ _19826_/A _19826_/B _20043_/B vssd1 vssd1 vccd1 vccd1 _19828_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_120_1061 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18461__B2 _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17282__B _17741_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19757_ _19756_/B _19756_/C _19756_/A vssd1 vssd1 vccd1 vccd1 _19758_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_155_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16969_ _17145_/A _17013_/D vssd1 vssd1 vccd1 vccd1 _16971_/B sky130_fd_sc_hd__and2_1
XANTENNA__13018__D _21768_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18708_ _18708_/A _18708_/B vssd1 vssd1 vccd1 vccd1 _18725_/A sky130_fd_sc_hd__or2_1
XFILLER_0_155_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15514__C _16173_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19688_ _19823_/A _20671_/B vssd1 vssd1 vccd1 vccd1 _19689_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18639_ _18789_/A _18640_/B _18640_/C _18784_/A vssd1 vssd1 vccd1 vccd1 _18641_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17972__B1 _17970_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21650_ _21722_/CLK hold284/X fanout643/X vssd1 vssd1 vccd1 vccd1 mstream_o[113]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__13034__C _15076_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_315 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20859__B1 _21305_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20601_ _20601_/A _20601_/B vssd1 vssd1 vccd1 vccd1 _20621_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_117_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19002__B _21373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21581_ _22106_/CLK _21581_/D _11089_/A vssd1 vssd1 vccd1 vccd1 mstream_o[44] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_89_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20532_ _20533_/A _20533_/B vssd1 vssd1 vccd1 vccd1 _20532_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_145_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20463_ _20462_/D _21293_/B _21261_/B _18008_/A vssd1 vssd1 vccd1 vccd1 _20464_/B
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__19477__B1 _14605_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout404_A _13155_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13761__A1 _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13985__B _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20394_ _21831_/Q _20394_/B _21056_/B vssd1 vssd1 vccd1 vccd1 _20650_/B sky130_fd_sc_hd__and3_1
XFILLER_0_15_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21036__B1 _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_22064_ _22069_/CLK _22064_/D fanout639/X vssd1 vssd1 vccd1 vccd1 mstream_o[0] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_100_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14312__D _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21015_ _21016_/A _21016_/B _21016_/C vssd1 vssd1 vccd1 vccd1 _21129_/A sky130_fd_sc_hd__o21a_1
XANTENNA__20477__A1_N _20583_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1045 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17192__B _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10980_ hold92/A hold171/A vssd1 vssd1 vccd1 vccd1 _10982_/A sky130_fd_sc_hd__or2_1
XANTENNA__19952__A1 _19951_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21917_ _21948_/CLK _21917_/D vssd1 vssd1 vccd1 vccd1 hold121/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__13225__B _21355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16766__A1 _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16766__B2 _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12650_ _12651_/A _12651_/B vssd1 vssd1 vccd1 vccd1 _12650_/X sky130_fd_sc_hd__and2_2
X_21848_ _21853_/CLK _21848_/D vssd1 vssd1 vccd1 vccd1 _21848_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_0_139_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14241__A2 _14557_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19704__A1 _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11601_ _11602_/A _11602_/B vssd1 vssd1 vccd1 vccd1 _11601_/X sky130_fd_sc_hd__and2_1
XFILLER_0_155_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12581_ _12577_/X _12579_/Y _12471_/B _12471_/Y vssd1 vssd1 vccd1 vccd1 _12583_/D
+ sky130_fd_sc_hd__o211a_1
X_21779_ _21789_/CLK _21779_/D vssd1 vssd1 vccd1 vccd1 hold333/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_148_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14320_ _14321_/B vssd1 vssd1 vccd1 vccd1 _14320_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_1103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11532_ _11544_/A1 t2x[27] v1z[27] fanout21/X _11531_/X vssd1 vssd1 vccd1 vccd1 _11532_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_1274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18751__B _19240_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14251_ _14251_/A _14251_/B _14251_/C vssd1 vssd1 vccd1 vccd1 _14418_/A sky130_fd_sc_hd__and3_4
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11463_ _21718_/D t2x[4] v1z[4] fanout17/X _11462_/X vssd1 vssd1 vccd1 vccd1 _11463_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13202_ _13198_/X _13200_/Y _13062_/B _13062_/Y vssd1 vssd1 vccd1 vccd1 _13204_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14182_ _14508_/A _14813_/A _14817_/C _14817_/D vssd1 vssd1 vccd1 vccd1 _14185_/D
+ sky130_fd_sc_hd__nand4_1
XANTENNA__13895__B _14537_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11394_ hold292/X fanout28/X _11393_/X vssd1 vssd1 vccd1 vccd1 _11394_/X sky130_fd_sc_hd__a21o_1
XANTENNA__16271__B _16371_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13133_ _13858_/B _13573_/D _13267_/A _13132_/D vssd1 vssd1 vccd1 vccd1 _13134_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__17494__A2 _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18990_ _18987_/X _18988_/X _18826_/C _18826_/Y vssd1 vssd1 vccd1 vccd1 _18991_/C
+ sky130_fd_sc_hd__a211oi_1
XANTENNA__17086__C _17086_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ _12924_/B _12924_/Y _13061_/X _13063_/Y vssd1 vssd1 vccd1 vccd1 _13067_/B
+ sky130_fd_sc_hd__a211oi_4
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17941_ _17940_/A _17940_/B _17940_/C vssd1 vssd1 vccd1 vccd1 _17943_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_40_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21578__A1 _11063_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12015_ _12015_/A _12015_/B vssd1 vssd1 vccd1 vccd1 _12017_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__18443__A1 _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17872_ _18008_/B _18010_/A _19906_/A _20146_/B vssd1 vssd1 vccd1 vccd1 _18006_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__18443__B2 _19373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13119__C _21776_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19611_ _19612_/A _19612_/B vssd1 vssd1 vccd1 vccd1 _19611_/Y sky130_fd_sc_hd__nor2_1
X_16823_ _16823_/A _16823_/B _16823_/C vssd1 vssd1 vccd1 vccd1 _16823_/X sky130_fd_sc_hd__and3_1
XFILLER_0_75_1118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19542_ _19542_/A _19542_/B vssd1 vssd1 vccd1 vccd1 _19556_/A sky130_fd_sc_hd__xnor2_1
X_13966_ _13966_/A _13966_/B vssd1 vssd1 vccd1 vccd1 _13967_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16754_ _16754_/A _16754_/B _16754_/C vssd1 vssd1 vccd1 vccd1 _16754_/Y sky130_fd_sc_hd__nand3_4
XFILLER_0_88_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18746__A2 _19529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15705_ _15705_/A _15705_/B vssd1 vssd1 vccd1 vccd1 _15706_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12917_ _12916_/A _12916_/B _12916_/C vssd1 vssd1 vccd1 vccd1 _12918_/C sky130_fd_sc_hd__a21o_1
X_16685_ _16657_/X _16658_/Y _16682_/A _16681_/Y vssd1 vssd1 vccd1 vccd1 _16686_/C
+ sky130_fd_sc_hd__a211o_1
X_19473_ _19161_/Y _19319_/X _19321_/B vssd1 vssd1 vccd1 vccd1 _19475_/A sky130_fd_sc_hd__o21ai_2
X_13897_ _15514_/B _14212_/D _14218_/B _15514_/A vssd1 vssd1 vccd1 vccd1 _13901_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18424_ _18269_/Y _18272_/X _18542_/A _18423_/X vssd1 vssd1 vccd1 vccd1 _18542_/B
+ sky130_fd_sc_hd__a211oi_2
X_15636_ _15640_/A _15803_/B vssd1 vssd1 vccd1 vccd1 _15641_/A sky130_fd_sc_hd__or2_2
XANTENNA__21352__B _21352_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ _12984_/A _12848_/B _13682_/C _14018_/C vssd1 vssd1 vccd1 vccd1 _12984_/B
+ sky130_fd_sc_hd__and4b_1
XFILLER_0_5_1225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14232__A2 _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_944 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20249__A _20249_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15567_ _15567_/A _15567_/B _15567_/C vssd1 vssd1 vccd1 vccd1 _15567_/X sky130_fd_sc_hd__or3_4
XFILLER_0_5_1269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_18355_ _18355_/A _18355_/B _18355_/C vssd1 vssd1 vccd1 vccd1 _18357_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_139_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12779_ _12780_/B _13034_/D _14386_/B _12780_/A vssd1 vssd1 vccd1 vccd1 _12779_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_29_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__14247__A _14248_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19171__A2 _19169_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_999 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14518_ _21743_/Q _15808_/C _14518_/C _14671_/A vssd1 vssd1 vccd1 vccd1 _14671_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_86_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17306_ _17520_/B _20249_/A vssd1 vssd1 vccd1 vccd1 _17310_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15498_ _21720_/Q hold95/X _10941_/X fanout5/X vssd1 vssd1 vccd1 vccd1 _15498_/X
+ sky130_fd_sc_hd__a22o_1
X_18286_ _18286_/A _18286_/B vssd1 vssd1 vccd1 vccd1 _18287_/B sky130_fd_sc_hd__nand2_1
XANTENNA__17182__A1 _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_662 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__17182__B2 _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_14449_ fanout9/X _14449_/B vssd1 vssd1 vccd1 vccd1 _14449_/Y sky130_fd_sc_hd__nor2_1
X_17237_ _17657_/A _19445_/A vssd1 vssd1 vccd1 vccd1 _17240_/A sky130_fd_sc_hd__and2_1
XFILLER_0_43_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_17168_ _17168_/A _17168_/B _17168_/C vssd1 vssd1 vccd1 vccd1 _17169_/C sky130_fd_sc_hd__or3_1
XFILLER_0_4_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17277__B _17387_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16119_ _16119_/A _16119_/B _16119_/C vssd1 vssd1 vccd1 vccd1 _16120_/A sky130_fd_sc_hd__or3_2
XANTENNA__17485__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_17099_ _17099_/A _17099_/B _17099_/C vssd1 vssd1 vccd1 vccd1 _17134_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_12_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_110_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21569__A1 _11043_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_985 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__15806__A _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20431__B _21169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20241__A1 _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20241__B2 _20774_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19809_ _19809_/A _19809_/B vssd1 vssd1 vccd1 vccd1 _19814_/A sky130_fd_sc_hd__or2_1
XANTENNA__13259__B1 _13258_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17443__D _17443_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11545__S _11545_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout187_A _21824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18198__B1 _19868_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16748__A1 _17096_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout354_A _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16637__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_1241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21702_ _22096_/CLK _21702_/D vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfxtp_1
XANTENNA__19013__A _19493_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_922 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_933 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_1079 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21633_ _21682_/CLK _21633_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[96] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_47_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout521_A _13877_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14157__A _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18257__A1_N _18857_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11280__S _11352_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout619_A _21717_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13982__A1 _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13982__B2 _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21564_ mstream_o[27] hold45/X _21579_/S vssd1 vssd1 vccd1 vccd1 _22091_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_74_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_20515_ hold185/X fanout7/X _15626_/Y _11550_/B vssd1 vssd1 vccd1 vccd1 _20515_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21495_ hold298/X sstream_i[72] _21507_/S vssd1 vssd1 vccd1 vccd1 _22022_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_31_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20606__B _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20446_ _20446_/A _20446_/B vssd1 vssd1 vccd1 vccd1 _20449_/C sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20377_ _20770_/B _20377_/B vssd1 vssd1 vccd1 vccd1 _20377_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_63_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__22102__RESET_B _11089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17915__B _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_1229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22047_ _22049_/CLK _22047_/D vssd1 vssd1 vccd1 vccd1 hold258/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__15435__B _15698_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21156__C _21256_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11455__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13820_ _14312_/D _16399_/B _16409_/B _14133_/D vssd1 vssd1 vccd1 vccd1 _13824_/D
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15161__A2_N _15838_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13751_ _13751_/A _13751_/B vssd1 vssd1 vccd1 vccd1 _13754_/A sky130_fd_sc_hd__nand2_1
X_10963_ _10961_/X _10967_/C vssd1 vssd1 vccd1 vccd1 _10965_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13670__B1 _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12702_ _12701_/B _12701_/C _12701_/A vssd1 vssd1 vccd1 vccd1 _12702_/X sky130_fd_sc_hd__a21o_1
X_16470_ _17300_/C _17520_/D _17124_/C _17282_/A vssd1 vssd1 vccd1 vccd1 _16471_/A
+ sky130_fd_sc_hd__and4_1
X_13682_ _13679_/Y _13835_/A _13682_/C _16328_/B vssd1 vssd1 vccd1 vccd1 _13835_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_85_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10894_ hold83/A hold137/A vssd1 vssd1 vccd1 vccd1 _10897_/A sky130_fd_sc_hd__or2_1
XANTENNA__16266__B _16414_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15421_ _15420_/B _15420_/C _15420_/A vssd1 vssd1 vccd1 vccd1 _15421_/X sky130_fd_sc_hd__a21o_1
X_12633_ _12543_/X _12546_/Y _12631_/A _12632_/Y vssd1 vssd1 vccd1 vccd1 _12716_/A
+ sky130_fd_sc_hd__a211o_2
XFILLER_0_156_949 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19477__A2_N fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15352_ _15354_/A _15354_/B vssd1 vssd1 vccd1 vccd1 _15352_/Y sky130_fd_sc_hd__nand2b_1
X_18140_ _18288_/B _18140_/B _18140_/C vssd1 vssd1 vccd1 vccd1 _18142_/A sky130_fd_sc_hd__and3_1
XFILLER_0_109_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12564_ _12784_/A _13034_/D vssd1 vssd1 vccd1 vccd1 _12567_/A sky130_fd_sc_hd__and2_1
XANTENNA__13402__C _13858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1060 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14303_ _14303_/A _14303_/B vssd1 vssd1 vccd1 vccd1 _14345_/A sky130_fd_sc_hd__nor2_2
XFILLER_0_81_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11515_ _11514_/X _18732_/C _11521_/S vssd1 vssd1 vccd1 vccd1 _21843_/D sky130_fd_sc_hd__mux2_1
X_18071_ _18071_/A _18071_/B _18071_/C vssd1 vssd1 vccd1 vccd1 _18074_/A sky130_fd_sc_hd__nand3_2
X_15283_ _15284_/A _15284_/B vssd1 vssd1 vccd1 vccd1 _15283_/Y sky130_fd_sc_hd__nand2b_1
XANTENNA__14217__D _14217_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17378__A _21142_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12495_ hold113/X _12494_/X fanout3/X vssd1 vssd1 vccd1 vccd1 hold114/A sky130_fd_sc_hd__mux2_1
X_17022_ _17096_/A _17145_/B vssd1 vssd1 vccd1 vccd1 _17023_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_1177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14234_ _14557_/A _14557_/B _14234_/C _15001_/B vssd1 vssd1 vccd1 vccd1 _14403_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_0_1188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11446_ _11445_/X hold294/X _11446_/S vssd1 vssd1 vccd1 vccd1 _21820_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_145_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_1253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_14165_ _14162_/X _14163_/Y _14002_/B _14004_/B vssd1 vssd1 vccd1 vccd1 _14165_/Y
+ sky130_fd_sc_hd__o211ai_2
XFILLER_0_106_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11377_ _11376_/X _17619_/A _11401_/S vssd1 vssd1 vccd1 vccd1 _21797_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13116_ _14133_/D _13997_/C vssd1 vssd1 vccd1 vccd1 _13117_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_81_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14096_ _14095_/B _14095_/C _14095_/A vssd1 vssd1 vccd1 vccd1 _14098_/B sky130_fd_sc_hd__a21o_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18973_ _18972_/A _18972_/B _18972_/C vssd1 vssd1 vccd1 vccd1 _18975_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ _13047_/A _13047_/B vssd1 vssd1 vccd1 vccd1 _13056_/A sky130_fd_sc_hd__xnor2_2
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17924_ _18058_/A _17924_/B vssd1 vssd1 vccd1 vccd1 _17928_/A sky130_fd_sc_hd__nand2_1
X_17855_ _17980_/A vssd1 vssd1 vccd1 vccd1 _17857_/C sky130_fd_sc_hd__inv_2
XANTENNA__11365__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16806_ _16806_/A _16806_/B _16806_/C vssd1 vssd1 vccd1 vccd1 _16876_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_89_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17786_ _19439_/A _17915_/D vssd1 vssd1 vccd1 vccd1 _17790_/A sky130_fd_sc_hd__nand2_1
X_14998_ _15373_/A _15373_/B _15510_/B _15368_/D vssd1 vssd1 vccd1 vccd1 _14998_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_152_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19525_ _19526_/A _19526_/B vssd1 vssd1 vccd1 vccd1 _19640_/B sky130_fd_sc_hd__and2b_1
X_16737_ _16737_/A _16737_/B vssd1 vssd1 vccd1 vccd1 _16738_/C sky130_fd_sc_hd__xnor2_1
X_13949_ _13948_/A _13948_/B _13948_/C _13948_/D vssd1 vssd1 vccd1 vccd1 _13949_/Y
+ sky130_fd_sc_hd__o22ai_2
XFILLER_0_72_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_1000 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19456_ _19456_/A _19456_/B vssd1 vssd1 vccd1 vccd1 _19457_/B sky130_fd_sc_hd__xor2_4
X_16668_ _16668_/A _16668_/B vssd1 vssd1 vccd1 vccd1 _16669_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_146_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18407_ _18281_/D _18282_/B _18405_/X _18552_/B vssd1 vssd1 vccd1 vccd1 _18409_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15619_ _15616_/Y _15617_/X _15477_/Y _15481_/A vssd1 vssd1 vccd1 vccd1 _15619_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19387_ _19387_/A _19387_/B vssd1 vssd1 vccd1 vccd1 _19395_/A sky130_fd_sc_hd__nand2_1
X_16599_ _16599_/A _16599_/B vssd1 vssd1 vccd1 vccd1 _16634_/A sky130_fd_sc_hd__xor2_2
XFILLER_0_57_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18338_ _18789_/A _18773_/B _18338_/C _18338_/D vssd1 vssd1 vccd1 vccd1 _18481_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__13312__C _15217_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19487__B _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18391__B _21361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_969 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18269_ _18270_/A _18270_/B vssd1 vssd1 vccd1 vccd1 _18269_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_142_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20300_ _20301_/A _20301_/B vssd1 vssd1 vccd1 vccd1 _20300_/X sky130_fd_sc_hd__and2_1
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_1039 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21280_ _21280_/A _21280_/B vssd1 vssd1 vccd1 vccd1 _21281_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout5 fanout6/X vssd1 vssd1 vccd1 vccd1 fanout5/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20231_ hold158/X _20230_/X fanout4/X vssd1 vssd1 vccd1 vccd1 hold159/A sky130_fd_sc_hd__mux2_1
XFILLER_0_12_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout102_A _21841_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20162_ _20163_/A _20163_/B vssd1 vssd1 vccd1 vccd1 _20162_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_110_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_20093_ _20093_/A _20235_/A vssd1 vssd1 vccd1 vccd1 _20094_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__14692__A2 _16326_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1083 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_44_clk_i _21822_/CLK vssd1 vssd1 vccd1 vccd1 _21963_/CLK sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout471_A _15091_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_1162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout569_A _12403_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_1146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__19907__A1 _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20995_ _20996_/A _20996_/B vssd1 vssd1 vccd1 vccd1 _20997_/A sky130_fd_sc_hd__nand2_1
XANTENNA__18285__C _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15702__C _16314_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_949 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21616_ _21906_/CLK _21616_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[79] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_30_1032 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_1043 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout15_A wire16/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_1242 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_1076 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21547_ mstream_o[10] hold82/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22074_/D sky130_fd_sc_hd__mux2_1
XANTENNA__18732__D _18894_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_1106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14615__A _15159_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11300_ _13258_/C _11299_/X _11352_/S vssd1 vssd1 vccd1 vccd1 _21776_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12280_ _12207_/X _12210_/Y _12235_/X vssd1 vssd1 vccd1 vccd1 _12280_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_50_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_21478_ hold164/X sstream_i[55] _21481_/S vssd1 vssd1 vccd1 vccd1 _22005_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_132_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12780__D _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11231_ fanout59/X v0z[1] fanout19/X _11230_/X vssd1 vssd1 vccd1 vccd1 _11231_/X
+ sky130_fd_sc_hd__a31o_1
XANTENNA__17449__A2 _17924_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20429_ _21169_/A _21264_/B _21046_/B _21056_/A vssd1 vssd1 vccd1 vccd1 _20433_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_132_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11162_ _12443_/A _11161_/X _11195_/S vssd1 vssd1 vccd1 vccd1 _21737_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_1184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15970_ _15971_/A _15970_/B vssd1 vssd1 vccd1 vccd1 _15970_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__14350__A _15153_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11093_ _11051_/Y hold21/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21687_/D sky130_fd_sc_hd__mux2_1
XANTENNA__21402__A0 _15626_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_1172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14921_ hold102/X _14920_/X fanout4/X vssd1 vssd1 vccd1 vccd1 hold103/A sky130_fd_sc_hd__mux2_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__18149__A1_N _19644_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
X_17640_ _17640_/A _17640_/B vssd1 vssd1 vccd1 vccd1 _17650_/A sky130_fd_sc_hd__xor2_2
Xhold72 hold72/A vssd1 vssd1 vccd1 vccd1 hold72/X sky130_fd_sc_hd__dlygate4sd3_1
X_14852_ _14974_/A _14718_/X _14974_/B _14971_/C vssd1 vssd1 vccd1 vccd1 _14865_/A
+ sky130_fd_sc_hd__o211ai_1
Xhold83 hold83/A vssd1 vssd1 vccd1 vccd1 hold83/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 hold94/A vssd1 vssd1 vccd1 vccd1 hold94/X sky130_fd_sc_hd__dlygate4sd3_1
X_13803_ _13800_/X _13801_/Y _13648_/C _13647_/Y vssd1 vssd1 vccd1 vccd1 _13803_/X
+ sky130_fd_sc_hd__a211o_1
X_14783_ _14783_/A _14783_/B vssd1 vssd1 vccd1 vccd1 _14804_/A sky130_fd_sc_hd__or2_1
X_17571_ _17570_/B _17570_/C _17570_/A vssd1 vssd1 vccd1 vccd1 _17571_/Y sky130_fd_sc_hd__a21oi_2
X_11995_ _11989_/A _11989_/C _11989_/B vssd1 vssd1 vccd1 vccd1 _11996_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_97_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19310_ _19311_/B _19311_/A vssd1 vssd1 vccd1 vccd1 _19467_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_58_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13734_ _13734_/A _13734_/B _13734_/C vssd1 vssd1 vccd1 vccd1 _13734_/Y sky130_fd_sc_hd__nand3_2
X_16522_ _16522_/A _16522_/B _16522_/C vssd1 vssd1 vccd1 vccd1 _16525_/A sky130_fd_sc_hd__nand3_1
XANTENNA__12020__D _12312_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10946_ _10946_/A _10946_/B vssd1 vssd1 vccd1 vccd1 _10946_/Y sky130_fd_sc_hd__nor2_2
XFILLER_0_133_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17385__A1 _17282_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_156_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19241_ _19241_/A _19241_/B _19387_/B vssd1 vssd1 vccd1 vccd1 _19243_/B sky130_fd_sc_hd__nand3_1
X_13665_ fanout9/A _21364_/B vssd1 vssd1 vccd1 vccd1 _13665_/Y sky130_fd_sc_hd__nor2_1
X_16453_ _17029_/A _16968_/C _16743_/C _17029_/B vssd1 vssd1 vccd1 vccd1 _16454_/B
+ sky130_fd_sc_hd__a22o_1
X_10877_ hold157/A hold188/A vssd1 vssd1 vccd1 vccd1 _10885_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_1217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18492__A _19723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15404_ _15404_/A _15404_/B vssd1 vssd1 vccd1 vccd1 _15405_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_128_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12616_ _13394_/A _14176_/C vssd1 vssd1 vccd1 vccd1 _12617_/B sky130_fd_sc_hd__nand2_1
X_16384_ _16384_/A _16384_/B vssd1 vssd1 vccd1 vccd1 _16394_/A sky130_fd_sc_hd__xnor2_2
X_19172_ hold188/X _19171_/X fanout4/X vssd1 vssd1 vccd1 vccd1 _21901_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_26_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_947 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13596_ _13593_/Y _13752_/A _14365_/A _15763_/A vssd1 vssd1 vccd1 vccd1 _13752_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_109_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18334__B1 _19906_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16724__B _17146_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15335_ _15334_/B _15334_/C _15334_/A vssd1 vssd1 vccd1 vccd1 _15336_/C sky130_fd_sc_hd__o21ai_1
X_18123_ _18127_/C _18122_/C _18122_/B vssd1 vssd1 vccd1 vccd1 _18124_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12547_ _12543_/X _12544_/Y _12432_/X _12434_/X vssd1 vssd1 vccd1 vccd1 _12583_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_124_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16443__C _16870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15266_ _15266_/A _15266_/B vssd1 vssd1 vccd1 vccd1 _15268_/B sky130_fd_sc_hd__nand2_1
X_18054_ _18055_/A _18185_/B _18054_/C vssd1 vssd1 vccd1 vccd1 _18181_/A sky130_fd_sc_hd__or3_1
XFILLER_0_35_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12478_ _12475_/Y _12476_/X _12373_/Y _12375_/X vssd1 vssd1 vccd1 vccd1 _12479_/D
+ sky130_fd_sc_hd__o211a_1
XANTENNA_3 _10792_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14244__B _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14217_ _15373_/A _15373_/B _14873_/B _14217_/D vssd1 vssd1 vccd1 vccd1 _14220_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_111_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17005_ _17005_/A _17005_/B _17005_/C vssd1 vssd1 vccd1 vccd1 _17005_/Y sky130_fd_sc_hd__nor3_1
X_11429_ _11447_/A1 hold293/A fanout48/X hold207/A vssd1 vssd1 vccd1 vccd1 _11429_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__18637__A1 _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15197_ _15060_/A _15060_/B _15058_/Y vssd1 vssd1 vccd1 vccd1 _15199_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18637__B2 _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11587__C _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14148_ _14149_/A _14149_/B _14149_/C vssd1 vssd1 vccd1 vccd1 _14148_/X sky130_fd_sc_hd__a21o_1
XANTENNA__21358__A _21420_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11884__A _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14079_ _14076_/X _14231_/B _13921_/X _13924_/A vssd1 vssd1 vccd1 vccd1 _14080_/B
+ sky130_fd_sc_hd__a211o_1
X_18956_ _19587_/B _20242_/C vssd1 vssd1 vccd1 vccd1 _18960_/A sky130_fd_sc_hd__nand2_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17907_ _18026_/A _17906_/C _17906_/A vssd1 vssd1 vccd1 vccd1 _17908_/C sky130_fd_sc_hd__a21o_1
X_18887_ _18760_/Y _18763_/Y _19006_/B _18886_/X vssd1 vssd1 vccd1 vccd1 _18889_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17612__A2 _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17838_ _17830_/A _17837_/B _17705_/X _17830_/B vssd1 vssd1 vccd1 vccd1 _17838_/X
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_1033 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17769_ _17768_/A _17768_/B _17768_/C vssd1 vssd1 vccd1 vccd1 _17770_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_156_1093 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__15091__A _15892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_1128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19508_ _20178_/D _20193_/D _19509_/C _19661_/A vssd1 vssd1 vccd1 vccd1 _19510_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_117_1077 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_20780_ _20912_/A _20780_/B vssd1 vssd1 vccd1 vccd1 _20781_/B sky130_fd_sc_hd__and2_1
XFILLER_0_49_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_1200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19474__C_N _19169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19439_ _19439_/A _20249_/B vssd1 vssd1 vccd1 vccd1 _19441_/C sky130_fd_sc_hd__and2_1
XANTENNA__11660__A2 _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_1244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_925 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14138__C _16084_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17128__A1 _17144_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17128__B2 _17129_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_993 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21401_ hold95/X fanout40/X _21400_/X vssd1 vssd1 vccd1 vccd1 _21941_/D sky130_fd_sc_hd__a21bo_1
XFILLER_0_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20132__B1 _20270_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13977__C _14312_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout317_A _21792_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21332_ _21407_/S _17173_/B _21421_/S vssd1 vssd1 vccd1 vccd1 _21332_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_130_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19945__B fanout8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21263_ _21263_/A _21263_/B vssd1 vssd1 vccd1 vccd1 _21265_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_1037 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19664__C _20733_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_1161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12912__A2 _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20214_ _20215_/A _20215_/B vssd1 vssd1 vccd1 vccd1 _20214_/X sky130_fd_sc_hd__and2b_1
XANTENNA__16103__A2 _16396_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21194_ _21194_/A _21194_/B vssd1 vssd1 vccd1 vccd1 _21196_/B sky130_fd_sc_hd__or2_1
XFILLER_0_60_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_1009 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_20145_ _20562_/B _21305_/A _21153_/B _19906_/A vssd1 vssd1 vccd1 vccd1 _20145_/Y
+ sky130_fd_sc_hd__a22oi_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20076_ _19939_/A _19938_/B _19936_/Y vssd1 vssd1 vccd1 vccd1 _20078_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12402__B _12402_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18800__A1 _19123_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_3437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12428__A1 _12642_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12428__B2 _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__15090__A2 _15091_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10800_ mstream_o[114] mstream_i sstream_o _10792_/Y vssd1 vssd1 vccd1 vccd1 _21716_/D
+ sky130_fd_sc_hd__a22o_1
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13514__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11780_ _12261_/A _13017_/A _12444_/B _12269_/B vssd1 vssd1 vccd1 vccd1 _11781_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__15432__C _15829_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20978_ _20978_/A _21095_/A _20978_/C vssd1 vssd1 vccd1 vccd1 _21091_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_1154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15131__A1_N _15933_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_1127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_1149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19108__A2 _19753_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13450_ _13451_/A _13451_/B _13451_/C vssd1 vssd1 vccd1 vccd1 _13450_/X sky130_fd_sc_hd__a21o_4
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ _12401_/A _12401_/B vssd1 vssd1 vccd1 vccd1 _12408_/A sky130_fd_sc_hd__or2_1
XFILLER_0_91_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12849__A1_N _13682_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13381_ _13378_/Y _13527_/A _13381_/C _16328_/B vssd1 vssd1 vccd1 vccd1 _13527_/B
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__18462__D _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_939 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15120_ _16196_/A _16369_/A _15120_/C _15266_/A vssd1 vssd1 vccd1 vccd1 _15266_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_133_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12332_ _12332_/A _12332_/B vssd1 vssd1 vccd1 vccd1 _12334_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11688__B _12319_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_15051_ _15013_/X _15014_/Y _15050_/C _15050_/D vssd1 vssd1 vccd1 vccd1 _15052_/B
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13156__A2 _13155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_1273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12263_ _12268_/A _12269_/D _12262_/X _12261_/X vssd1 vssd1 vccd1 vccd1 _12264_/C
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_972 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16560__A _16813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14999__B _15373_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14002_ _14002_/A _14002_/B _14002_/C vssd1 vssd1 vccd1 vccd1 _14004_/B sky130_fd_sc_hd__nand3_2
X_11214_ hold175/X fanout51/X fanout48/X hold236/A vssd1 vssd1 vccd1 vccd1 _11214_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12194_ _12193_/B _12193_/C _12193_/A vssd1 vssd1 vccd1 vccd1 _12195_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_120_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18810_ _18810_/A _18810_/B _18810_/C vssd1 vssd1 vccd1 vccd1 _18813_/B sky130_fd_sc_hd__nand3_4
X_11145_ hold231/X _11122_/X fanout45/X hold179/X vssd1 vssd1 vccd1 vccd1 _11145_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19871__A _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19790_ _19169_/B _19788_/Y _19789_/Y vssd1 vssd1 vccd1 vccd1 _19792_/B sky130_fd_sc_hd__a21oi_4
X_18741_ _20317_/D _19382_/B _18741_/C _18741_/D vssd1 vssd1 vccd1 vccd1 _18741_/Y
+ sky130_fd_sc_hd__nand4_1
X_15953_ _16084_/A _21785_/Q _15954_/D _16203_/D vssd1 vssd1 vccd1 vccd1 _15957_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__13408__B _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11076_ _10912_/X hold69/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21671_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19590__B _21171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12312__B _13258_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14904_ _14904_/A _14904_/B vssd1 vssd1 vccd1 vccd1 _14906_/B sky130_fd_sc_hd__xor2_1
X_18672_ _18669_/X _18670_/Y _18516_/C _18515_/Y vssd1 vssd1 vccd1 vccd1 _18674_/D
+ sky130_fd_sc_hd__a211oi_2
X_15884_ _16011_/B _15883_/X _15749_/A _15751_/X vssd1 vssd1 vccd1 vccd1 _16016_/B
+ sky130_fd_sc_hd__o211a_1
X_17623_ _17522_/C _17524_/A _17737_/B _17622_/X vssd1 vssd1 vccd1 vccd1 _17749_/A
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_37_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14835_ _14679_/A _14679_/C _14679_/B vssd1 vssd1 vccd1 vccd1 _14836_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_153_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_1217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17554_ _17657_/A _19439_/A _17551_/Y _17552_/X vssd1 vssd1 vccd1 vccd1 _17555_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_14766_ _14689_/A _14689_/B _14688_/A vssd1 vssd1 vccd1 vccd1 _14806_/A sky130_fd_sc_hd__a21oi_2
X_11978_ _11976_/A _11977_/X _11905_/Y _11910_/X vssd1 vssd1 vccd1 vccd1 _12388_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_86_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18934__B _19092_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16505_ _16553_/A _16505_/B vssd1 vssd1 vccd1 vccd1 _16715_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_156_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13717_ _13718_/A _13718_/B vssd1 vssd1 vccd1 vccd1 _13846_/B sky130_fd_sc_hd__or2_1
X_10929_ hold109/A hold158/A vssd1 vssd1 vccd1 vccd1 _10931_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_129_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_14697_ _21768_/Q _16266_/C _14698_/D _15514_/A vssd1 vssd1 vccd1 vccd1 _14702_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__11642__A2 _12403_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17485_ hold125/A fanout7/X _17484_/X _11550_/A _17378_/Y vssd1 vssd1 vccd1 vccd1
+ _17485_/X sky130_fd_sc_hd__a221o_1
XFILLER_0_86_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_1183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19111__A _19432_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19224_ _19224_/A _19224_/B vssd1 vssd1 vccd1 vccd1 _19234_/A sky130_fd_sc_hd__xor2_1
X_16436_ _16436_/A _16436_/B vssd1 vssd1 vccd1 vccd1 _16437_/B sky130_fd_sc_hd__xnor2_4
X_13648_ _13648_/A _13648_/B _13648_/C _13648_/D vssd1 vssd1 vccd1 vccd1 _13648_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_6_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19155_ _18991_/B _19155_/B vssd1 vssd1 vccd1 vccd1 _19157_/B sky130_fd_sc_hd__and2b_1
XANTENNA__18858__A1 _18859_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16367_ _16361_/B _16362_/A _16366_/X _16360_/B vssd1 vssd1 vccd1 vccd1 _16437_/A
+ sky130_fd_sc_hd__a211o_1
X_13579_ _13580_/A _13580_/B _13580_/C vssd1 vssd1 vccd1 vccd1 _13581_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_6_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18106_ _18106_/A vssd1 vssd1 vccd1 vccd1 _18234_/A sky130_fd_sc_hd__inv_2
XFILLER_0_48_1123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15318_ _16092_/D _15717_/C _15976_/D _15961_/D vssd1 vssd1 vccd1 vccd1 _15318_/Y
+ sky130_fd_sc_hd__a22oi_1
XFILLER_0_54_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16298_ _16298_/A _16298_/B vssd1 vssd1 vccd1 vccd1 _16300_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_81_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19086_ _20101_/B _19705_/B _19546_/D _20101_/A vssd1 vssd1 vccd1 vccd1 _19088_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_1145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17530__A1 _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_1047 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18037_ _17901_/A _17901_/C _17901_/B vssd1 vssd1 vccd1 vccd1 _18038_/C sky130_fd_sc_hd__a21bo_1
XFILLER_0_23_961 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15249_ _15249_/A _15249_/B vssd1 vssd1 vccd1 vccd1 _15252_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_78_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__16470__A _17300_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout307 _21794_/Q vssd1 vssd1 vccd1 vccd1 _19337_/D sky130_fd_sc_hd__buf_4
Xfanout318 _17493_/A vssd1 vssd1 vccd1 vccd1 _17146_/C sky130_fd_sc_hd__buf_4
Xfanout329 _16404_/B vssd1 vssd1 vccd1 vccd1 _15698_/B sky130_fd_sc_hd__buf_4
X_19988_ _21199_/A _20838_/B _20265_/D vssd1 vssd1 vccd1 vccd1 _19988_/X sky130_fd_sc_hd__and3_1
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_1020 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_18939_ _18938_/A _18938_/B _18938_/C vssd1 vssd1 vccd1 vccd1 _18940_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21950_ _21963_/CLK _21950_/D vssd1 vssd1 vccd1 vccd1 hold225/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_27_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__18794__B1 _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17597__B2 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20901_ _20901_/A _20901_/B _20902_/B _20643_/A vssd1 vssd1 vccd1 vccd1 _20904_/B
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_96_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21881_ _21945_/CLK hold37/X vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_55_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14938__A1_N _21733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout267_A _21802_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20832_ _20667_/B _20710_/A _20830_/Y _20831_/X vssd1 vssd1 vccd1 vccd1 _21016_/A
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_76_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11094__A0 _11053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11633__A2 _12619_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20763_ _20596_/Y _20601_/A _20896_/A _20762_/X vssd1 vssd1 vccd1 vccd1 _20896_/B
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_77_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout434_A _21762_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20694_ _20694_/A _20694_/B vssd1 vssd1 vccd1 vccd1 _20696_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_135_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_1085 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19378__D _19691_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout601_A _11459_/B2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20105__B1 _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20317__D _20317_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17521__A1 _17520_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17521__B2 _17520_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21315_ _21056_/A _21169_/A _10796_/Y _21056_/B vssd1 vssd1 vccd1 vccd1 _21316_/B
+ sky130_fd_sc_hd__o211a_1
XANTENNA__16380__A _16380_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21246_ _21246_/A _21246_/B vssd1 vssd1 vccd1 vccd1 _21248_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__21581__RESET_B _11089_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20333__C _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19691__A _21199_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21177_ _21178_/A _21178_/B vssd1 vssd1 vccd1 vccd1 _21179_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_102_1132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout82_A _21846_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_1065 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20128_ _21199_/A _20863_/C _21278_/A _20265_/D vssd1 vssd1 vccd1 vccd1 _20330_/A
+ sky130_fd_sc_hd__nand4_2
XANTENNA__13310__A2 _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18738__C _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12950_ _13091_/A _12950_/B _12950_/C vssd1 vssd1 vccd1 vccd1 _12951_/B sky130_fd_sc_hd__and3_1
XTAP_3201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20059_ _20059_/A _20167_/A _20059_/C vssd1 vssd1 vccd1 vccd1 _20167_/B sky130_fd_sc_hd__nor3_1
XTAP_3212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11321__A1 _11325_/A1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17642__C _18622_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11321__B2 _21723_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11901_ _11901_/A _11901_/B _11901_/C vssd1 vssd1 vccd1 vccd1 _11901_/X sky130_fd_sc_hd__and3_2
XTAP_3234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ _13013_/A _13157_/B vssd1 vssd1 vccd1 vccd1 _12884_/A sky130_fd_sc_hd__and2_1
XTAP_3256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20592__B1 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_201 hold268/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_212 hold275/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_223 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14620_ _14620_/A _14620_/B vssd1 vssd1 vccd1 vccd1 _14625_/A sky130_fd_sc_hd__xnor2_2
X_11832_ _11826_/Y _11829_/X _11831_/Y _11801_/X vssd1 vssd1 vccd1 vccd1 _11836_/A
+ sky130_fd_sc_hd__o211ai_4
XANTENNA_234 hold299/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_245 _11347_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11085__A0 _10972_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_256 v2z[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_267 hold288/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14551_ _14551_/A _14551_/B _14551_/C vssd1 vssd1 vccd1 vccd1 _14553_/A sky130_fd_sc_hd__and3_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_278 hold283/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18001__A2 _19060_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11763_ _11763_/A _11763_/B vssd1 vssd1 vccd1 vccd1 _11764_/C sky130_fd_sc_hd__xnor2_2
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_289 hold274/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16555__A _16870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_839 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13502_ _13523_/B _13501_/B _13500_/C _13500_/D vssd1 vssd1 vccd1 vccd1 _13502_/Y
+ sky130_fd_sc_hd__a2bb2oi_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13898__B _15514_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14482_ _14482_/A _14482_/B _14482_/C vssd1 vssd1 vccd1 vccd1 _14484_/B sky130_fd_sc_hd__nand3_2
X_17270_ _17372_/A _16912_/Y _17171_/A _17171_/B vssd1 vssd1 vccd1 vccd1 _17381_/B
+ sky130_fd_sc_hd__o22a_4
XFILLER_0_67_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11694_ _12426_/B _12619_/A _12330_/A _11694_/D vssd1 vssd1 vccd1 vccd1 _12330_/B
+ sky130_fd_sc_hd__nand4_1
XANTENNA__17760__A1 _18767_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16221_ _16221_/A _16221_/B vssd1 vssd1 vccd1 vccd1 _16223_/B sky130_fd_sc_hd__xnor2_1
X_13433_ _13280_/A _13280_/Y _13430_/X _13431_/Y vssd1 vssd1 vccd1 vccd1 _13433_/Y
+ sky130_fd_sc_hd__o211ai_4
XANTENNA__13377__A2 _13997_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19866__A _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14075__A _14848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16152_ _16152_/A _16152_/B vssd1 vssd1 vccd1 vccd1 _16191_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20647__B2 _11547_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13364_ _13091_/A _13087_/X _13223_/A vssd1 vssd1 vccd1 vccd1 _13365_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15103_ _15103_/A _15226_/B _15103_/C vssd1 vssd1 vccd1 vccd1 _15254_/A sky130_fd_sc_hd__and3_1
XANTENNA__13129__A2 _15768_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12315_ _12315_/A _12315_/B vssd1 vssd1 vccd1 vccd1 _12317_/A sky130_fd_sc_hd__xnor2_2
X_16083_ _16196_/A _16084_/C _16084_/D _16084_/A vssd1 vssd1 vccd1 vccd1 _16087_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13295_ _13293_/Y _13445_/A _14195_/A _15763_/A vssd1 vssd1 vccd1 vccd1 _13445_/B
+ sky130_fd_sc_hd__and4bb_1
XANTENNA__14877__A2 _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15034_ _15933_/C _16409_/A _15034_/C _15127_/A vssd1 vssd1 vccd1 vccd1 _15127_/B
+ sky130_fd_sc_hd__nand4_1
X_19911_ _19911_/A _19911_/B _19911_/C vssd1 vssd1 vccd1 vccd1 _19914_/A sky130_fd_sc_hd__nand3_1
X_12246_ _12261_/A _12269_/B _12246_/C _12246_/D vssd1 vssd1 vccd1 vccd1 _12249_/C
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_139_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_1087 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17276__B1 _21258_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19842_ _19843_/A _19843_/B vssd1 vssd1 vccd1 vccd1 _19842_/X sky130_fd_sc_hd__and2b_1
XFILLER_0_102_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12177_ _12160_/A _12160_/C _12160_/B vssd1 vssd1 vccd1 vccd1 _12177_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_1075 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__18929__B _18929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11128_ hold160/X fanout23/X _11127_/X vssd1 vssd1 vccd1 vccd1 _11128_/X sky130_fd_sc_hd__a21o_1
XANTENNA__17833__B _21349_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19773_ _19773_/A _19773_/B vssd1 vssd1 vccd1 vccd1 _19776_/A sky130_fd_sc_hd__xor2_1
X_16985_ _16986_/A _16986_/B vssd1 vssd1 vccd1 vccd1 _16999_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_78_1138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18724_ _18721_/Y _18722_/X _18563_/Y _18566_/X vssd1 vssd1 vccd1 vccd1 _18725_/C
+ sky130_fd_sc_hd__o211a_1
X_15936_ _15936_/A _15936_/B vssd1 vssd1 vccd1 vccd1 _15938_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__21355__B _21355_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11059_ _11059_/A _11059_/B vssd1 vssd1 vccd1 vccd1 _11059_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__18010__A _18010_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21375__A2 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18655_ _18500_/A _18500_/C _18500_/B vssd1 vssd1 vccd1 vccd1 _18656_/C sky130_fd_sc_hd__a21bo_1
X_15867_ _15867_/A _15867_/B _15867_/C vssd1 vssd1 vccd1 vccd1 _15952_/B sky130_fd_sc_hd__or3_1
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11863__A2 _12621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_1161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17606_ _18857_/B _18703_/A _21151_/A _18894_/B vssd1 vssd1 vccd1 vccd1 _17715_/A
+ sky130_fd_sc_hd__and4_2
XANTENNA__19339__A1_N _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14818_ _16203_/D _15022_/B _14820_/C _14820_/D vssd1 vssd1 vccd1 vccd1 _14818_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_153_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_942 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18586_ _18583_/Y _18584_/X _19644_/A _19060_/B vssd1 vssd1 vccd1 vccd1 _18587_/B
+ sky130_fd_sc_hd__and4bb_1
XTAP_3790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_15798_ _15798_/A _15798_/B vssd1 vssd1 vccd1 vccd1 _15800_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_87_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11076__A0 _10912_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17537_ _17422_/X _17424_/X _17535_/X _17536_/Y vssd1 vssd1 vccd1 vccd1 _17575_/A
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_59_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14749_ _14750_/B _14750_/A vssd1 vssd1 vccd1 vccd1 _14749_/Y sky130_fd_sc_hd__nand2b_1
XFILLER_0_15_1133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11615__A2 _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12993__A _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_1177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17468_ _17356_/C _17355_/Y _17466_/X _17467_/Y vssd1 vssd1 vccd1 vccd1 _17468_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_50_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19207_ _19206_/B _19206_/C _19195_/Y vssd1 vssd1 vccd1 vccd1 _19207_/Y sky130_fd_sc_hd__a21boi_1
X_16419_ _16278_/A _16278_/B _16276_/Y vssd1 vssd1 vccd1 vccd1 _16420_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_104_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_958 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17399_ _17400_/A _17400_/B vssd1 vssd1 vccd1 vccd1 _17512_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19138_ _19135_/X _19136_/Y _18975_/B _18975_/Y vssd1 vssd1 vccd1 vccd1 _19139_/C
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13320__C _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17503__A1 _17619_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17503__B2 _17621_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_933 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19069_ _19379_/B _19240_/B _19070_/C _19235_/A vssd1 vssd1 vccd1 vccd1 _19071_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14713__A _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_1121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_977 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21100_ _21208_/A vssd1 vssd1 vccd1 vccd1 _21102_/D sky130_fd_sc_hd__inv_2
XFILLER_0_1_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_22080_ _22080_/CLK _22080_/D fanout636/X vssd1 vssd1 vccd1 vccd1 mstream_o[16] sky130_fd_sc_hd__dfrtp_4
XANTENNA__19256__A1 _20101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15528__B _15529_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12879__A1 _13152_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__19256__B2 _20101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_1007 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21031_ _20918_/A _20918_/B _20788_/A vssd1 vssd1 vccd1 vccd1 _21035_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_10_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout104 _19691_/D vssd1 vssd1 vccd1 vccd1 _19057_/D sky130_fd_sc_hd__buf_2
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout115 _20148_/C vssd1 vssd1 vccd1 vccd1 _19240_/B sky130_fd_sc_hd__buf_4
Xfanout126 _21837_/Q vssd1 vssd1 vccd1 vccd1 _20689_/A sky130_fd_sc_hd__buf_4
XFILLER_0_22_1137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__20810__A1 _20562_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout137 _21834_/Q vssd1 vssd1 vccd1 vccd1 _20774_/A sky130_fd_sc_hd__clkbuf_8
XANTENNA__13048__B _14391_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20810__B2 _21056_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout148 _19092_/B vssd1 vssd1 vccd1 vccd1 _20394_/B sky130_fd_sc_hd__buf_6
XFILLER_0_129_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout159 _16743_/B vssd1 vssd1 vccd1 vccd1 _17029_/B sky130_fd_sc_hd__buf_4
XANTENNA_fanout384_A _16173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16490__A1 _17636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__21366__A2 fanout40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21933_ _21942_/CLK _21933_/D vssd1 vssd1 vccd1 vccd1 hold118/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_fanout551_A _21733_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17181__D _17739_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21864_ _21932_/CLK _21864_/D vssd1 vssd1 vccd1 vccd1 hold88/A sky130_fd_sc_hd__dfxtp_1
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11067__A0 _11066_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13999__A _14306_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20815_ _20815_/A _20938_/B vssd1 vssd1 vccd1 vccd1 _20817_/B sky130_fd_sc_hd__or2_1
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_132_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_986 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_1233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21795_ _22020_/CLK _21795_/D vssd1 vssd1 vccd1 vccd1 _21795_/Q sky130_fd_sc_hd__dfxtp_4
XFILLER_0_65_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19731__A2 _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20746_ _20743_/Y _20744_/X _20615_/X _20617_/X vssd1 vssd1 vccd1 vccd1 _20747_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17742__A1 _21796_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__14556__A1 _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__14556__B2 _14557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19686__A _19686_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20677_ _21256_/A _21040_/A _20677_/C _20677_/D vssd1 vssd1 vccd1 vccd1 _20801_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__14326__C _14477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19495__B2 _18849_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_991 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_1004 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__17637__C _18616_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_977 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12100_ _12100_/A _12100_/B _12100_/C vssd1 vssd1 vccd1 vccd1 _12150_/A sky130_fd_sc_hd__nand3_1
XANTENNA__16541__C _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_1097 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13080_ _13083_/B vssd1 vssd1 vccd1 vccd1 _13080_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_131_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11458__S _11470_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ _12036_/A _12036_/B _12036_/C vssd1 vssd1 vccd1 vccd1 _12286_/C sky130_fd_sc_hd__a21oi_2
X_21229_ _21229_/A _21229_/B vssd1 vssd1 vccd1 vccd1 _21230_/B sky130_fd_sc_hd__nor2_1
Xhold180 hold180/A vssd1 vssd1 vccd1 vccd1 hold180/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 hold191/A vssd1 vssd1 vccd1 vccd1 hold191/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12143__A _12267_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19852__C _20247_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11542__A1 _19185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18749__B _19686_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19571__D _19874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16770_ _16838_/A _16838_/B vssd1 vssd1 vccd1 vccd1 _16770_/X sky130_fd_sc_hd__and2_1
X_13982_ _14133_/D _16404_/B _16406_/B _13983_/B vssd1 vssd1 vccd1 vccd1 _13985_/C
+ sky130_fd_sc_hd__a22oi_2
XANTENNA__21357__A2 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15721_ _15722_/B _15722_/A vssd1 vssd1 vccd1 vccd1 _15721_/Y sky130_fd_sc_hd__nand2b_1
XTAP_3020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12933_ _12929_/X _12930_/Y _12803_/C _12802_/Y vssd1 vssd1 vccd1 vccd1 _12934_/D
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_73_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_1144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18440_ _18440_/A _18440_/B vssd1 vssd1 vccd1 vccd1 _18441_/B sky130_fd_sc_hd__nand2_1
X_15652_ _16399_/A _15911_/A _15911_/C _16305_/B vssd1 vssd1 vccd1 vccd1 _15655_/C
+ sky130_fd_sc_hd__a22o_1
XTAP_3075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_150_1203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_3086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ _12862_/X _12864_/B vssd1 vssd1 vccd1 vccd1 _12865_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_69_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11058__A0 _11057_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18484__B _19732_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14603_ _14911_/A _14603_/B _14603_/C vssd1 vssd1 vccd1 vccd1 _14604_/B sky130_fd_sc_hd__nor3_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18371_ _18368_/X _18369_/Y _18220_/C _18219_/Y vssd1 vssd1 vccd1 vccd1 _18373_/D
+ sky130_fd_sc_hd__a211oi_2
X_11815_ _11815_/A _11815_/B vssd1 vssd1 vccd1 vccd1 _11816_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_56_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_15583_ _15443_/A _15442_/A _15442_/B _15438_/B _15438_/A vssd1 vssd1 vccd1 vccd1
+ _15585_/B sky130_fd_sc_hd__o32ai_4
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12795_ _12795_/A _12795_/B _12795_/C vssd1 vssd1 vccd1 vccd1 _12798_/B sky130_fd_sc_hd__nand3_4
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_327 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17322_ _17236_/A _17235_/A _17235_/B vssd1 vssd1 vccd1 vccd1 _17329_/A sky130_fd_sc_hd__o21ba_1
XANTENNA__19722__A2 _20247_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_14534_ _14212_/B _16328_/A _16326_/A _14993_/A vssd1 vssd1 vccd1 vccd1 _14534_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_84_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11746_ _12781_/D _12443_/A _11709_/A _11707_/Y vssd1 vssd1 vccd1 vccd1 _11747_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_141_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17253_ _16634_/B _16634_/Y _17250_/X _17252_/Y vssd1 vssd1 vccd1 vccd1 _17256_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_71_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14465_ _14463_/D _16406_/B _16374_/B _14312_/D vssd1 vssd1 vccd1 vccd1 _14466_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_43_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11677_ _12223_/A _12877_/B _11676_/B _11673_/X vssd1 vssd1 vccd1 vccd1 _11682_/A
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16204_ _16203_/D _16406_/B _16374_/B _15695_/A vssd1 vssd1 vccd1 vccd1 _16205_/B
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_52_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13416_ _13416_/A _13416_/B vssd1 vssd1 vccd1 vccd1 _13425_/A sky130_fd_sc_hd__or2_1
XFILLER_0_10_1052 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14396_ _14532_/A _14395_/C _14395_/A vssd1 vssd1 vccd1 vccd1 _14398_/C sky130_fd_sc_hd__a21o_1
X_17184_ _17277_/A _17741_/B _17183_/C _17183_/D vssd1 vssd1 vccd1 vccd1 _17185_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__19486__A1 _19487_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19486__B2 _19487_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_1029 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16135_ _16001_/X _16003_/Y _16133_/Y _16134_/X vssd1 vssd1 vccd1 vccd1 _16251_/A
+ sky130_fd_sc_hd__a211oi_4
X_13347_ _13348_/A _13348_/B _13348_/C vssd1 vssd1 vccd1 vccd1 _13347_/Y sky130_fd_sc_hd__nor3_2
XFILLER_0_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_18_clk_i_A clkbuf_2_3__f_clk_i/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_1006 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_1186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_16066_ _16064_/X _16066_/B vssd1 vssd1 vccd1 vccd1 _16067_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_110_925 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13278_ _13427_/B _13278_/B _13278_/C vssd1 vssd1 vccd1 vccd1 _13280_/A sky130_fd_sc_hd__and3_2
XFILLER_0_59_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21045__A1 _21256_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11368__S _11401_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15017_ _15017_/A _15017_/B vssd1 vssd1 vccd1 vccd1 _15019_/A sky130_fd_sc_hd__nand2_1
X_12229_ _12229_/A _12269_/D vssd1 vssd1 vccd1 vccd1 _12232_/A sky130_fd_sc_hd__nand2_1
XANTENNA__11533__A1 _19013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15592__A1_N _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19825_ _20462_/D _20193_/D _19825_/C _20043_/A vssd1 vssd1 vccd1 vccd1 _20043_/B
+ sky130_fd_sc_hd__nand4_2
XANTENNA__18461__A2 _18929_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20270__A _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_1073 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19756_ _19756_/A _19756_/B _19756_/C vssd1 vssd1 vccd1 vccd1 _19758_/B sky130_fd_sc_hd__nand3_2
X_16968_ _17141_/A _17141_/B _16968_/C _17013_/C vssd1 vssd1 vccd1 vccd1 _16971_/A
+ sky130_fd_sc_hd__nand4_1
XANTENNA__21348__A2 _21381_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18707_ _18707_/A _18707_/B vssd1 vssd1 vccd1 vccd1 _18708_/B sky130_fd_sc_hd__nor2_1
X_15919_ _16369_/A _16396_/A _15919_/C _15919_/D vssd1 vssd1 vccd1 vccd1 _16050_/B
+ sky130_fd_sc_hd__and4_1
X_19687_ fanout96/X _19686_/X _19685_/X vssd1 vssd1 vccd1 vccd1 _19689_/A sky130_fd_sc_hd__a21bo_1
X_16899_ _17041_/A _16899_/B _17493_/A _18859_/A vssd1 vssd1 vccd1 vccd1 _16997_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_155_1169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18638_ _19732_/A _18787_/B _19092_/C _19262_/C vssd1 vssd1 vccd1 vccd1 _18784_/A
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_59_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11049__A0 _11048_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17972__B2 _11550_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14786__A1 _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_1064 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18569_ _18572_/B vssd1 vssd1 vccd1 vccd1 _18569_/Y sky130_fd_sc_hd__inv_2
XANTENNA__13034__D _13034_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__20859__A1 _21296_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20600_ _20600_/A _20600_/B vssd1 vssd1 vccd1 vccd1 _20601_/B sky130_fd_sc_hd__or2_1
XANTENNA__20859__B2 _20991_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21580_ _22106_/CLK _21580_/D fanout637/X vssd1 vssd1 vccd1 vccd1 mstream_o[43] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_129_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_1053 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__20148__C _20148_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20531_ _20914_/A _20531_/B vssd1 vssd1 vccd1 vccd1 _20533_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_156_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout132_A _19087_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_1205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20462_ _18008_/A _21293_/B _20721_/C _20462_/D vssd1 vssd1 vccd1 vccd1 _20600_/A
+ sky130_fd_sc_hd__and4b_2
XANTENNA__19477__B2 _19636_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_1216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__15539__A _16369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13761__A2 _14557_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20393_ _20650_/A _21171_/B vssd1 vssd1 vccd1 vccd1 _20397_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_936 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__21036__A1 _21301_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout599_A _16363_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_22063_ _22063_/CLK _22063_/D vssd1 vssd1 vccd1 vccd1 hold283/A sky130_fd_sc_hd__dfxtp_4
XANTENNA__21036__B2 _21151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11524__A1 _19199_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21014_ _21014_/A _21014_/B vssd1 vssd1 vccd1 vccd1 _21016_/C sky130_fd_sc_hd__and2_1
XFILLER_0_96_1002 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15274__A _15931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__21339__A2 _21421_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11288__A0 _12858_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17412__B1 _20774_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19952__A2 _19951_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13823__A2_N _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21916_ _21948_/CLK hold172/X vssd1 vssd1 vccd1 vccd1 hold171/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_136_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21847_ _21853_/CLK _21847_/D vssd1 vssd1 vccd1 vccd1 _21847_/Q sky130_fd_sc_hd__dfxtp_4
XANTENNA__15974__B1 _16418_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_1041 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11600_ _12426_/B _12402_/A _11599_/B _11596_/X vssd1 vssd1 vccd1 vccd1 _11602_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_66_945 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12580_ _12471_/B _12471_/Y _12577_/X _12579_/Y vssd1 vssd1 vccd1 vccd1 _12583_/C
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_37_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21778_ _21816_/CLK _21778_/D vssd1 vssd1 vccd1 vccd1 _21778_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11531_ _11089_/B t1y[27] t0x[27] _11223_/A vssd1 vssd1 vccd1 vccd1 _11531_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_147_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20729_ _20729_/A _20729_/B vssd1 vssd1 vccd1 vccd1 _20740_/A sky130_fd_sc_hd__or2_1
XANTENNA__17929__A _21824_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_1126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14250_ _14572_/A _14250_/B vssd1 vssd1 vccd1 vccd1 _14251_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11462_ _11123_/A t1y[4] t0x[4] _21724_/D vssd1 vssd1 vccd1 vccd1 _11462_/X sky130_fd_sc_hd__a22o_1
XFILLER_0_135_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13201_ _13062_/B _13062_/Y _13198_/X _13200_/Y vssd1 vssd1 vccd1 vccd1 _13204_/B
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_33_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_14181_ _14508_/A _14813_/A _14354_/C _14817_/D vssd1 vssd1 vccd1 vccd1 _14181_/X
+ sky130_fd_sc_hd__and4_1
X_11393_ _11124_/A hold254/X _11126_/B hold170/X vssd1 vssd1 vccd1 vccd1 _11393_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__14353__A _15695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16271__C _16369_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13132_ _13858_/B _13573_/D _13267_/A _13132_/D vssd1 vssd1 vccd1 vccd1 _13267_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_0_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_1013 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__17086__D _17123_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_1035 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13063_ _13062_/B _13062_/C _13062_/A vssd1 vssd1 vccd1 vccd1 _13063_/Y sky130_fd_sc_hd__a21oi_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17940_ _17940_/A _17940_/B _17940_/C vssd1 vssd1 vccd1 vccd1 _17943_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_44_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11515__A1 _18732_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ _12009_/A _12009_/B _12002_/X vssd1 vssd1 vccd1 vccd1 _12017_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__12712__B1 _11053_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17871_ _18008_/B _18769_/B _17759_/X _17758_/X _18767_/B vssd1 vssd1 vccd1 vccd1
+ _17876_/A sky130_fd_sc_hd__a32o_1
XANTENNA__18443__A2 _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13119__D _21777_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_19610_ _19449_/A _19449_/B _19447_/X vssd1 vssd1 vccd1 vccd1 _19612_/B sky130_fd_sc_hd__a21oi_4
X_16822_ _16822_/A _16822_/B vssd1 vssd1 vccd1 vccd1 _16823_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__12601__A fanout9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14465__B1 _16374_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout490 _21746_/Q vssd1 vssd1 vccd1 vccd1 _14384_/C sky130_fd_sc_hd__clkbuf_8
XANTENNA__11279__B1 _11278_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19541_ _19539_/X _19541_/B vssd1 vssd1 vccd1 vccd1 _19542_/B sky130_fd_sc_hd__nand2b_1
X_16753_ _16753_/A _16753_/B vssd1 vssd1 vccd1 vccd1 _16754_/C sky130_fd_sc_hd__xor2_2
X_13965_ _13664_/A _14294_/B vssd1 vssd1 vccd1 vccd1 _13966_/B sky130_fd_sc_hd__and2b_1
X_15704_ _15702_/D _15838_/B _16374_/B _15435_/A vssd1 vssd1 vccd1 vccd1 _15705_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_12916_ _12916_/A _12916_/B _12916_/C vssd1 vssd1 vccd1 vccd1 _12918_/B sky130_fd_sc_hd__nand3_1
XANTENNA__18746__A3 _19068_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19472_ _19472_/A _19472_/B vssd1 vssd1 vccd1 vccd1 _19476_/A sky130_fd_sc_hd__xnor2_2
X_16684_ _16686_/B vssd1 vssd1 vccd1 vccd1 _16684_/Y sky130_fd_sc_hd__inv_2
X_13896_ _13896_/A _13896_/B vssd1 vssd1 vccd1 vccd1 _13904_/A sky130_fd_sc_hd__xor2_1
X_18423_ _18543_/B _18421_/X _18307_/X _18310_/Y vssd1 vssd1 vccd1 vccd1 _18423_/X
+ sky130_fd_sc_hd__o211a_1
X_15635_ _16027_/A _16369_/B _15635_/C _15635_/D vssd1 vssd1 vccd1 vccd1 _15803_/B
+ sky130_fd_sc_hd__and4_1
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ _12848_/B vssd1 vssd1 vccd1 vccd1 _12847_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_69_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__20249__B _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_1175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12779__B1 _14386_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_1261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18354_ _18204_/A _18204_/C _18204_/B vssd1 vssd1 vccd1 vccd1 _18355_/C sky130_fd_sc_hd__a21bo_1
X_15566_ _15563_/Y _15564_/X _15420_/B _15420_/Y vssd1 vssd1 vccd1 vccd1 _15567_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_967 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12778_ _12778_/A _12778_/B vssd1 vssd1 vccd1 vccd1 _12798_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14247__B _21759_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_17305_ _17393_/B _17305_/B vssd1 vssd1 vccd1 vccd1 _17315_/A sky130_fd_sc_hd__nor2_1
X_14517_ _14365_/A _15808_/C _14518_/C _14671_/A vssd1 vssd1 vccd1 vccd1 _14519_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_1147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18285_ _19644_/A _19487_/A _19227_/C _19227_/D vssd1 vssd1 vccd1 vccd1 _18286_/B
+ sky130_fd_sc_hd__nand4_1
X_11729_ _12458_/A _12357_/C _13155_/A _13155_/B vssd1 vssd1 vccd1 vccd1 _11732_/A
+ sky130_fd_sc_hd__nand4_2
X_15497_ _15625_/B _15497_/B vssd1 vssd1 vccd1 vccd1 _21399_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16743__A _16813_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17182__A2 _17739_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_674 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17236_ _17236_/A _17236_/B vssd1 vssd1 vccd1 vccd1 _17245_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_142_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14448_ _14448_/A _14601_/B vssd1 vssd1 vccd1 vccd1 _14449_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__20265__A _20863_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17167_ _17167_/A _17167_/B vssd1 vssd1 vccd1 vccd1 _17168_/C sky130_fd_sc_hd__xnor2_1
XANTENNA__10791__A _11122_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14379_ _14379_/A _14379_/B _14379_/C vssd1 vssd1 vccd1 vccd1 _14381_/A sky130_fd_sc_hd__and3_1
XANTENNA__17277__C _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16118_ _16115_/Y _16116_/X _15985_/X _15987_/X vssd1 vssd1 vccd1 vccd1 _16119_/C
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_122_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17098_ _17091_/A _17091_/B _17091_/C vssd1 vssd1 vccd1 vccd1 _17099_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_10_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16049_ _16049_/A _16165_/B vssd1 vssd1 vccd1 vccd1 _16052_/A sky130_fd_sc_hd__or2_1
XFILLER_0_0_953 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_1270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11506__A1 _19227_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12214__C _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15806__B _15931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20241__A2 _20242_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20431__C _21264_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19808_ _19808_/A _19808_/B _19808_/C vssd1 vssd1 vccd1 vccd1 _19809_/B sky130_fd_sc_hd__and3_1
XANTENNA__13259__A1 _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12511__A _12511_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14456__B1 _16084_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13259__B2 _13860_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__16996__A2 _17493_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11809__A2 _12444_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19739_ _19740_/A _19740_/B _19740_/C _19740_/D vssd1 vssd1 vccd1 vccd1 _19743_/A
+ sky130_fd_sc_hd__a22o_1
XANTENNA__16918__A _17145_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16637__B _17433_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21701_ _22096_/CLK _21701_/D vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_149_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19013__B _19337_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_1275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_21632_ _21682_/CLK _21632_/D fanout644/X vssd1 vssd1 vccd1 vccd1 mstream_o[95] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_978 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__14157__B _16328_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13982__A2 _16404_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_21563_ mstream_o[26] hold12/X _21579_/S vssd1 vssd1 vccd1 vccd1 _22090_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout514_A _21741_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20514_ _20643_/B _20514_/B vssd1 vssd1 vccd1 vccd1 _20514_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_0_132_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21494_ hold149/X sstream_i[71] _21494_/S vssd1 vssd1 vccd1 vccd1 _22021_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_43_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__20606__C _21283_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20445_ _20446_/A _20446_/B vssd1 vssd1 vccd1 vccd1 _20445_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_1057 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_1154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20376_ _20643_/A _20901_/A vssd1 vssd1 vccd1 vccd1 _20377_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19870__A1 _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19870__B2 _19972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__14312__A_N _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__17915__C _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_22046_ _22049_/CLK _22046_/D vssd1 vssd1 vccd1 vccd1 hold234/A sky130_fd_sc_hd__dfxtp_4
XFILLER_0_134_1017 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13750_ _15763_/A _14365_/D _13750_/C _13750_/D vssd1 vssd1 vccd1 vccd1 _13751_/B
+ sky130_fd_sc_hd__nand4_2
X_10962_ hold36/A hold145/A vssd1 vssd1 vccd1 vccd1 _10967_/C sky130_fd_sc_hd__or2_1
XFILLER_0_138_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13670__A1 _14133_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13670__B2 _13983_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12701_ _12701_/A _12701_/B _12701_/C vssd1 vssd1 vccd1 vccd1 _12701_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_70_1016 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__14993__D _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13681_ _13682_/C _16328_/B _13679_/Y _13835_/A vssd1 vssd1 vccd1 vccd1 _13681_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_10893_ mstream_o[49] _10892_/Y _10992_/S vssd1 vssd1 vccd1 vccd1 _21586_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14348__A _14659_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_15420_ _15420_/A _15420_/B _15420_/C vssd1 vssd1 vccd1 vccd1 _15420_/Y sky130_fd_sc_hd__nand3_2
XANTENNA__16266__C _16266_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_956 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12632_ _12630_/B _12630_/C _12630_/A vssd1 vssd1 vccd1 vccd1 _12632_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_0_38_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_989 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15351_ _15351_/A _15351_/B vssd1 vssd1 vccd1 vccd1 _15354_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__17659__A _19892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12563_ _12563_/A _12563_/B vssd1 vssd1 vccd1 vccd1 _12572_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_1101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13402__D _13402_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14302_ _14171_/A _14303_/B _14170_/B _14172_/Y vssd1 vssd1 vccd1 vccd1 _14439_/A
+ sky130_fd_sc_hd__o31ai_4
X_11514_ _11224_/A t2x[21] v1z[21] fanout21/X _11513_/X vssd1 vssd1 vccd1 vccd1 _11514_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_1072 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18070_ _18069_/A _18069_/B _18069_/C vssd1 vssd1 vccd1 vccd1 _18071_/C sky130_fd_sc_hd__a21o_1
XFILLER_0_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15282_ _15282_/A _15282_/B vssd1 vssd1 vccd1 vccd1 _15284_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_124_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12494_ _21725_/D hold193/A _11048_/Y fanout6/X _12493_/Y vssd1 vssd1 vccd1 vccd1
+ _12494_/X sky130_fd_sc_hd__a221o_1
XANTENNA__17378__B _21340_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_17021_ _17019_/X _17021_/B vssd1 vssd1 vccd1 vccd1 _17023_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_150_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14233_ _14557_/B _15091_/C _15001_/B _14557_/A vssd1 vssd1 vccd1 vccd1 _14236_/C
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11445_ hold237/A fanout29/X _11444_/X vssd1 vssd1 vccd1 vccd1 _11445_/X sky130_fd_sc_hd__a21o_2
XANTENNA__19874__A _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_1157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14164_ _14002_/B _14004_/B _14162_/X _14163_/Y vssd1 vssd1 vccd1 vccd1 _14338_/B
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_0_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11376_ hold149/X fanout29/X _11375_/X vssd1 vssd1 vccd1 vccd1 _11376_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_46_1276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13115_ _13113_/X _13115_/B vssd1 vssd1 vccd1 vccd1 _13117_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__17394__A _17490_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15907__A _15907_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14095_ _14095_/A _14095_/B _14095_/C vssd1 vssd1 vccd1 vccd1 _14098_/A sky130_fd_sc_hd__nand3_2
X_18972_ _18972_/A _18972_/B _18972_/C vssd1 vssd1 vccd1 vccd1 _18975_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_81_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ _13046_/A _13046_/B vssd1 vssd1 vccd1 vccd1 _13047_/B sky130_fd_sc_hd__nor2_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17923_ _17923_/A _17923_/B vssd1 vssd1 vccd1 vccd1 _17943_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_147_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__14805__A_N _14806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_1030 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17854_ _18851_/C _17854_/B _19051_/C _19221_/C vssd1 vssd1 vccd1 vccd1 _17980_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_79_1063 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16805_ _16805_/A _16805_/B vssd1 vssd1 vccd1 vccd1 _16806_/C sky130_fd_sc_hd__xor2_1
X_17785_ _17785_/A _17785_/B vssd1 vssd1 vccd1 vccd1 _17805_/A sky130_fd_sc_hd__xnor2_2
X_14997_ _15373_/B _15098_/B _15368_/D _15373_/A vssd1 vssd1 vccd1 vccd1 _15001_/C
+ sky130_fd_sc_hd__a22o_1
XANTENNA__19377__B1 _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__15642__A _16031_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19524_ _19524_/A _19524_/B vssd1 vssd1 vccd1 vccd1 _19526_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_152_1117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13272__A1_N _13858_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_16736_ _16734_/X _16736_/B vssd1 vssd1 vccd1 vccd1 _16737_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_117_1237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13948_ _13948_/A _13948_/B _13948_/C _13948_/D vssd1 vssd1 vccd1 vccd1 _13948_/X
+ sky130_fd_sc_hd__or4_1
XFILLER_0_88_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19455_ _19456_/A _19456_/B vssd1 vssd1 vccd1 vccd1 _19455_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_9_1170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_16667_ _17096_/A _16860_/C _16507_/X _16508_/Y vssd1 vssd1 vccd1 vccd1 _16668_/B
+ sky130_fd_sc_hd__o2bb2a_1
X_13879_ _13878_/B _14032_/B _13878_/A vssd1 vssd1 vccd1 vccd1 _13880_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_9_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18406_ _18403_/Y _18552_/A _19008_/D _19201_/B vssd1 vssd1 vccd1 vccd1 _18552_/B
+ sky130_fd_sc_hd__and4bb_1
XFILLER_0_5_1023 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15618_ _15477_/Y _15481_/A _15616_/Y _15617_/X vssd1 vssd1 vccd1 vccd1 _15753_/A
+ sky130_fd_sc_hd__a211oi_4
XANTENNA__12216__A2 _12214_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_19386_ _19386_/A _19386_/B vssd1 vssd1 vccd1 vccd1 _19400_/A sky130_fd_sc_hd__xnor2_1
X_16598_ _16599_/A _16599_/B vssd1 vssd1 vccd1 vccd1 _17217_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_1091 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_1078 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18337_ _18789_/A _18773_/B _18338_/C _18338_/D vssd1 vssd1 vccd1 vccd1 _18339_/A
+ sky130_fd_sc_hd__a22oi_1
X_15549_ _15931_/B _16266_/C _14698_/D _15931_/A vssd1 vssd1 vccd1 vccd1 _15553_/D
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13312__D _14365_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__19487__C _20838_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_18268_ _18120_/A _18120_/B _18118_/X vssd1 vssd1 vccd1 vccd1 _18270_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_1018 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17219_ _17219_/A _17297_/A _17219_/C vssd1 vssd1 vccd1 vccd1 _17297_/B sky130_fd_sc_hd__nand3_1
X_18199_ _18197_/X _18199_/B vssd1 vssd1 vccd1 vccd1 _18200_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_142_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20230_ hold167/A fanout7/X _15356_/X _11550_/B _20229_/Y vssd1 vssd1 vccd1 vccd1
+ _20230_/X sky130_fd_sc_hd__a221o_1
Xfanout6 fanout6/A vssd1 vssd1 vccd1 vccd1 fanout6/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_12_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_20161_ _20161_/A _20161_/B vssd1 vssd1 vccd1 vccd1 _20163_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_0_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15536__B _15916_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19008__B _19185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20092_ _20235_/A _20093_/A vssd1 vssd1 vccd1 vccd1 _20240_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout297_A _21796_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_1095 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_1174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_1005 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_3608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_1196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout464_A _21753_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_1109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_1158 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_1049 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20994_ _20994_/A _20994_/B vssd1 vssd1 vccd1 vccd1 _20996_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__17918__A1 _21087_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__18285__D _19227_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout631_A _21776_/Q vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__15702__D _15702_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_1011 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_21615_ _21906_/CLK _21615_/D fanout641/X vssd1 vssd1 vccd1 vccd1 mstream_o[78] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_1210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_948 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_1119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_21546_ mstream_o[9] hold173/X _21554_/S vssd1 vssd1 vccd1 vccd1 _22073_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_63_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_1088 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__14615__B _14936_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_981 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__19694__A _19695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21477_ hold116/X sstream_i[54] _21481_/S vssd1 vssd1 vccd1 vccd1 _22004_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_133_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11230_ _21718_/D t1x[1] v2z[1] _21724_/D _11229_/X vssd1 vssd1 vccd1 vccd1 _11230_/X
+ sky130_fd_sc_hd__a221o_2
XFILLER_0_121_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20428_ _20428_/A _20428_/B vssd1 vssd1 vccd1 vccd1 _20436_/A sky130_fd_sc_hd__nand2_1
XANTENNA__18646__A2 _19866_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11161_ hold211/X fanout23/X _11160_/X vssd1 vssd1 vccd1 vccd1 _11161_/X sky130_fd_sc_hd__a21o_1
X_20359_ _20207_/X _20209_/X _20357_/Y _20358_/X vssd1 vssd1 vccd1 vccd1 _20359_/Y
+ sky130_fd_sc_hd__o211ai_4
X_11092_ _11048_/Y hold85/X _11108_/S vssd1 vssd1 vccd1 vccd1 _21686_/D sky130_fd_sc_hd__mux2_1
XANTENNA__14350__B _15788_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_1038 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_14920_ _12291_/B _14918_/Y _14919_/X vssd1 vssd1 vccd1 vccd1 _14920_/X sky130_fd_sc_hd__a21o_1
X_22029_ _22038_/CLK _22029_/D vssd1 vssd1 vccd1 vccd1 hold269/A sky130_fd_sc_hd__dfxtp_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_14851_ _14974_/A _14718_/X _14974_/B _14971_/C vssd1 vssd1 vccd1 vccd1 _14851_/X
+ sky130_fd_sc_hd__o211a_1
Xhold73 hold73/A vssd1 vssd1 vccd1 vccd1 hold73/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold84 hold84/A vssd1 vssd1 vccd1 vccd1 hold84/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_76_1258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold95 hold95/A vssd1 vssd1 vccd1 vccd1 hold95/X sky130_fd_sc_hd__dlygate4sd3_1
X_13802_ _13648_/C _13647_/Y _13800_/X _13801_/Y vssd1 vssd1 vccd1 vccd1 _13802_/Y
+ sky130_fd_sc_hd__o211ai_4
X_17570_ _17570_/A _17570_/B _17570_/C vssd1 vssd1 vccd1 vccd1 _17570_/Y sky130_fd_sc_hd__nand3_2
X_14782_ _14782_/A _14782_/B vssd1 vssd1 vccd1 vccd1 _14783_/B sky130_fd_sc_hd__and2_1
X_11994_ _11994_/A _11994_/B vssd1 vssd1 vccd1 vccd1 _11996_/B sky130_fd_sc_hd__xnor2_1
X_16521_ _17619_/A _17041_/A _16899_/B _17619_/B vssd1 vssd1 vccd1 vccd1 _16522_/C
+ sky130_fd_sc_hd__nand4_1
X_13733_ _13734_/A _13734_/B _13734_/C vssd1 vssd1 vccd1 vccd1 _13733_/X sky130_fd_sc_hd__and3_1
X_10945_ _10945_/A _10945_/B _10945_/C vssd1 vssd1 vccd1 vccd1 _10946_/B sky130_fd_sc_hd__and3_1
XFILLER_0_86_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__18773__A _20650_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__17385__A2 _20797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_19240_ _19535_/B _19240_/B _19240_/C _19387_/A vssd1 vssd1 vccd1 vccd1 _19387_/B
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_156_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_16452_ _16989_/C _17013_/D vssd1 vssd1 vccd1 vccd1 _16749_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13664_ _13664_/A _13964_/B vssd1 vssd1 vccd1 vccd1 _21364_/B sky130_fd_sc_hd__xor2_4
XANTENNA__16593__B1 _16743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10876_ hold157/A hold188/A vssd1 vssd1 vccd1 vccd1 _10878_/A sky130_fd_sc_hd__or2_1
XFILLER_0_27_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15403_ _15404_/A _15404_/B vssd1 vssd1 vccd1 vccd1 _15600_/B sky130_fd_sc_hd__or2_2
XFILLER_0_13_1231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_156_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19171_ _11550_/A _19169_/Y _19170_/X vssd1 vssd1 vccd1 vccd1 _19171_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_2_1229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12615_ _12615_/A _12615_/B vssd1 vssd1 vccd1 vccd1 _12617_/A sky130_fd_sc_hd__xnor2_2
X_16383_ _16289_/A _16289_/B _16383_/S vssd1 vssd1 vccd1 vccd1 _16384_/B sky130_fd_sc_hd__mux2_1
X_13595_ _14365_/A _15763_/A _13593_/Y _13752_/A vssd1 vssd1 vccd1 vccd1 _13597_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__18334__A1 _18787_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14806__A _14806_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__18334__B2 _18787_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13710__A _13864_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18122_ _18127_/C _18122_/B _18122_/C vssd1 vssd1 vccd1 vccd1 _18277_/A sky130_fd_sc_hd__and3_1
X_15334_ _15334_/A _15334_/B _15334_/C vssd1 vssd1 vccd1 vccd1 _15430_/B sky130_fd_sc_hd__or3_1
XANTENNA__16724__C _17526_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12546_ _12432_/X _12434_/X _12543_/X _12544_/Y vssd1 vssd1 vccd1 vccd1 _12546_/Y
+ sky130_fd_sc_hd__o211ai_4
XFILLER_0_42_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_18053_ _18185_/B _18054_/C vssd1 vssd1 vccd1 vccd1 _18055_/B sky130_fd_sc_hd__nor2_1
X_15265_ _15267_/A _15400_/B vssd1 vssd1 vccd1 vccd1 _15268_/A sky130_fd_sc_hd__or2_1
XANTENNA__16443__D _16917_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12326__A _12637_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12477_ _12373_/Y _12375_/X _12475_/Y _12476_/X vssd1 vssd1 vccd1 vccd1 _12479_/C
+ sky130_fd_sc_hd__a211oi_4
XANTENNA_4 _10792_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12906__B1 _14384_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17004_ _16956_/Y _16964_/X _17002_/A _17002_/Y vssd1 vssd1 vccd1 vccd1 _17005_/C
+ sky130_fd_sc_hd__a211oi_1
X_14216_ _15373_/B _14873_/B _14217_/D _15373_/A vssd1 vssd1 vccd1 vccd1 _14220_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11428_ _11427_/X _21283_/A _11470_/S vssd1 vssd1 vccd1 vccd1 _21814_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_123_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15196_ _15196_/A _15196_/B vssd1 vssd1 vccd1 vccd1 _15199_/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11587__D _12268_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_1062 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_686 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_14147_ _14149_/A _14149_/B _14149_/C vssd1 vssd1 vccd1 vccd1 _14301_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11359_ _11358_/X _17146_/C _11401_/S vssd1 vssd1 vccd1 vccd1 _21791_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19109__A _19430_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__21358__B _21358_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__22064__RESET_B fanout639/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11884__B _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14078_ _13921_/X _13924_/A _14076_/X _14231_/B vssd1 vssd1 vccd1 vccd1 _14078_/X
+ sky130_fd_sc_hd__o211a_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_18955_ _18955_/A _18955_/B vssd1 vssd1 vccd1 vccd1 _18975_/A sky130_fd_sc_hd__xnor2_2
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13157__A _13157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13029_ _13029_/A _13029_/B _13029_/C vssd1 vssd1 vccd1 vccd1 _13031_/A sky130_fd_sc_hd__nand3_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_17906_ _17906_/A _18026_/A _17906_/C vssd1 vssd1 vccd1 vccd1 _18026_/B sky130_fd_sc_hd__nand3_2
X_18886_ _19159_/A _18885_/B _19006_/A _18885_/D vssd1 vssd1 vccd1 vccd1 _18886_/X
+ sky130_fd_sc_hd__o22a_1
X_17837_ _17837_/A _17837_/B vssd1 vssd1 vccd1 vccd1 _17837_/X sky130_fd_sc_hd__or2_2
XFILLER_0_117_1001 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_156_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_17768_ _17768_/A _17768_/B _17768_/C vssd1 vssd1 vccd1 vccd1 _17891_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_117_1045 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15091__B _15632_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_16719_ _16718_/A _16718_/Y _16686_/X _16687_/Y vssd1 vssd1 vccd1 vccd1 _16721_/B
+ sky130_fd_sc_hd__a211o_1
X_19507_ _20462_/D _20026_/B _20733_/C _20606_/D vssd1 vssd1 vccd1 vccd1 _19661_/A
+ sky130_fd_sc_hd__nand4_2
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_17699_ _17698_/B _17698_/C _17698_/A vssd1 vssd1 vccd1 vccd1 _17700_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_117_1089 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17376__A2 fanout7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19438_ _19438_/A _19438_/B _21171_/B _21056_/B vssd1 vssd1 vccd1 vccd1 _19441_/B
+ sky130_fd_sc_hd__nand4_1
XFILLER_0_119_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_1077 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_1197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19369_ _19370_/A _19370_/B vssd1 vssd1 vccd1 vccd1 _19483_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_128_961 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_1129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__14716__A _14716_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__17128__A2 _17146_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_21400_ _21420_/S _20377_/B _21381_/B _21399_/Y vssd1 vssd1 vccd1 vccd1 _21400_/X
+ sky130_fd_sc_hd__a211o_1
XANTENNA__13620__A _14713_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__20132__A1 _20416_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__20132__B2 _20416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13977__D _16409_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21331_ _21349_/A _21331_/B vssd1 vssd1 vccd1 vccd1 _21331_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_981 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout212_A _21283_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11778__C _13017_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_1141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_1005 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21262_ _21218_/A _21217_/B _21215_/Y vssd1 vssd1 vccd1 vccd1 _21263_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_4_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_1185 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_973 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__19664__D _20606_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13570__B1 _14365_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_20213_ _20066_/A _20066_/B _20024_/A vssd1 vssd1 vccd1 vccd1 _20215_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_1049 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__17836__B1 fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_1124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_1173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_21193_ _21193_/A _21193_/B vssd1 vssd1 vccd1 vccd1 _21195_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_40_483 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_1037 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_20144_ _19874_/B _19967_/X _19970_/A _19970_/B vssd1 vssd1 vccd1 vccd1 _20151_/A
+ sky130_fd_sc_hd__o2bb2a_1
XANTENNA_fanout581_A _12269_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__17762__A _18030_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_20075_ _20075_/A _20075_/B vssd1 vssd1 vccd1 vccd1 _20078_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__13873__A1 _14195_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__18800__A2 _20249_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_3427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1101 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_1093 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_3438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_3449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12428__A2 _14698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_135_1145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13514__B _21361_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_20977_ _21095_/A _20978_/C _20978_/A vssd1 vssd1 vccd1 vccd1 _20979_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_71_1133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_1009 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15432__D _15954_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_1189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13233__C _14155_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__19201__B _19201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12400_ _12511_/A _12402_/A _12858_/C _12991_/D _12305_/B vssd1 vssd1 vccd1 vccd1
+ _12410_/A sky130_fd_sc_hd__a41o_1
X_13380_ _13381_/C _16328_/B _13378_/Y _13527_/A vssd1 vssd1 vccd1 vccd1 _13382_/A
+ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_24_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_929 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__16878__A1 _16989_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ _12332_/B _12332_/A vssd1 vssd1 vccd1 vccd1 _12331_/X sky130_fd_sc_hd__and2b_1
X_21529_ hold299/X sstream_i[106] _21536_/S vssd1 vssd1 vccd1 vccd1 _22056_/D sky130_fd_sc_hd__mux2_1
XFILLER_0_90_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_1241 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11688__C _12420_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_15050_ _15013_/X _15014_/Y _15050_/C _15050_/D vssd1 vssd1 vccd1 vccd1 _15050_/X
+ sky130_fd_sc_hd__and4bb_1
X_12262_ _12261_/A _12268_/B _21727_/Q _12269_/B vssd1 vssd1 vccd1 vccd1 _12262_/X
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_1105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__16560__B _16743_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11167__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11213_ _14557_/D _11212_/X _11284_/S vssd1 vssd1 vccd1 vccd1 _21754_/D sky130_fd_sc_hd__mux2_1
X_14001_ _14000_/B _14153_/B _14000_/A vssd1 vssd1 vccd1 vccd1 _14002_/C sky130_fd_sc_hd__a21o_1
XANTENNA__14999__C _15098_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_995 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_1149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12193_ _12193_/A _12193_/B _12193_/C vssd1 vssd1 vccd1 vccd1 _12228_/A sky130_fd_sc_hd__nand3_1
XANTENNA__15302__A1 _15439_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11144_ _12512_/A _11143_/X _11260_/S vssd1 vssd1 vccd1 vccd1 _21731_/D sky130_fd_sc_hd__mux2_1
XANTENNA__19871__B _20394_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__15891__S fanout2/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_18740_ _20317_/D _19382_/B _18741_/C _18741_/D vssd1 vssd1 vccd1 vccd1 _18740_/X
+ sky130_fd_sc_hd__and4_1
X_15952_ _15867_/B _15952_/B vssd1 vssd1 vccd1 vccd1 _15996_/A sky130_fd_sc_hd__nand2b_1
X_11075_ _10903_/Y hold70/X _11088_/S vssd1 vssd1 vccd1 vccd1 _21670_/D sky130_fd_sc_hd__mux2_1
XANTENNA__13408__C _14354_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_14903_ _14904_/A _14904_/B vssd1 vssd1 vccd1 vccd1 _15067_/A sky130_fd_sc_hd__or2_1
X_18671_ _18516_/C _18515_/Y _18669_/X _18670_/Y vssd1 vssd1 vccd1 vccd1 _18674_/C
+ sky130_fd_sc_hd__o211a_2
X_15883_ _16011_/A _15881_/X _15708_/Y _15711_/Y vssd1 vssd1 vccd1 vccd1 _15883_/X
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_1044 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_1201 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__15192__A _15192_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_17622_ _17621_/C _17741_/B _17737_/A _17620_/Y vssd1 vssd1 vccd1 vccd1 _17622_/X
+ sky130_fd_sc_hd__o2bb2a_1
X_14834_ _14833_/B _14833_/C _14833_/A vssd1 vssd1 vccd1 vccd1 _14836_/B sky130_fd_sc_hd__a21o_1
XANTENNA__13705__A _13858_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_1028 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_1245 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17553_ _17551_/Y _17552_/X _17657_/A _19439_/A vssd1 vssd1 vccd1 vccd1 _17555_/A
+ sky130_fd_sc_hd__and4bb_1
X_14765_ _14650_/A _14650_/B _14648_/Y vssd1 vssd1 vccd1 vccd1 _14808_/A sky130_fd_sc_hd__o21ba_1
XFILLER_0_98_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11977_ _11977_/A _11979_/A _11976_/A vssd1 vssd1 vccd1 vccd1 _11977_/X sky130_fd_sc_hd__or3b_1
XFILLER_0_86_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_16504_ _17197_/A _16503_/C _16503_/A vssd1 vssd1 vccd1 vccd1 _16505_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__15369__A1 _16027_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13716_ _13716_/A _13716_/B vssd1 vssd1 vccd1 vccd1 _13718_/B sky130_fd_sc_hd__xnor2_1
X_10928_ hold109/A hold158/A vssd1 vssd1 vccd1 vccd1 _10931_/A sky130_fd_sc_hd__or2_1
XFILLER_0_6_1140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_17484_ _17594_/A _17484_/B vssd1 vssd1 vccd1 vccd1 _17484_/X sky130_fd_sc_hd__and2_4
X_14696_ _14696_/A _14696_/B vssd1 vssd1 vccd1 vccd1 _14705_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_74_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_156_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_19223_ _20026_/B _19223_/B vssd1 vssd1 vccd1 vccd1 _19224_/B sky130_fd_sc_hd__nand2_1
X_16435_ _16435_/A _16435_/B vssd1 vssd1 vccd1 vccd1 _16436_/B sky130_fd_sc_hd__xnor2_2
XFILLER_0_117_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__16627__A1_N _16870_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13647_ _13648_/A _13648_/B _13648_/C _13648_/D vssd1 vssd1 vccd1 vccd1 _13647_/Y
+ sky130_fd_sc_hd__nor4_2
XANTENNA__19111__B _19866_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10859_ _10859_/A _10859_/B _10859_/C vssd1 vssd1 vccd1 vccd1 _10860_/B sky130_fd_sc_hd__and3_1
XFILLER_0_6_1195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_1026 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_1050 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__18008__A _18008_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13440__A _14367_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_1061 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_1048 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_19154_ _19154_/A _19154_/B vssd1 vssd1 vccd1 vccd1 _19157_/A sky130_fd_sc_hd__or2_1
X_16366_ _16360_/A _16366_/B vssd1 vssd1 vccd1 vccd1 _16366_/X sky130_fd_sc_hd__and2b_1
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_43_clk_i _21822_/CLK vssd1 vssd1 vccd1 vccd1 _21724_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13578_ _13578_/A _13578_/B vssd1 vssd1 vccd1 vccd1 _13580_/C sky130_fd_sc_hd__xnor2_2
XANTENNA__18858__A2 _21261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_953 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_18105_ _17850_/A _17850_/B _17990_/B _17988_/Y vssd1 vssd1 vccd1 vccd1 _18106_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__16869__A1 _17013_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_1113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_15317_ _16092_/D _15788_/B _15115_/C _15113_/A vssd1 vssd1 vccd1 vccd1 _15324_/A
+ sky130_fd_sc_hd__a31oi_4
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_1173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_19085_ _18955_/A _18954_/B _18952_/X vssd1 vssd1 vccd1 vccd1 _19101_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_42_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12529_ _12750_/A _13152_/C _13152_/D _12528_/B vssd1 vssd1 vccd1 vccd1 _12530_/D
+ sky130_fd_sc_hd__a22o_1
X_16297_ _16297_/A _16297_/B vssd1 vssd1 vccd1 vccd1 _16298_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__17530__A2 _17206_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_923 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_18036_ _19892_/A _18624_/A _18175_/A _18035_/D vssd1 vssd1 vccd1 vccd1 _18038_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_951 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_15248_ _15249_/A _15249_/B vssd1 vssd1 vccd1 vccd1 _15248_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_300 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_258 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__16470__B _17520_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11158__A2 fanout23/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_15179_ _15179_/A _15179_/B _15179_/C vssd1 vssd1 vccd1 vccd1 _15179_/X sky130_fd_sc_hd__and3_1
XFILLER_0_111_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout308 _17123_/C vssd1 vssd1 vccd1 vccd1 _17124_/C sky130_fd_sc_hd__buf_4
Xfanout319 _17493_/A vssd1 vssd1 vccd1 vccd1 _17277_/A sky130_fd_sc_hd__buf_4
X_19987_ _21199_/A fanout96/X _20265_/D _20838_/B vssd1 vssd1 vccd1 vccd1 _19987_/X
+ sky130_fd_sc_hd__a22o_1
X_18938_ _18938_/A _18938_/B _18938_/C vssd1 vssd1 vccd1 vccd1 _19084_/A sky130_fd_sc_hd__nand3_1
.ends

