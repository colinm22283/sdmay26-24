VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vga
  CLASS BLOCK ;
  FOREIGN vga ;
  ORIGIN 0.000 0.000 ;
  SIZE 600.000 BY 600.000 ;
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 149.590 596.000 149.870 600.000 ;
    END
  END clk_i
  PIN enable_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 469.240 600.000 469.840 ;
    END
  END enable_i
  PIN fb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 591.640 600.000 592.240 ;
    END
  END fb_i
  PIN hsync_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END hsync_o
  PIN mport_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 6.840 600.000 7.440 ;
    END
  END mport_i[0]
  PIN mport_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 142.840 600.000 143.440 ;
    END
  END mport_i[10]
  PIN mport_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 156.440 600.000 157.040 ;
    END
  END mport_i[11]
  PIN mport_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 170.040 600.000 170.640 ;
    END
  END mport_i[12]
  PIN mport_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 183.640 600.000 184.240 ;
    END
  END mport_i[13]
  PIN mport_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 197.240 600.000 197.840 ;
    END
  END mport_i[14]
  PIN mport_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 210.840 600.000 211.440 ;
    END
  END mport_i[15]
  PIN mport_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 224.440 600.000 225.040 ;
    END
  END mport_i[16]
  PIN mport_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 238.040 600.000 238.640 ;
    END
  END mport_i[17]
  PIN mport_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 251.640 600.000 252.240 ;
    END
  END mport_i[18]
  PIN mport_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 265.240 600.000 265.840 ;
    END
  END mport_i[19]
  PIN mport_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 20.440 600.000 21.040 ;
    END
  END mport_i[1]
  PIN mport_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 278.840 600.000 279.440 ;
    END
  END mport_i[20]
  PIN mport_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 292.440 600.000 293.040 ;
    END
  END mport_i[21]
  PIN mport_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 306.040 600.000 306.640 ;
    END
  END mport_i[22]
  PIN mport_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 319.640 600.000 320.240 ;
    END
  END mport_i[23]
  PIN mport_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 333.240 600.000 333.840 ;
    END
  END mport_i[24]
  PIN mport_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 346.840 600.000 347.440 ;
    END
  END mport_i[25]
  PIN mport_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 360.440 600.000 361.040 ;
    END
  END mport_i[26]
  PIN mport_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 374.040 600.000 374.640 ;
    END
  END mport_i[27]
  PIN mport_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 387.640 600.000 388.240 ;
    END
  END mport_i[28]
  PIN mport_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 401.240 600.000 401.840 ;
    END
  END mport_i[29]
  PIN mport_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 34.040 600.000 34.640 ;
    END
  END mport_i[2]
  PIN mport_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 414.840 600.000 415.440 ;
    END
  END mport_i[30]
  PIN mport_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 428.440 600.000 429.040 ;
    END
  END mport_i[31]
  PIN mport_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 442.040 600.000 442.640 ;
    END
  END mport_i[32]
  PIN mport_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 455.640 600.000 456.240 ;
    END
  END mport_i[33]
  PIN mport_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 47.640 600.000 48.240 ;
    END
  END mport_i[3]
  PIN mport_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 61.240 600.000 61.840 ;
    END
  END mport_i[4]
  PIN mport_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 74.840 600.000 75.440 ;
    END
  END mport_i[5]
  PIN mport_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 88.440 600.000 89.040 ;
    END
  END mport_i[6]
  PIN mport_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 102.040 600.000 102.640 ;
    END
  END mport_i[7]
  PIN mport_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 596.000 115.640 600.000 116.240 ;
    END
  END mport_i[8]
  PIN mport_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 129.240 600.000 129.840 ;
    END
  END mport_i[9]
  PIN mport_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END mport_o[0]
  PIN mport_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END mport_o[10]
  PIN mport_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END mport_o[11]
  PIN mport_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END mport_o[12]
  PIN mport_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END mport_o[13]
  PIN mport_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END mport_o[14]
  PIN mport_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END mport_o[15]
  PIN mport_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END mport_o[16]
  PIN mport_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END mport_o[17]
  PIN mport_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END mport_o[18]
  PIN mport_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END mport_o[19]
  PIN mport_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END mport_o[1]
  PIN mport_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END mport_o[20]
  PIN mport_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END mport_o[21]
  PIN mport_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 201.320 4.000 201.920 ;
    END
  END mport_o[22]
  PIN mport_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END mport_o[23]
  PIN mport_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END mport_o[24]
  PIN mport_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END mport_o[25]
  PIN mport_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.960 4.000 234.560 ;
    END
  END mport_o[26]
  PIN mport_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END mport_o[27]
  PIN mport_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 250.280 4.000 250.880 ;
    END
  END mport_o[28]
  PIN mport_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END mport_o[29]
  PIN mport_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END mport_o[2]
  PIN mport_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 266.600 4.000 267.200 ;
    END
  END mport_o[30]
  PIN mport_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END mport_o[31]
  PIN mport_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END mport_o[32]
  PIN mport_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END mport_o[33]
  PIN mport_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END mport_o[34]
  PIN mport_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END mport_o[35]
  PIN mport_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END mport_o[36]
  PIN mport_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END mport_o[37]
  PIN mport_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END mport_o[38]
  PIN mport_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END mport_o[39]
  PIN mport_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END mport_o[3]
  PIN mport_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.200 4.000 348.800 ;
    END
  END mport_o[40]
  PIN mport_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END mport_o[41]
  PIN mport_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END mport_o[42]
  PIN mport_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 372.680 4.000 373.280 ;
    END
  END mport_o[43]
  PIN mport_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END mport_o[44]
  PIN mport_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END mport_o[45]
  PIN mport_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.160 4.000 397.760 ;
    END
  END mport_o[46]
  PIN mport_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END mport_o[47]
  PIN mport_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 413.480 4.000 414.080 ;
    END
  END mport_o[48]
  PIN mport_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END mport_o[49]
  PIN mport_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END mport_o[4]
  PIN mport_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END mport_o[50]
  PIN mport_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.960 4.000 438.560 ;
    END
  END mport_o[51]
  PIN mport_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END mport_o[52]
  PIN mport_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END mport_o[53]
  PIN mport_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END mport_o[54]
  PIN mport_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 470.600 4.000 471.200 ;
    END
  END mport_o[55]
  PIN mport_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END mport_o[56]
  PIN mport_o[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END mport_o[57]
  PIN mport_o[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END mport_o[58]
  PIN mport_o[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END mport_o[59]
  PIN mport_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END mport_o[5]
  PIN mport_o[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END mport_o[60]
  PIN mport_o[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 519.560 4.000 520.160 ;
    END
  END mport_o[61]
  PIN mport_o[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END mport_o[62]
  PIN mport_o[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END mport_o[63]
  PIN mport_o[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 544.040 4.000 544.640 ;
    END
  END mport_o[64]
  PIN mport_o[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END mport_o[65]
  PIN mport_o[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 560.360 4.000 560.960 ;
    END
  END mport_o[66]
  PIN mport_o[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 568.520 4.000 569.120 ;
    END
  END mport_o[67]
  PIN mport_o[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.680 4.000 577.280 ;
    END
  END mport_o[68]
  PIN mport_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END mport_o[6]
  PIN mport_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.920 4.000 79.520 ;
    END
  END mport_o[7]
  PIN mport_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END mport_o[8]
  PIN mport_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END mport_o[9]
  PIN nrst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 449.510 596.000 449.790 600.000 ;
    END
  END nrst_i
  PIN pixel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END pixel_o[0]
  PIN pixel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END pixel_o[1]
  PIN pixel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END pixel_o[2]
  PIN pixel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END pixel_o[3]
  PIN pixel_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END pixel_o[4]
  PIN pixel_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END pixel_o[5]
  PIN pixel_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END pixel_o[6]
  PIN pixel_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END pixel_o[7]
  PIN prescaler_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 482.840 600.000 483.440 ;
    END
  END prescaler_i[0]
  PIN prescaler_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 496.440 600.000 497.040 ;
    END
  END prescaler_i[1]
  PIN prescaler_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 510.040 600.000 510.640 ;
    END
  END prescaler_i[2]
  PIN prescaler_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 596.000 523.640 600.000 524.240 ;
    END
  END prescaler_i[3]
  PIN resolution_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 537.240 600.000 537.840 ;
    END
  END resolution_i[0]
  PIN resolution_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 550.840 600.000 551.440 ;
    END
  END resolution_i[1]
  PIN resolution_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 564.440 600.000 565.040 ;
    END
  END resolution_i[2]
  PIN resolution_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 596.000 578.040 600.000 578.640 ;
    END
  END resolution_i[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN vsync_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END vsync_o
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 594.320 587.605 ;
      LAYER met1 ;
        RECT 4.670 9.220 597.930 588.160 ;
      LAYER met2 ;
        RECT 4.690 595.720 149.310 596.000 ;
        RECT 150.150 595.720 449.230 596.000 ;
        RECT 450.070 595.720 597.900 596.000 ;
        RECT 4.690 4.280 597.900 595.720 ;
        RECT 4.690 3.670 30.170 4.280 ;
        RECT 31.010 3.670 89.970 4.280 ;
        RECT 90.810 3.670 149.770 4.280 ;
        RECT 150.610 3.670 209.570 4.280 ;
        RECT 210.410 3.670 269.370 4.280 ;
        RECT 270.210 3.670 329.170 4.280 ;
        RECT 330.010 3.670 388.970 4.280 ;
        RECT 389.810 3.670 448.770 4.280 ;
        RECT 449.610 3.670 508.570 4.280 ;
        RECT 509.410 3.670 568.370 4.280 ;
        RECT 569.210 3.670 597.900 4.280 ;
      LAYER met3 ;
        RECT 3.990 579.040 596.095 587.685 ;
        RECT 3.990 577.680 595.600 579.040 ;
        RECT 4.400 577.640 595.600 577.680 ;
        RECT 4.400 576.280 596.095 577.640 ;
        RECT 3.990 569.520 596.095 576.280 ;
        RECT 4.400 568.120 596.095 569.520 ;
        RECT 3.990 565.440 596.095 568.120 ;
        RECT 3.990 564.040 595.600 565.440 ;
        RECT 3.990 561.360 596.095 564.040 ;
        RECT 4.400 559.960 596.095 561.360 ;
        RECT 3.990 553.200 596.095 559.960 ;
        RECT 4.400 551.840 596.095 553.200 ;
        RECT 4.400 551.800 595.600 551.840 ;
        RECT 3.990 550.440 595.600 551.800 ;
        RECT 3.990 545.040 596.095 550.440 ;
        RECT 4.400 543.640 596.095 545.040 ;
        RECT 3.990 538.240 596.095 543.640 ;
        RECT 3.990 536.880 595.600 538.240 ;
        RECT 4.400 536.840 595.600 536.880 ;
        RECT 4.400 535.480 596.095 536.840 ;
        RECT 3.990 528.720 596.095 535.480 ;
        RECT 4.400 527.320 596.095 528.720 ;
        RECT 3.990 524.640 596.095 527.320 ;
        RECT 3.990 523.240 595.600 524.640 ;
        RECT 3.990 520.560 596.095 523.240 ;
        RECT 4.400 519.160 596.095 520.560 ;
        RECT 3.990 512.400 596.095 519.160 ;
        RECT 4.400 511.040 596.095 512.400 ;
        RECT 4.400 511.000 595.600 511.040 ;
        RECT 3.990 509.640 595.600 511.000 ;
        RECT 3.990 504.240 596.095 509.640 ;
        RECT 4.400 502.840 596.095 504.240 ;
        RECT 3.990 497.440 596.095 502.840 ;
        RECT 3.990 496.080 595.600 497.440 ;
        RECT 4.400 496.040 595.600 496.080 ;
        RECT 4.400 494.680 596.095 496.040 ;
        RECT 3.990 487.920 596.095 494.680 ;
        RECT 4.400 486.520 596.095 487.920 ;
        RECT 3.990 483.840 596.095 486.520 ;
        RECT 3.990 482.440 595.600 483.840 ;
        RECT 3.990 479.760 596.095 482.440 ;
        RECT 4.400 478.360 596.095 479.760 ;
        RECT 3.990 471.600 596.095 478.360 ;
        RECT 4.400 470.240 596.095 471.600 ;
        RECT 4.400 470.200 595.600 470.240 ;
        RECT 3.990 468.840 595.600 470.200 ;
        RECT 3.990 463.440 596.095 468.840 ;
        RECT 4.400 462.040 596.095 463.440 ;
        RECT 3.990 456.640 596.095 462.040 ;
        RECT 3.990 455.280 595.600 456.640 ;
        RECT 4.400 455.240 595.600 455.280 ;
        RECT 4.400 453.880 596.095 455.240 ;
        RECT 3.990 447.120 596.095 453.880 ;
        RECT 4.400 445.720 596.095 447.120 ;
        RECT 3.990 443.040 596.095 445.720 ;
        RECT 3.990 441.640 595.600 443.040 ;
        RECT 3.990 438.960 596.095 441.640 ;
        RECT 4.400 437.560 596.095 438.960 ;
        RECT 3.990 430.800 596.095 437.560 ;
        RECT 4.400 429.440 596.095 430.800 ;
        RECT 4.400 429.400 595.600 429.440 ;
        RECT 3.990 428.040 595.600 429.400 ;
        RECT 3.990 422.640 596.095 428.040 ;
        RECT 4.400 421.240 596.095 422.640 ;
        RECT 3.990 415.840 596.095 421.240 ;
        RECT 3.990 414.480 595.600 415.840 ;
        RECT 4.400 414.440 595.600 414.480 ;
        RECT 4.400 413.080 596.095 414.440 ;
        RECT 3.990 406.320 596.095 413.080 ;
        RECT 4.400 404.920 596.095 406.320 ;
        RECT 3.990 402.240 596.095 404.920 ;
        RECT 3.990 400.840 595.600 402.240 ;
        RECT 3.990 398.160 596.095 400.840 ;
        RECT 4.400 396.760 596.095 398.160 ;
        RECT 3.990 390.000 596.095 396.760 ;
        RECT 4.400 388.640 596.095 390.000 ;
        RECT 4.400 388.600 595.600 388.640 ;
        RECT 3.990 387.240 595.600 388.600 ;
        RECT 3.990 381.840 596.095 387.240 ;
        RECT 4.400 380.440 596.095 381.840 ;
        RECT 3.990 375.040 596.095 380.440 ;
        RECT 3.990 373.680 595.600 375.040 ;
        RECT 4.400 373.640 595.600 373.680 ;
        RECT 4.400 372.280 596.095 373.640 ;
        RECT 3.990 365.520 596.095 372.280 ;
        RECT 4.400 364.120 596.095 365.520 ;
        RECT 3.990 361.440 596.095 364.120 ;
        RECT 3.990 360.040 595.600 361.440 ;
        RECT 3.990 357.360 596.095 360.040 ;
        RECT 4.400 355.960 596.095 357.360 ;
        RECT 3.990 349.200 596.095 355.960 ;
        RECT 4.400 347.840 596.095 349.200 ;
        RECT 4.400 347.800 595.600 347.840 ;
        RECT 3.990 346.440 595.600 347.800 ;
        RECT 3.990 341.040 596.095 346.440 ;
        RECT 4.400 339.640 596.095 341.040 ;
        RECT 3.990 334.240 596.095 339.640 ;
        RECT 3.990 332.880 595.600 334.240 ;
        RECT 4.400 332.840 595.600 332.880 ;
        RECT 4.400 331.480 596.095 332.840 ;
        RECT 3.990 324.720 596.095 331.480 ;
        RECT 4.400 323.320 596.095 324.720 ;
        RECT 3.990 320.640 596.095 323.320 ;
        RECT 3.990 319.240 595.600 320.640 ;
        RECT 3.990 316.560 596.095 319.240 ;
        RECT 4.400 315.160 596.095 316.560 ;
        RECT 3.990 308.400 596.095 315.160 ;
        RECT 4.400 307.040 596.095 308.400 ;
        RECT 4.400 307.000 595.600 307.040 ;
        RECT 3.990 305.640 595.600 307.000 ;
        RECT 3.990 300.240 596.095 305.640 ;
        RECT 4.400 298.840 596.095 300.240 ;
        RECT 3.990 293.440 596.095 298.840 ;
        RECT 3.990 292.080 595.600 293.440 ;
        RECT 4.400 292.040 595.600 292.080 ;
        RECT 4.400 290.680 596.095 292.040 ;
        RECT 3.990 283.920 596.095 290.680 ;
        RECT 4.400 282.520 596.095 283.920 ;
        RECT 3.990 279.840 596.095 282.520 ;
        RECT 3.990 278.440 595.600 279.840 ;
        RECT 3.990 275.760 596.095 278.440 ;
        RECT 4.400 274.360 596.095 275.760 ;
        RECT 3.990 267.600 596.095 274.360 ;
        RECT 4.400 266.240 596.095 267.600 ;
        RECT 4.400 266.200 595.600 266.240 ;
        RECT 3.990 264.840 595.600 266.200 ;
        RECT 3.990 259.440 596.095 264.840 ;
        RECT 4.400 258.040 596.095 259.440 ;
        RECT 3.990 252.640 596.095 258.040 ;
        RECT 3.990 251.280 595.600 252.640 ;
        RECT 4.400 251.240 595.600 251.280 ;
        RECT 4.400 249.880 596.095 251.240 ;
        RECT 3.990 243.120 596.095 249.880 ;
        RECT 4.400 241.720 596.095 243.120 ;
        RECT 3.990 239.040 596.095 241.720 ;
        RECT 3.990 237.640 595.600 239.040 ;
        RECT 3.990 234.960 596.095 237.640 ;
        RECT 4.400 233.560 596.095 234.960 ;
        RECT 3.990 226.800 596.095 233.560 ;
        RECT 4.400 225.440 596.095 226.800 ;
        RECT 4.400 225.400 595.600 225.440 ;
        RECT 3.990 224.040 595.600 225.400 ;
        RECT 3.990 218.640 596.095 224.040 ;
        RECT 4.400 217.240 596.095 218.640 ;
        RECT 3.990 211.840 596.095 217.240 ;
        RECT 3.990 210.480 595.600 211.840 ;
        RECT 4.400 210.440 595.600 210.480 ;
        RECT 4.400 209.080 596.095 210.440 ;
        RECT 3.990 202.320 596.095 209.080 ;
        RECT 4.400 200.920 596.095 202.320 ;
        RECT 3.990 198.240 596.095 200.920 ;
        RECT 3.990 196.840 595.600 198.240 ;
        RECT 3.990 194.160 596.095 196.840 ;
        RECT 4.400 192.760 596.095 194.160 ;
        RECT 3.990 186.000 596.095 192.760 ;
        RECT 4.400 184.640 596.095 186.000 ;
        RECT 4.400 184.600 595.600 184.640 ;
        RECT 3.990 183.240 595.600 184.600 ;
        RECT 3.990 177.840 596.095 183.240 ;
        RECT 4.400 176.440 596.095 177.840 ;
        RECT 3.990 171.040 596.095 176.440 ;
        RECT 3.990 169.680 595.600 171.040 ;
        RECT 4.400 169.640 595.600 169.680 ;
        RECT 4.400 168.280 596.095 169.640 ;
        RECT 3.990 161.520 596.095 168.280 ;
        RECT 4.400 160.120 596.095 161.520 ;
        RECT 3.990 157.440 596.095 160.120 ;
        RECT 3.990 156.040 595.600 157.440 ;
        RECT 3.990 153.360 596.095 156.040 ;
        RECT 4.400 151.960 596.095 153.360 ;
        RECT 3.990 145.200 596.095 151.960 ;
        RECT 4.400 143.840 596.095 145.200 ;
        RECT 4.400 143.800 595.600 143.840 ;
        RECT 3.990 142.440 595.600 143.800 ;
        RECT 3.990 137.040 596.095 142.440 ;
        RECT 4.400 135.640 596.095 137.040 ;
        RECT 3.990 130.240 596.095 135.640 ;
        RECT 3.990 128.880 595.600 130.240 ;
        RECT 4.400 128.840 595.600 128.880 ;
        RECT 4.400 127.480 596.095 128.840 ;
        RECT 3.990 120.720 596.095 127.480 ;
        RECT 4.400 119.320 596.095 120.720 ;
        RECT 3.990 116.640 596.095 119.320 ;
        RECT 3.990 115.240 595.600 116.640 ;
        RECT 3.990 112.560 596.095 115.240 ;
        RECT 4.400 111.160 596.095 112.560 ;
        RECT 3.990 104.400 596.095 111.160 ;
        RECT 4.400 103.040 596.095 104.400 ;
        RECT 4.400 103.000 595.600 103.040 ;
        RECT 3.990 101.640 595.600 103.000 ;
        RECT 3.990 96.240 596.095 101.640 ;
        RECT 4.400 94.840 596.095 96.240 ;
        RECT 3.990 89.440 596.095 94.840 ;
        RECT 3.990 88.080 595.600 89.440 ;
        RECT 4.400 88.040 595.600 88.080 ;
        RECT 4.400 86.680 596.095 88.040 ;
        RECT 3.990 79.920 596.095 86.680 ;
        RECT 4.400 78.520 596.095 79.920 ;
        RECT 3.990 75.840 596.095 78.520 ;
        RECT 3.990 74.440 595.600 75.840 ;
        RECT 3.990 71.760 596.095 74.440 ;
        RECT 4.400 70.360 596.095 71.760 ;
        RECT 3.990 63.600 596.095 70.360 ;
        RECT 4.400 62.240 596.095 63.600 ;
        RECT 4.400 62.200 595.600 62.240 ;
        RECT 3.990 60.840 595.600 62.200 ;
        RECT 3.990 55.440 596.095 60.840 ;
        RECT 4.400 54.040 596.095 55.440 ;
        RECT 3.990 48.640 596.095 54.040 ;
        RECT 3.990 47.280 595.600 48.640 ;
        RECT 4.400 47.240 595.600 47.280 ;
        RECT 4.400 45.880 596.095 47.240 ;
        RECT 3.990 39.120 596.095 45.880 ;
        RECT 4.400 37.720 596.095 39.120 ;
        RECT 3.990 35.040 596.095 37.720 ;
        RECT 3.990 33.640 595.600 35.040 ;
        RECT 3.990 30.960 596.095 33.640 ;
        RECT 4.400 29.560 596.095 30.960 ;
        RECT 3.990 22.800 596.095 29.560 ;
        RECT 4.400 21.440 596.095 22.800 ;
        RECT 4.400 21.400 595.600 21.440 ;
        RECT 3.990 20.040 595.600 21.400 ;
        RECT 3.990 7.840 596.095 20.040 ;
        RECT 3.990 6.975 595.600 7.840 ;
      LAYER met4 ;
        RECT 15.935 15.135 20.640 585.985 ;
        RECT 23.040 15.135 97.440 585.985 ;
        RECT 99.840 15.135 174.240 585.985 ;
        RECT 176.640 15.135 251.040 585.985 ;
        RECT 253.440 15.135 327.840 585.985 ;
        RECT 330.240 15.135 404.640 585.985 ;
        RECT 407.040 15.135 481.440 585.985 ;
        RECT 483.840 15.135 558.240 585.985 ;
        RECT 560.640 15.135 585.745 585.985 ;
  END
END vga
END LIBRARY

