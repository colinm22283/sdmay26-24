* NGSPICE file created from mac.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

.subckt mac a_i[0] a_i[10] a_i[11] a_i[12] a_i[13] a_i[14] a_i[15] a_i[16] a_i[17]
+ a_i[18] a_i[19] a_i[1] a_i[20] a_i[21] a_i[22] a_i[23] a_i[24] a_i[25] a_i[26] a_i[27]
+ a_i[28] a_i[29] a_i[2] a_i[30] a_i[31] a_i[3] a_i[4] a_i[5] a_i[6] a_i[7] a_i[8]
+ a_i[9] b_i[0] b_i[10] b_i[11] b_i[12] b_i[13] b_i[14] b_i[15] b_i[16] b_i[17] b_i[18]
+ b_i[19] b_i[1] b_i[20] b_i[21] b_i[22] b_i[23] b_i[24] b_i[25] b_i[26] b_i[27] b_i[28]
+ b_i[29] b_i[2] b_i[30] b_i[31] b_i[3] b_i[4] b_i[5] b_i[6] b_i[7] b_i[8] b_i[9]
+ clk nrst vccd1 vssd1 y_o[0] y_o[10] y_o[11] y_o[12] y_o[13] y_o[14] y_o[15] y_o[16]
+ y_o[17] y_o[18] y_o[19] y_o[1] y_o[20] y_o[21] y_o[22] y_o[23] y_o[24] y_o[25] y_o[26]
+ y_o[27] y_o[28] y_o[29] y_o[2] y_o[30] y_o[31] y_o[3] y_o[4] y_o[5] y_o[6] y_o[7]
+ y_o[8] y_o[9]
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05903_ _08574_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _05906_/B sky130_fd_sc_hd__nand2_1
X_09671_ _09673_/A vssd1 vssd1 vccd1 vccd1 _09672_/B sky130_fd_sc_hd__inv_2
X_06883_ _06884_/B _06884_/A vssd1 vssd1 vccd1 vccd1 _06883_/Y sky130_fd_sc_hd__nand2_1
X_08622_ _08622_/A vssd1 vssd1 vccd1 vccd1 _08623_/C sky130_fd_sc_hd__inv_2
X_05834_ _05836_/C vssd1 vssd1 vccd1 vccd1 _05835_/B sky130_fd_sc_hd__inv_2
X_05765_ _05855_/A _05854_/A vssd1 vssd1 vccd1 vccd1 _05765_/Y sky130_fd_sc_hd__nand2_1
X_08553_ _08562_/B vssd1 vssd1 vccd1 vccd1 _08554_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07504_ _07504_/A _07504_/B vssd1 vssd1 vccd1 vccd1 _07614_/B sky130_fd_sc_hd__nand2_1
X_08484_ _08485_/A _08485_/B vssd1 vssd1 vccd1 vccd1 _08486_/A sky130_fd_sc_hd__or2_1
XFILLER_0_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07435_ _07436_/B _07435_/B _07435_/C vssd1 vssd1 vccd1 vccd1 _07713_/B sky130_fd_sc_hd__nand3_1
X_05696_ _05696_/A _05696_/B vssd1 vssd1 vccd1 vccd1 _05697_/A sky130_fd_sc_hd__nand2_1
X_07366_ _07453_/B _07452_/A _07452_/B vssd1 vssd1 vccd1 vccd1 _07545_/B sky130_fd_sc_hd__nand3b_2
X_09105_ _09105_/A _09105_/B vssd1 vssd1 vccd1 vccd1 _09105_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_72_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07297_ _07297_/A _07297_/B vssd1 vssd1 vccd1 vccd1 _07301_/A sky130_fd_sc_hd__nand2_1
X_06317_ _06317_/A _06317_/B vssd1 vssd1 vccd1 vccd1 _06688_/B sky130_fd_sc_hd__nand2_1
X_09036_ _09036_/A _09036_/B _09036_/C vssd1 vssd1 vccd1 vccd1 _09037_/B sky130_fd_sc_hd__nand3_1
X_06248_ _06248_/A _06248_/B _06248_/C vssd1 vssd1 vccd1 vccd1 _06413_/C sky130_fd_sc_hd__nand3_1
X_06179_ _06299_/A _06179_/B _06179_/C vssd1 vssd1 vccd1 vccd1 _06221_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_40_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09938_ _09936_/Y _09938_/B _09938_/C vssd1 vssd1 vccd1 vccd1 _09939_/B sky130_fd_sc_hd__nand3b_1
X_09869_ _10305_/B _09869_/B vssd1 vssd1 vccd1 vccd1 _09893_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07523__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_67_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10713_ _10718_/CLK _10713_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold58/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10644_ _10644_/A _10644_/B vssd1 vssd1 vccd1 vccd1 _10712_/D sky130_fd_sc_hd__xor2_1
X_10575_ _10575_/A vssd1 vssd1 vccd1 vccd1 _10707_/A sky130_fd_sc_hd__inv_4
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10108__B _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09202__A1 _09201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10009_ _10010_/B _10010_/A vssd1 vssd1 vccd1 vccd1 _10184_/A sky130_fd_sc_hd__or2_1
XANTENNA__09632__B _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08529__A _09971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05550_ _05600_/A vssd1 vssd1 vccd1 vccd1 _05553_/A sky130_fd_sc_hd__inv_2
XANTENNA__07152__B _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06049__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_328 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05481_ _05497_/A _05497_/B vssd1 vssd1 vccd1 vccd1 _05496_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07220_ _10275_/B _10156_/A vssd1 vssd1 vccd1 vccd1 _07221_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_54_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07151_ _07319_/A _07320_/B vssd1 vssd1 vccd1 vccd1 _07323_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_6_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06102_ _06921_/B _06102_/B vssd1 vssd1 vccd1 vccd1 _06104_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05400__B _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07082_ _07084_/B vssd1 vssd1 vccd1 vccd1 _07083_/B sky130_fd_sc_hd__inv_2
X_06033_ _06032_/B _06841_/B _06033_/C vssd1 vssd1 vccd1 vccd1 _06841_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_1_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06512__A _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07984_ _07986_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07985_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09723_ _10060_/A _09729_/B vssd1 vssd1 vccd1 vccd1 _09896_/B sky130_fd_sc_hd__nand2_1
X_06935_ _07284_/B _06935_/B vssd1 vssd1 vccd1 vccd1 _06937_/A sky130_fd_sc_hd__nand2_1
X_06866_ _06866_/A _06866_/B vssd1 vssd1 vccd1 vccd1 _06867_/B sky130_fd_sc_hd__nand2_1
X_09654_ _09654_/A vssd1 vssd1 vccd1 vccd1 _09932_/B sky130_fd_sc_hd__inv_2
X_05817_ _05827_/B _06057_/A vssd1 vssd1 vccd1 vccd1 _05826_/A sky130_fd_sc_hd__nand2_1
X_08605_ _10128_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _08606_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09585_ _09588_/A _09831_/A vssd1 vssd1 vccd1 vccd1 _09586_/A sky130_fd_sc_hd__nand2_1
X_06797_ _06800_/A _06799_/B _08442_/A vssd1 vssd1 vccd1 vccd1 _08822_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08158__B _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08536_ _08488_/B _08488_/A _08486_/A vssd1 vssd1 vccd1 vccd1 _08630_/A sky130_fd_sc_hd__o21a_1
X_05748_ _06227_/C _06227_/B _05747_/Y vssd1 vssd1 vccd1 vccd1 _06106_/A sky130_fd_sc_hd__a21oi_1
X_08467_ _08467_/A _08467_/B vssd1 vssd1 vccd1 vccd1 _08869_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09680__A1 _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05679_ _05683_/B _05680_/A vssd1 vssd1 vccd1 vccd1 _05682_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09680__B2 _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08398_ _09602_/B vssd1 vssd1 vccd1 vccd1 _10188_/A sky130_fd_sc_hd__inv_2
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07418_ _07418_/A _07418_/B vssd1 vssd1 vccd1 vccd1 _07441_/B sky130_fd_sc_hd__nand2_1
X_07349_ _07349_/A _07349_/B vssd1 vssd1 vccd1 vccd1 _07351_/A sky130_fd_sc_hd__nand2_1
X_10360_ _10385_/A _10360_/B vssd1 vssd1 vccd1 vccd1 _10361_/A sky130_fd_sc_hd__nand2_1
X_10291_ _10294_/B _10294_/C vssd1 vssd1 vccd1 vccd1 _10293_/A sky130_fd_sc_hd__nand2_1
X_09019_ _09021_/C vssd1 vssd1 vccd1 vccd1 _09020_/B sky130_fd_sc_hd__inv_2
XFILLER_0_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06182__B1 _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10627_ _10627_/A vssd1 vssd1 vccd1 vccd1 _10630_/B sky130_fd_sc_hd__inv_2
XFILLER_0_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10558_ _10558_/A _10558_/B vssd1 vssd1 vccd1 vccd1 _10559_/A sky130_fd_sc_hd__nand2_1
X_10489_ _10504_/B _10493_/B vssd1 vssd1 vccd1 vccd1 _10492_/A sky130_fd_sc_hd__nand2_1
X_06720_ _10101_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _06722_/A sky130_fd_sc_hd__nand2_1
X_06651_ _06653_/C _06651_/B _06651_/C vssd1 vssd1 vccd1 vccd1 _06654_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__08259__A _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05602_ _05604_/B vssd1 vssd1 vccd1 vccd1 _05603_/B sky130_fd_sc_hd__inv_2
X_09370_ _10101_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _09376_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06582_ _10284_/B _10148_/A vssd1 vssd1 vccd1 vccd1 _07061_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05533_ _05533_/A _05533_/B _05533_/C vssd1 vssd1 vccd1 vccd1 _05631_/C sky130_fd_sc_hd__nand3_1
X_08321_ _08321_/A _08321_/B vssd1 vssd1 vccd1 vccd1 _08355_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08252_ _08252_/A _08252_/B _08252_/C vssd1 vssd1 vccd1 vccd1 _08253_/B sky130_fd_sc_hd__nand3_1
X_05464_ _05913_/B vssd1 vssd1 vccd1 vccd1 _05471_/B sky130_fd_sc_hd__inv_2
XFILLER_0_61_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07203_ _07203_/A _07203_/B _07203_/C vssd1 vssd1 vccd1 vccd1 _07205_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08183_ _08197_/B _08185_/B vssd1 vssd1 vccd1 vccd1 _08184_/A sky130_fd_sc_hd__nand2_1
X_05395_ _05395_/A _05395_/B vssd1 vssd1 vccd1 vccd1 _05396_/A sky130_fd_sc_hd__nand2_1
X_07134_ _07134_/A _07134_/B vssd1 vssd1 vccd1 vccd1 _07298_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07065_ _07065_/A _07065_/B _07065_/C vssd1 vssd1 vccd1 vccd1 _07066_/B sky130_fd_sc_hd__nand3_1
X_06016_ _06106_/B _06016_/B vssd1 vssd1 vccd1 vccd1 _06017_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07967_ _07967_/A _07967_/B vssd1 vssd1 vccd1 vccd1 _07971_/A sky130_fd_sc_hd__nand2_1
X_09706_ _09708_/B vssd1 vssd1 vccd1 vccd1 _09707_/B sky130_fd_sc_hd__inv_2
X_06918_ _06918_/A _06918_/B vssd1 vssd1 vccd1 vccd1 _06925_/B sky130_fd_sc_hd__nand2_1
X_07898_ _07898_/A vssd1 vssd1 vccd1 vccd1 _07899_/C sky130_fd_sc_hd__inv_2
XANTENNA__10211__B _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06849_ _08983_/B _06849_/B vssd1 vssd1 vccd1 vccd1 _06881_/B sky130_fd_sc_hd__nand2_1
X_09637_ _09637_/A _09637_/B vssd1 vssd1 vccd1 vccd1 _09642_/A sky130_fd_sc_hd__nand2_1
X_09568_ _09568_/A _09569_/A vssd1 vssd1 vccd1 vccd1 _09574_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08519_ _08519_/A _08520_/A vssd1 vssd1 vccd1 vccd1 _08523_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09499_ _09213_/A _09214_/C _09219_/A vssd1 vssd1 vccd1 vccd1 _09793_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_80_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08632__A _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10412_ hold62/X vssd1 vssd1 vccd1 vccd1 _10413_/B sky130_fd_sc_hd__inv_2
XFILLER_0_33_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10343_ _10343_/A hold52/X _10343_/C vssd1 vssd1 vccd1 vccd1 _10591_/C sky130_fd_sc_hd__nand3_1
XANTENNA__05975__B _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08351__B _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10274_ _10274_/A _10274_/B vssd1 vssd1 vccd1 vccd1 _10274_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06152__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10712__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09910__B _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06327__A _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08870_ _08964_/B _08964_/C vssd1 vssd1 vccd1 vccd1 _08963_/A sky130_fd_sc_hd__nand2_1
X_07821_ _07821_/A _07824_/A _07821_/C vssd1 vssd1 vccd1 vccd1 _08066_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_19_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09092__B _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10335__A_N _10334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ _07919_/B _07945_/B _07751_/Y vssd1 vssd1 vccd1 vccd1 _07767_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__10031__B _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07683_ _07689_/A _07690_/A _07689_/B vssd1 vssd1 vccd1 vccd1 _07800_/C sky130_fd_sc_hd__nand3_2
X_06703_ _10414_/B vssd1 vssd1 vccd1 vccd1 _10406_/B sky130_fd_sc_hd__inv_2
XANTENNA__09820__B _09835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09422_ _09422_/A _09598_/A vssd1 vssd1 vccd1 vccd1 _09424_/A sky130_fd_sc_hd__nand2_1
X_06634_ _06977_/C _06977_/B _06633_/Y vssd1 vssd1 vccd1 vccd1 _06968_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__08717__A _08725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09353_ _09353_/A _09353_/B vssd1 vssd1 vccd1 vccd1 _09353_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_74_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08304_ _08304_/A _08304_/B _08304_/C vssd1 vssd1 vccd1 vccd1 _08312_/A sky130_fd_sc_hd__or3_1
X_06565_ _06567_/A vssd1 vssd1 vccd1 vccd1 _06566_/B sky130_fd_sc_hd__inv_2
XFILLER_0_74_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09284_ _09557_/B _09284_/B vssd1 vssd1 vccd1 vccd1 _09292_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07340__B _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06496_ _06498_/B _06498_/C vssd1 vssd1 vccd1 vccd1 _06497_/A sky130_fd_sc_hd__nand2_1
X_05516_ _05515_/B _05954_/B _05516_/C vssd1 vssd1 vccd1 vccd1 _05954_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_74_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08235_ _08372_/A _08373_/A vssd1 vssd1 vccd1 vccd1 _08235_/Y sky130_fd_sc_hd__nand2_1
X_05447_ _07891_/B input4/X vssd1 vssd1 vccd1 vccd1 _05454_/B sky130_fd_sc_hd__nand2_1
X_08166_ _08166_/A _08166_/B vssd1 vssd1 vccd1 vccd1 _08167_/A sky130_fd_sc_hd__nand2_1
X_05378_ _05518_/A _05518_/B vssd1 vssd1 vccd1 vccd1 _05384_/C sky130_fd_sc_hd__nand2_2
XANTENNA__08452__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07117_ _07117_/A _07117_/B vssd1 vssd1 vccd1 vccd1 _07427_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09267__B _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08097_ _09710_/B _08337_/A vssd1 vssd1 vccd1 vccd1 _08100_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08171__B _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07048_ _10247_/B _10158_/A vssd1 vssd1 vccd1 vccd1 _07211_/A sky130_fd_sc_hd__nand2_1
X_08999_ _08999_/A vssd1 vssd1 vccd1 vccd1 _09006_/A sky130_fd_sc_hd__inv_2
XFILLER_0_65_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05986__A _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10326_ _10087_/C _10087_/B _10079_/A vssd1 vssd1 vccd1 vccd1 _10329_/B sky130_fd_sc_hd__a21oi_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ _10256_/B _10257_/B _10257_/C vssd1 vssd1 vccd1 vccd1 _10263_/C sky130_fd_sc_hd__nand3b_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10188_ _10188_/A _10188_/B _10188_/C _10188_/D vssd1 vssd1 vccd1 vccd1 _10190_/A
+ sky130_fd_sc_hd__or4_1
XFILLER_0_56_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_339 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06350_ _06546_/B _06545_/A vssd1 vssd1 vccd1 vccd1 _06549_/C sky130_fd_sc_hd__nand2_1
X_06281_ _06283_/A _06281_/B vssd1 vssd1 vccd1 vccd1 _06282_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08020_ input1/X _10129_/A vssd1 vssd1 vccd1 vccd1 _08021_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09971_ _09971_/A _09971_/B _09971_/C vssd1 vssd1 vccd1 vccd1 _09972_/A sky130_fd_sc_hd__nor3_1
X_08922_ _08927_/B _08927_/A vssd1 vssd1 vccd1 vccd1 _08925_/B sky130_fd_sc_hd__nor2_1
X_08853_ _09268_/A _10276_/D _08852_/C vssd1 vssd1 vccd1 vccd1 _08854_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08784_ _09710_/B vssd1 vssd1 vccd1 vccd1 _10248_/D sky130_fd_sc_hd__inv_2
XANTENNA__10042__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05996_ _05996_/A _05996_/B vssd1 vssd1 vccd1 vccd1 _05997_/B sky130_fd_sc_hd__nand2_1
X_07804_ _07804_/A _07804_/B vssd1 vssd1 vccd1 vccd1 _07943_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07335__B _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07735_ _07735_/A _07735_/B vssd1 vssd1 vccd1 vccd1 _07736_/C sky130_fd_sc_hd__nand2_1
X_09405_ _09405_/A _09406_/A vssd1 vssd1 vccd1 vccd1 _09411_/B sky130_fd_sc_hd__nand2_1
X_07666_ _07666_/A _07666_/B vssd1 vssd1 vccd1 vccd1 _07668_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07597_ _07857_/B _07597_/B _07599_/B vssd1 vssd1 vccd1 vccd1 _07598_/B sky130_fd_sc_hd__nand3_1
X_06617_ _06617_/A _06617_/B _06617_/C vssd1 vssd1 vccd1 vccd1 _06957_/C sky130_fd_sc_hd__nand3_1
X_09336_ _09336_/A _09336_/B _09336_/C vssd1 vssd1 vccd1 vccd1 _09354_/C sky130_fd_sc_hd__nand3_1
X_06548_ _06548_/A _06548_/B vssd1 vssd1 vccd1 vccd1 _06549_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09267_ _10211_/A _10247_/B vssd1 vssd1 vccd1 vccd1 _09268_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08218_ _08218_/A vssd1 vssd1 vccd1 vccd1 _08219_/B sky130_fd_sc_hd__inv_2
X_06479_ _06479_/A _06479_/B vssd1 vssd1 vccd1 vccd1 _06480_/A sky130_fd_sc_hd__nand2_1
X_09198_ _09207_/B _09441_/B vssd1 vssd1 vccd1 vccd1 _09206_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08149_ _08149_/A _08149_/B _08149_/C vssd1 vssd1 vccd1 vccd1 _08212_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_30_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08910__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10111_ _10111_/A vssd1 vssd1 vccd1 vccd1 _10120_/B sky130_fd_sc_hd__inv_2
XFILLER_0_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10042_ input46/X _10211_/A _10211_/B _10210_/B vssd1 vssd1 vccd1 vccd1 _10044_/A
+ sky130_fd_sc_hd__and4_1
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 hold30/A vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 hold52/A vssd1 vssd1 vccd1 vccd1 hold52/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold63 hold63/A vssd1 vssd1 vccd1 vccd1 hold63/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09188__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10309_ _10309_/A _10309_/B vssd1 vssd1 vccd1 vccd1 _10311_/A sky130_fd_sc_hd__nand2_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05850_ _05850_/A _06183_/A vssd1 vssd1 vccd1 vccd1 _05851_/B sky130_fd_sc_hd__nand2_1
X_05781_ _08739_/A input40/X vssd1 vssd1 vccd1 vccd1 _05786_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07520_ _07520_/A _07520_/B _07520_/C vssd1 vssd1 vccd1 vccd1 _07667_/C sky130_fd_sc_hd__nand3_2
X_07451_ _07477_/B _07477_/C vssd1 vssd1 vccd1 vccd1 _07476_/A sky130_fd_sc_hd__nand2_1
X_07382_ _10284_/B _10156_/A vssd1 vssd1 vccd1 vccd1 _07383_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06402_ _06579_/C _06579_/B _06575_/A vssd1 vssd1 vccd1 vccd1 _06567_/A sky130_fd_sc_hd__a21oi_2
X_09121_ input52/X _10292_/B vssd1 vssd1 vccd1 vccd1 _09122_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06333_ _06465_/A _06466_/A vssd1 vssd1 vccd1 vccd1 _06333_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09052_ _09052_/A _09052_/B vssd1 vssd1 vccd1 vccd1 _09351_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_25_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06264_ _06264_/A vssd1 vssd1 vccd1 vccd1 _06267_/A sky130_fd_sc_hd__inv_2
XANTENNA__06515__A _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08003_ _08006_/A _08006_/B vssd1 vssd1 vccd1 vccd1 _08109_/B sky130_fd_sc_hd__nand2_1
X_06195_ _06195_/A vssd1 vssd1 vccd1 vccd1 _06369_/B sky130_fd_sc_hd__inv_2
XFILLER_0_4_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09954_ _10103_/A _10103_/B input19/X input24/X vssd1 vssd1 vccd1 vccd1 _09955_/A
+ sky130_fd_sc_hd__and4_1
X_08905_ _08905_/A vssd1 vssd1 vccd1 vccd1 _08905_/Y sky130_fd_sc_hd__inv_2
X_09885_ _10274_/A _10274_/B vssd1 vssd1 vccd1 vccd1 _09889_/B sky130_fd_sc_hd__or2_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _08835_/B _08836_/B _08836_/C vssd1 vssd1 vccd1 vccd1 _08840_/B sky130_fd_sc_hd__nand3b_1
X_08767_ _08767_/A _08767_/B vssd1 vssd1 vccd1 vccd1 _08833_/C sky130_fd_sc_hd__nand2_1
X_05979_ _05979_/A _05980_/A _06796_/A vssd1 vssd1 vccd1 vccd1 _06810_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_67_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08698_ _10201_/A _09678_/C vssd1 vssd1 vccd1 vccd1 _08699_/B sky130_fd_sc_hd__nand2_1
X_07718_ _07717_/B _07718_/B _07718_/C vssd1 vssd1 vccd1 vccd1 _07828_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_67_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07649_ _07649_/A _07649_/B vssd1 vssd1 vccd1 vccd1 _07808_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_82_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10660_ _10660_/A _10660_/B vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__nand2_1
X_09319_ _09351_/A vssd1 vssd1 vccd1 vccd1 _09320_/B sky130_fd_sc_hd__inv_2
XFILLER_0_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10591_ _10591_/A _10707_/A _10591_/C vssd1 vssd1 vccd1 vccd1 _10592_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_35_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput75 hold61/A vssd1 vssd1 vccd1 vccd1 y_o[18] sky130_fd_sc_hd__buf_12
Xoutput86 hold39/A vssd1 vssd1 vccd1 vccd1 y_o[28] sky130_fd_sc_hd__buf_12
Xoutput97 hold59/A vssd1 vssd1 vccd1 vccd1 y_o[9] sky130_fd_sc_hd__buf_12
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10025_ _10025_/A _10183_/A _10229_/A vssd1 vssd1 vccd1 vccd1 _10052_/C sky130_fd_sc_hd__nand3_1
XANTENNA__09190__B _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08256__B1 _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09646__A _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06989__B _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ _06953_/B _06954_/B _06954_/C vssd1 vssd1 vccd1 vccd1 _06952_/A sky130_fd_sc_hd__nand3_1
X_09670_ _09670_/A _09670_/B vssd1 vssd1 vccd1 vccd1 _09673_/A sky130_fd_sc_hd__nand2_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05902_ _05906_/A vssd1 vssd1 vccd1 vccd1 _05905_/A sky130_fd_sc_hd__inv_2
X_06882_ _08984_/A _06888_/B vssd1 vssd1 vccd1 vccd1 _06887_/A sky130_fd_sc_hd__nand2_1
X_08621_ _08621_/A _08622_/A vssd1 vssd1 vccd1 vccd1 _08625_/A sky130_fd_sc_hd__nand2_1
X_05833_ _05833_/A _06091_/A vssd1 vssd1 vccd1 vccd1 _05836_/C sky130_fd_sc_hd__nand2_1
X_05764_ _05738_/C _05738_/B _05730_/Y vssd1 vssd1 vccd1 vccd1 _05854_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08552_ _08552_/A _08552_/B vssd1 vssd1 vccd1 vccd1 _08562_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07503_ _07505_/A _07505_/B vssd1 vssd1 vccd1 vccd1 _07504_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05414__A _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08483_ _10103_/A input17/X vssd1 vssd1 vccd1 vccd1 _08485_/B sky130_fd_sc_hd__nand2_1
X_07434_ _07444_/B _07445_/B _07445_/C vssd1 vssd1 vccd1 vccd1 _07436_/B sky130_fd_sc_hd__nand3_1
X_05695_ _05695_/A _05695_/B vssd1 vssd1 vccd1 vccd1 _05696_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06229__B _06229_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08725__A _08725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07365_ _07365_/A _07365_/B vssd1 vssd1 vccd1 vccd1 _07452_/B sky130_fd_sc_hd__nand2_1
X_09104_ _09105_/A _09104_/B _09105_/B vssd1 vssd1 vccd1 vccd1 _09108_/B sky130_fd_sc_hd__nand3_1
X_07296_ _07298_/A vssd1 vssd1 vccd1 vccd1 _07297_/B sky130_fd_sc_hd__inv_2
XFILLER_0_17_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06316_ _06318_/A _06318_/B vssd1 vssd1 vccd1 vccd1 _06317_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09035_ _09056_/B _09056_/C vssd1 vssd1 vccd1 vccd1 _09055_/A sky130_fd_sc_hd__nand2_1
X_06247_ _06247_/A _06247_/B vssd1 vssd1 vccd1 vccd1 _06413_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09747__B1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06178_ _06299_/B _06178_/B vssd1 vssd1 vccd1 vccd1 _06221_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09937_ _09938_/B _09938_/C _09936_/Y vssd1 vssd1 vccd1 vccd1 _09939_/A sky130_fd_sc_hd__a21bo_1
X_09868_ _10305_/A vssd1 vssd1 vccd1 vccd1 _09869_/B sky130_fd_sc_hd__inv_2
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09799_ _09799_/A _09799_/B vssd1 vssd1 vccd1 vccd1 _09801_/A sky130_fd_sc_hd__nor2_1
X_08819_ _08819_/A _08819_/B vssd1 vssd1 vccd1 vccd1 _08871_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07523__B input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10712_ _10718_/CLK _10712_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold51/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10643_ _10643_/A _10529_/Y vssd1 vssd1 vccd1 vccd1 _10644_/B sky130_fd_sc_hd__or2b_1
XANTENNA__10737__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10574_ _10574_/A _10580_/A vssd1 vssd1 vccd1 vccd1 _10575_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10008_ _10184_/B _10008_/B vssd1 vssd1 vccd1 vccd1 _10010_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05480_ _05898_/A _05480_/B _05480_/C vssd1 vssd1 vccd1 vccd1 _05497_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_39_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07150_ _10211_/B _10112_/A vssd1 vssd1 vccd1 vccd1 _07320_/B sky130_fd_sc_hd__nand2_1
X_06101_ _06101_/A _06101_/B _06101_/C vssd1 vssd1 vccd1 vccd1 _06308_/B sky130_fd_sc_hd__nand3_1
X_07081_ _07081_/A _07081_/B vssd1 vssd1 vccd1 vccd1 _07084_/B sky130_fd_sc_hd__nand2_1
X_06032_ _06032_/A _06032_/B vssd1 vssd1 vccd1 vccd1 _06038_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05409__A _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ _09722_/A _09722_/B _09722_/C vssd1 vssd1 vccd1 vccd1 _09729_/B sky130_fd_sc_hd__nand3_1
X_07983_ _10040_/B _08337_/A vssd1 vssd1 vccd1 vccd1 _07986_/B sky130_fd_sc_hd__nand2_1
X_06934_ _07284_/A vssd1 vssd1 vccd1 vccd1 _06935_/B sky130_fd_sc_hd__inv_2
X_06865_ _06866_/A _06866_/B vssd1 vssd1 vccd1 vccd1 _08842_/B sky130_fd_sc_hd__or2_1
X_09653_ _09655_/B _09655_/A vssd1 vssd1 vccd1 vccd1 _09654_/A sky130_fd_sc_hd__nor2_1
XANTENNA__07624__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09584_ _09584_/A _09821_/A _09584_/C vssd1 vssd1 vccd1 vccd1 _09831_/A sky130_fd_sc_hd__nand3_2
X_05816_ _06057_/B _05816_/B _05816_/C vssd1 vssd1 vccd1 vccd1 _06057_/A sky130_fd_sc_hd__nand3_1
X_08604_ _08604_/A _08604_/B vssd1 vssd1 vccd1 vccd1 _08619_/B sky130_fd_sc_hd__nand2_1
X_06796_ _06796_/A _06796_/B vssd1 vssd1 vccd1 vccd1 _06799_/B sky130_fd_sc_hd__nand2_1
X_08535_ _08539_/A _08604_/A vssd1 vssd1 vccd1 vccd1 _08630_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05747_ _06228_/B _06229_/B vssd1 vssd1 vccd1 vccd1 _05747_/Y sky130_fd_sc_hd__nor2_1
X_08466_ _08465_/B _08466_/B _08466_/C vssd1 vssd1 vccd1 vccd1 _08467_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__09680__A2 _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05678_ _05681_/B vssd1 vssd1 vccd1 vccd1 _05683_/B sky130_fd_sc_hd__inv_2
X_08397_ input64/X vssd1 vssd1 vccd1 vccd1 _09912_/A sky130_fd_sc_hd__inv_2
X_07417_ _07418_/B _07418_/A vssd1 vssd1 vccd1 vccd1 _07835_/C sky130_fd_sc_hd__nor2_2
X_07348_ _07502_/B _07500_/A vssd1 vssd1 vccd1 vccd1 _07348_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07279_ _07279_/A _07279_/B vssd1 vssd1 vccd1 vccd1 _07859_/A sky130_fd_sc_hd__nand2_1
X_10290_ _10290_/A _10290_/B _10290_/C vssd1 vssd1 vccd1 vccd1 _10294_/C sky130_fd_sc_hd__nand3_1
X_09018_ _09018_/A _09018_/B vssd1 vssd1 vccd1 vccd1 _09021_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06182__A1 _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06182__B2 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10626_ hold2/X _10626_/B vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10557_ _10557_/A _10557_/B vssd1 vssd1 vccd1 vccd1 _10694_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_59_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10488_ _10497_/B _10497_/A vssd1 vssd1 vccd1 vccd1 _10504_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09924__A _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06650_ _06650_/A _06652_/C _06652_/B vssd1 vssd1 vccd1 vccd1 _06651_/C sky130_fd_sc_hd__nand3_1
XANTENNA__08259__B _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05601_ _05560_/C _05560_/B _05600_/Y vssd1 vssd1 vccd1 vccd1 _05604_/B sky130_fd_sc_hd__a21oi_2
X_06581_ _06581_/A _06581_/B vssd1 vssd1 vccd1 vccd1 _07096_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05532_ _05532_/A _05894_/B vssd1 vssd1 vccd1 vccd1 _05533_/C sky130_fd_sc_hd__nand2_1
X_08320_ _08320_/A _08320_/B vssd1 vssd1 vccd1 vccd1 _08321_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08251_ _08251_/A _08251_/B _08251_/C vssd1 vssd1 vccd1 vccd1 _08253_/A sky130_fd_sc_hd__nand3_1
X_05463_ _08573_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _05913_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07202_ _07195_/B _07195_/C _07201_/Y vssd1 vssd1 vccd1 vccd1 _07204_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08182_ _08252_/A _08252_/C _08252_/B vssd1 vssd1 vccd1 vccd1 _08195_/B sky130_fd_sc_hd__a21boi_1
X_05394_ _05394_/A _05394_/B _05394_/C vssd1 vssd1 vccd1 vccd1 _05673_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_40_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07133_ _07135_/A _07135_/B vssd1 vssd1 vccd1 vccd1 _07134_/A sky130_fd_sc_hd__nand2_1
X_07064_ _07064_/A _07064_/B vssd1 vssd1 vccd1 vccd1 _07205_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06523__A _07891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06015_ _06015_/A _06015_/B vssd1 vssd1 vccd1 vccd1 _06902_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07966_ _07968_/B _07968_/C vssd1 vssd1 vccd1 vccd1 _07967_/A sky130_fd_sc_hd__nand2_1
X_09705_ _09705_/A _09705_/B vssd1 vssd1 vccd1 vccd1 _09708_/B sky130_fd_sc_hd__nand2_1
X_06917_ _06919_/C vssd1 vssd1 vccd1 vccd1 _06918_/B sky130_fd_sc_hd__inv_2
X_07897_ _08897_/B _07897_/B vssd1 vssd1 vccd1 vccd1 _07898_/A sky130_fd_sc_hd__nand2_1
X_09636_ _09636_/A _09636_/B vssd1 vssd1 vccd1 vccd1 _09637_/B sky130_fd_sc_hd__xnor2_1
X_06848_ _08983_/A vssd1 vssd1 vccd1 vccd1 _06849_/B sky130_fd_sc_hd__inv_2
X_09567_ _09816_/A _09567_/B vssd1 vssd1 vccd1 vccd1 _09569_/A sky130_fd_sc_hd__nand2_1
X_06779_ _10211_/B _10148_/A vssd1 vssd1 vccd1 vccd1 _06780_/B sky130_fd_sc_hd__nand2_1
X_09498_ _09502_/A _09502_/B vssd1 vssd1 vccd1 vccd1 _09793_/B sky130_fd_sc_hd__nand2_1
X_08518_ _08518_/A _08518_/B vssd1 vssd1 vccd1 vccd1 _08520_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08449_ _08449_/A _08449_/B vssd1 vssd1 vccd1 vccd1 _08817_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_65_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10411_ _10419_/A _10419_/C vssd1 vssd1 vccd1 vccd1 _10413_/A sky130_fd_sc_hd__nand2_1
X_10342_ _10342_/A _10342_/B vssd1 vssd1 vccd1 vccd1 _10591_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08632__B _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08351__C _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10273_ _10298_/B _10298_/C vssd1 vssd1 vccd1 vccd1 _10297_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06152__B input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09644__A2 _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08095__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05512__A _07897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06327__B _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10609_ _10611_/A hold18/X vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__nor2_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07820_ _07822_/A _07823_/A vssd1 vssd1 vccd1 vccd1 _07821_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07751_ _07916_/A _07917_/A vssd1 vssd1 vccd1 vccd1 _07751_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06702_ _06702_/A _10410_/C vssd1 vssd1 vccd1 vccd1 _10414_/B sky130_fd_sc_hd__nand2_1
X_07682_ _07682_/A _07682_/B _07682_/C vssd1 vssd1 vccd1 vccd1 _07689_/B sky130_fd_sc_hd__nand3_1
X_09421_ _09421_/A _09421_/B vssd1 vssd1 vccd1 vccd1 _09598_/A sky130_fd_sc_hd__nand2_1
X_06633_ _06973_/A _06974_/B vssd1 vssd1 vccd1 vccd1 _06633_/Y sky130_fd_sc_hd__nor2_1
X_09352_ _09352_/A _09352_/B vssd1 vssd1 vccd1 vccd1 _09358_/A sky130_fd_sc_hd__nand2_1
X_06564_ _06573_/B vssd1 vssd1 vccd1 vccd1 _06571_/A sky130_fd_sc_hd__inv_2
XFILLER_0_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08303_ _08303_/A vssd1 vssd1 vccd1 vccd1 _08304_/C sky130_fd_sc_hd__inv_2
X_05515_ _05515_/A _05515_/B vssd1 vssd1 vccd1 vccd1 _05522_/A sky130_fd_sc_hd__nand2_1
X_09283_ _09557_/A vssd1 vssd1 vccd1 vccd1 _09284_/B sky130_fd_sc_hd__inv_2
XFILLER_0_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06495_ _06495_/A _06495_/B vssd1 vssd1 vccd1 vccd1 _06498_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_62_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08234_ _08373_/B _08373_/C vssd1 vssd1 vccd1 vccd1 _08372_/A sky130_fd_sc_hd__nand2_1
X_05446_ _05454_/A vssd1 vssd1 vccd1 vccd1 _05449_/A sky130_fd_sc_hd__inv_2
XFILLER_0_55_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08165_ _08165_/A vssd1 vssd1 vccd1 vccd1 _08166_/B sky130_fd_sc_hd__inv_2
X_05377_ _05377_/A _05377_/B vssd1 vssd1 vccd1 vccd1 _05384_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_151 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07116_ _07118_/A _07118_/B vssd1 vssd1 vccd1 vccd1 _07117_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08096_ _08100_/A vssd1 vssd1 vccd1 vccd1 _08099_/A sky130_fd_sc_hd__inv_2
XFILLER_0_30_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07047_ _07065_/C _07065_/B vssd1 vssd1 vccd1 vccd1 _07057_/A sky130_fd_sc_hd__nand2_1
X_08998_ _08998_/A _08998_/B vssd1 vssd1 vccd1 vccd1 _09000_/A sky130_fd_sc_hd__nand2_1
X_07949_ _08139_/B _07979_/A vssd1 vssd1 vccd1 vccd1 _07953_/A sky130_fd_sc_hd__nand2_1
X_09619_ _09668_/B vssd1 vssd1 vccd1 vccd1 _09666_/A sky130_fd_sc_hd__inv_2
XFILLER_0_38_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05986__B _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10325_ _10329_/A _10329_/C vssd1 vssd1 vccd1 vccd1 _10328_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10256_ _10256_/A _10256_/B vssd1 vssd1 vccd1 vccd1 _10263_/A sky130_fd_sc_hd__nand2_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10187_ _10187_/A _10187_/B vssd1 vssd1 vccd1 vccd1 _10191_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05507__A _07785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06280_ _06280_/A vssd1 vssd1 vccd1 vccd1 _06283_/A sky130_fd_sc_hd__inv_2
XFILLER_0_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09970_ _10129_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _09971_/C sky130_fd_sc_hd__nand2_1
X_08921_ _08856_/A _08855_/B _08855_/A vssd1 vssd1 vccd1 vccd1 _08927_/A sky130_fd_sc_hd__o21ba_1
X_08852_ _09268_/A _10276_/D _08852_/C vssd1 vssd1 vccd1 vccd1 _08855_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_20_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07803_ _07910_/B _07951_/A vssd1 vssd1 vccd1 vccd1 _07804_/B sky130_fd_sc_hd__nand2_1
X_08783_ _09840_/B _10201_/B vssd1 vssd1 vccd1 vccd1 _08783_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__10042__B _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05995_ _05995_/A _05995_/B _05995_/C vssd1 vssd1 vccd1 vccd1 _05996_/B sky130_fd_sc_hd__nand3_1
X_07734_ _07734_/A _07734_/B vssd1 vssd1 vccd1 vccd1 _07736_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07665_ _07724_/B _07724_/C vssd1 vssd1 vccd1 vccd1 _07723_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07632__A _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09404_ _09404_/A _09611_/A vssd1 vssd1 vccd1 vccd1 _09406_/A sky130_fd_sc_hd__nand2_1
X_06616_ _06616_/A _06616_/B _06616_/C vssd1 vssd1 vccd1 vccd1 _06617_/B sky130_fd_sc_hd__nand3_1
X_07596_ _07596_/A _07596_/B _07596_/C vssd1 vssd1 vccd1 vccd1 _07598_/A sky130_fd_sc_hd__nand3_1
X_09335_ _09335_/A _09335_/B vssd1 vssd1 vccd1 vccd1 _09354_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06547_ _06547_/A _06547_/B _06547_/C vssd1 vssd1 vccd1 vccd1 _06553_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_35_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09266_ _09266_/A vssd1 vssd1 vccd1 vccd1 _09271_/A sky130_fd_sc_hd__inv_2
X_06478_ _06480_/B _06479_/B _06479_/A vssd1 vssd1 vccd1 vccd1 _06481_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_62_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08217_ _08217_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08219_/A sky130_fd_sc_hd__nand2_1
X_05429_ _05429_/A _05429_/B vssd1 vssd1 vccd1 vccd1 _05524_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_62_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09197_ _09195_/Y _09197_/B _09197_/C vssd1 vssd1 vccd1 vccd1 _09441_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08148_ _08148_/A _08148_/B vssd1 vssd1 vccd1 vccd1 _08149_/A sky130_fd_sc_hd__nand2_1
X_08079_ _08079_/A _08079_/B vssd1 vssd1 vccd1 vccd1 _08080_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08910__B input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout98_A fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10110_ _10110_/A _10110_/B vssd1 vssd1 vccd1 vccd1 _10111_/A sky130_fd_sc_hd__nor2_1
X_10041_ _10041_/A vssd1 vssd1 vccd1 vccd1 _10045_/A sky130_fd_sc_hd__inv_2
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 hold31/A vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 hold64/A vssd1 vssd1 vccd1 vccd1 hold64/X sky130_fd_sc_hd__buf_1
Xhold53 hold53/A vssd1 vssd1 vccd1 vccd1 hold53/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08222__A_N _08245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09188__B _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10308_ _10310_/C vssd1 vssd1 vccd1 vccd1 _10309_/B sky130_fd_sc_hd__inv_2
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10239_ _10243_/B _10243_/C vssd1 vssd1 vccd1 vccd1 _10242_/A sky130_fd_sc_hd__nand2_1
X_05780_ _09517_/C _10187_/B vssd1 vssd1 vccd1 vccd1 _05789_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07450_ _07450_/A _07450_/B _07450_/C vssd1 vssd1 vccd1 vccd1 _07477_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_8_104 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07381_ _07384_/A _07384_/B vssd1 vssd1 vccd1 vccd1 _07482_/C sky130_fd_sc_hd__nand2_1
X_06401_ _06401_/A _06401_/B vssd1 vssd1 vccd1 vccd1 _06575_/A sky130_fd_sc_hd__nor2_1
X_09120_ _09123_/B _09564_/B vssd1 vssd1 vccd1 vccd1 _09122_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06332_ _06458_/C _06458_/B _06331_/Y vssd1 vssd1 vccd1 vccd1 _06466_/A sky130_fd_sc_hd__a21oi_2
X_09051_ _09053_/A vssd1 vssd1 vccd1 vccd1 _09052_/B sky130_fd_sc_hd__inv_2
XFILLER_0_44_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08002_ _09749_/B _08574_/A vssd1 vssd1 vccd1 vccd1 _08006_/B sky130_fd_sc_hd__nand2_1
X_06263_ _06267_/B _06264_/A vssd1 vssd1 vccd1 vccd1 _06266_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06194_ _09517_/D input38/X vssd1 vssd1 vccd1 vccd1 _06195_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07627__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09953_ _10101_/A input18/X vssd1 vssd1 vccd1 vccd1 _09958_/A sky130_fd_sc_hd__nand2_1
X_08904_ _08908_/B _09101_/A vssd1 vssd1 vccd1 vccd1 _08907_/A sky130_fd_sc_hd__nand2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _09884_/A _09884_/B vssd1 vssd1 vccd1 vccd1 _10274_/B sky130_fd_sc_hd__nand2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ _08835_/A _08835_/B vssd1 vssd1 vccd1 vccd1 _08840_/A sky130_fd_sc_hd__nand2_1
X_08766_ _08777_/A _08777_/C vssd1 vssd1 vccd1 vccd1 _08806_/B sky130_fd_sc_hd__nand2_1
X_05978_ _06796_/B _05978_/B _05978_/C vssd1 vssd1 vccd1 vccd1 _06796_/A sky130_fd_sc_hd__nand3_1
X_07717_ _07717_/A _07717_/B vssd1 vssd1 vccd1 vccd1 _07828_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07362__A _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08697_ _10212_/B _10005_/A vssd1 vssd1 vccd1 vccd1 _09228_/C sky130_fd_sc_hd__nand2_1
X_07648_ _07648_/A _07486_/Y vssd1 vssd1 vccd1 vccd1 _07649_/B sky130_fd_sc_hd__nor2b_1
X_07579_ _07579_/A _07579_/B _07579_/C vssd1 vssd1 vccd1 vccd1 _07580_/B sky130_fd_sc_hd__nand3_1
X_09318_ _09587_/A _09321_/B vssd1 vssd1 vccd1 vccd1 _09351_/B sky130_fd_sc_hd__nand2_1
X_10590_ hold15/X hold7/X vssd1 vssd1 vccd1 vccd1 _10594_/A sky130_fd_sc_hd__nand2_1
X_09249_ _09251_/B vssd1 vssd1 vccd1 vccd1 _09250_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput76 hold41/A vssd1 vssd1 vccd1 vccd1 y_o[19] sky130_fd_sc_hd__buf_12
Xoutput87 hold1/A vssd1 vssd1 vccd1 vccd1 y_o[29] sky130_fd_sc_hd__buf_12
X_10024_ _10024_/A vssd1 vssd1 vccd1 vccd1 _10229_/A sky130_fd_sc_hd__inv_2
XANTENNA__08368__A _10511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09199__A _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08256__B2 _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08256__A1 _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09646__B _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06351__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06950_ _06647_/Y _06964_/B _06656_/Y vssd1 vssd1 vccd1 vccd1 _06953_/B sky130_fd_sc_hd__a21o_1
X_06881_ _06881_/A _06881_/B _06881_/C vssd1 vssd1 vccd1 vccd1 _06888_/B sky130_fd_sc_hd__nand3_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05901_ input55/X _10156_/B vssd1 vssd1 vccd1 vccd1 _05906_/A sky130_fd_sc_hd__nand2_1
X_05832_ _05831_/B _05832_/B _06091_/B vssd1 vssd1 vccd1 vccd1 _06091_/A sky130_fd_sc_hd__nand3b_1
X_08620_ _08620_/A _08620_/B vssd1 vssd1 vccd1 vccd1 _08622_/A sky130_fd_sc_hd__nand2_1
X_05763_ _05853_/A _05853_/C vssd1 vssd1 vccd1 vccd1 _05855_/A sky130_fd_sc_hd__nand2_1
X_08551_ _08562_/A _08562_/C vssd1 vssd1 vccd1 vccd1 _08554_/A sky130_fd_sc_hd__nand2_1
X_07502_ _07502_/A _07502_/B vssd1 vssd1 vccd1 vccd1 _07505_/B sky130_fd_sc_hd__nand2_1
X_05694_ _06258_/A _06259_/A vssd1 vssd1 vccd1 vccd1 _06243_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05414__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08482_ _10103_/B _10156_/B vssd1 vssd1 vccd1 vccd1 _08485_/A sky130_fd_sc_hd__nand2_1
X_07433_ _07348_/Y _07504_/B _07372_/Y vssd1 vssd1 vccd1 vccd1 _07444_/B sky130_fd_sc_hd__a21o_1
XANTENNA__08725__B _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09103_ _09539_/A _09539_/B _09103_/C vssd1 vssd1 vccd1 vccd1 _09105_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07364_ _07364_/A _07364_/B vssd1 vssd1 vccd1 vccd1 _07452_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07295_ _07566_/B _07566_/C vssd1 vssd1 vccd1 vccd1 _07565_/A sky130_fd_sc_hd__nand2_1
X_06315_ _06315_/A _06315_/B _06315_/C vssd1 vssd1 vccd1 vccd1 _06318_/B sky130_fd_sc_hd__nand3_1
X_09034_ _09034_/A _09034_/B _09034_/C vssd1 vssd1 vccd1 vccd1 _09056_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_32_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06246_ _06248_/A _06248_/B vssd1 vssd1 vccd1 vccd1 _06247_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09747__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09747__B2 _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06177_ _06299_/A vssd1 vssd1 vccd1 vccd1 _06178_/B sky130_fd_sc_hd__inv_2
XFILLER_0_13_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09936_ _09936_/A _09936_/B vssd1 vssd1 vccd1 vccd1 _09936_/Y sky130_fd_sc_hd__nand2_1
X_09867_ _09768_/C _09768_/B _09763_/Y vssd1 vssd1 vccd1 vccd1 _10305_/A sky130_fd_sc_hd__a21oi_2
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09798_ _09804_/A _09804_/C vssd1 vssd1 vccd1 vccd1 _09803_/A sky130_fd_sc_hd__nand2_1
X_08818_ _08872_/A _08872_/B vssd1 vssd1 vccd1 vccd1 _08871_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08188__A _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08749_ _08749_/A vssd1 vssd1 vccd1 vccd1 _08750_/B sky130_fd_sc_hd__inv_2
XFILLER_0_67_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10711_ _10718_/CLK hold24/X fanout99/X vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__dfrtp_1
X_10642_ _10642_/A _10642_/B vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__xor2_1
X_10573_ _10573_/A _10573_/B hold64/X vssd1 vssd1 vccd1 vccd1 _10580_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10007_ _10187_/A _10005_/A _09602_/B _09678_/C vssd1 vssd1 vccd1 vccd1 _10008_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_39_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06100_ _06921_/B _06921_/A vssd1 vssd1 vccd1 vccd1 _06101_/C sky130_fd_sc_hd__nand2_1
X_07080_ _07080_/A _07097_/A vssd1 vssd1 vccd1 vccd1 _07081_/A sky130_fd_sc_hd__nand2_1
X_06031_ _10247_/B _10187_/B vssd1 vssd1 vccd1 vccd1 _06032_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07982_ _09517_/D _08171_/B vssd1 vssd1 vccd1 vccd1 _07986_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05409__B _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09721_ _09721_/A _09721_/B vssd1 vssd1 vccd1 vccd1 _10060_/A sky130_fd_sc_hd__nand2_1
X_06933_ _09353_/A _06936_/B vssd1 vssd1 vccd1 vccd1 _07284_/B sky130_fd_sc_hd__nand2_1
X_06864_ _08739_/A _09477_/C vssd1 vssd1 vccd1 vccd1 _06866_/B sky130_fd_sc_hd__nand2_1
X_09652_ _09982_/A _09652_/B vssd1 vssd1 vccd1 vccd1 _09655_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07624__B _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09583_ _09583_/A _09583_/B vssd1 vssd1 vccd1 vccd1 _09584_/C sky130_fd_sc_hd__nand2_1
X_05815_ _06057_/B _05816_/C _05816_/B vssd1 vssd1 vccd1 vccd1 _05827_/B sky130_fd_sc_hd__a21o_1
X_06795_ _06799_/A _06800_/B vssd1 vssd1 vccd1 vccd1 _06798_/B sky130_fd_sc_hd__nand2_1
X_08603_ _08623_/A _09185_/B vssd1 vssd1 vccd1 vccd1 _08621_/A sky130_fd_sc_hd__nand2_1
X_08534_ _08533_/B _08604_/B _08534_/C vssd1 vssd1 vccd1 vccd1 _08604_/A sky130_fd_sc_hd__nand3b_1
X_05746_ _06230_/B vssd1 vssd1 vccd1 vccd1 _06227_/B sky130_fd_sc_hd__inv_2
XFILLER_0_77_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08736__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08465_ _08465_/A _08465_/B vssd1 vssd1 vccd1 vccd1 _08467_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05677_ _06240_/B _06240_/C vssd1 vssd1 vccd1 vccd1 _06245_/A sky130_fd_sc_hd__nand2_1
X_08396_ _08703_/A _08396_/B vssd1 vssd1 vccd1 vccd1 _08421_/B sky130_fd_sc_hd__xor2_1
X_07416_ _07403_/A _07405_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07418_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07347_ _07332_/Y _07511_/B _07346_/Y vssd1 vssd1 vccd1 vccd1 _07500_/A sky130_fd_sc_hd__a21oi_1
X_09017_ _09021_/A _09021_/B vssd1 vssd1 vccd1 vccd1 _09020_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07278_ _07856_/B vssd1 vssd1 vccd1 vccd1 _07279_/B sky130_fd_sc_hd__inv_2
XANTENNA__08471__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06229_ _06229_/A _06229_/B vssd1 vssd1 vccd1 vccd1 _06230_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07087__A _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09919_ _09919_/A vssd1 vssd1 vccd1 vccd1 _09921_/A sky130_fd_sc_hd__inv_2
XFILLER_0_68_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06182__A2 _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08646__A _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10625_ hold1/X _10632_/A hold39/A vssd1 vssd1 vccd1 vccd1 _10626_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__09477__A _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10556_ _10678_/A _10556_/B vssd1 vssd1 vccd1 vccd1 _10557_/B sky130_fd_sc_hd__nand2_1
X_10487_ _10487_/A _10487_/B vssd1 vssd1 vccd1 vccd1 _10497_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09924__B _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10151__A _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08259__C _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05600_ _05600_/A _05600_/B vssd1 vssd1 vccd1 vccd1 _05600_/Y sky130_fd_sc_hd__nor2_1
X_06580_ _09551_/C _10188_/B _06400_/C vssd1 vssd1 vccd1 vccd1 _06581_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05531_ _05531_/A _05894_/A vssd1 vssd1 vccd1 vccd1 _05533_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08250_ _08252_/A _08252_/B vssd1 vssd1 vccd1 vccd1 _08251_/A sky130_fd_sc_hd__nand2_1
X_05462_ _05422_/Y _05638_/B _05461_/Y vssd1 vssd1 vccd1 vccd1 _05630_/B sky130_fd_sc_hd__a21o_1
X_07201_ _07201_/A _07201_/B vssd1 vssd1 vccd1 vccd1 _07201_/Y sky130_fd_sc_hd__nor2_1
X_08181_ _08181_/A _08181_/B vssd1 vssd1 vccd1 vccd1 _08252_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07132_ _07132_/A _07132_/B vssd1 vssd1 vccd1 vccd1 _07135_/B sky130_fd_sc_hd__nand2_1
X_05393_ _05395_/A _05393_/B vssd1 vssd1 vccd1 vccd1 _05394_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_40_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07063_ _07203_/C vssd1 vssd1 vccd1 vccd1 _07064_/B sky130_fd_sc_hd__inv_2
X_06014_ _06902_/A _06015_/A _06015_/B vssd1 vssd1 vccd1 vccd1 _06089_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_2_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07965_ _07965_/A _07965_/B vssd1 vssd1 vccd1 vccd1 _07968_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07635__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09704_ _10035_/A _09708_/C vssd1 vssd1 vccd1 vccd1 _09707_/A sky130_fd_sc_hd__nand2_1
X_06916_ _09330_/B _06916_/B vssd1 vssd1 vccd1 vccd1 _06919_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_4_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07896_ _07896_/A _07896_/B vssd1 vssd1 vccd1 vccd1 _07899_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09635_ _09635_/A _09635_/B vssd1 vssd1 vccd1 vccd1 _09636_/B sky130_fd_sc_hd__nand2_1
X_06847_ _06845_/Y _06041_/B _06846_/Y vssd1 vssd1 vccd1 vccd1 _08983_/A sky130_fd_sc_hd__a21oi_2
X_09566_ _09565_/B _09566_/B _09566_/C vssd1 vssd1 vccd1 vccd1 _09567_/B sky130_fd_sc_hd__nand3b_1
X_06778_ _08769_/B _06781_/C vssd1 vssd1 vccd1 vccd1 _06780_/A sky130_fd_sc_hd__nand2_1
X_09497_ _09497_/A _09497_/B _09497_/C vssd1 vssd1 vccd1 vccd1 _09502_/B sky130_fd_sc_hd__nand3_1
X_05729_ _08725_/A input36/X vssd1 vssd1 vccd1 vccd1 _05731_/B sky130_fd_sc_hd__nand2_1
X_08517_ _08517_/A _08517_/B vssd1 vssd1 vccd1 vccd1 _08518_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08448_ _08450_/A _08450_/C vssd1 vssd1 vccd1 vccd1 _08449_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08379_ _10525_/A _08379_/B vssd1 vssd1 vccd1 vccd1 _10467_/B sky130_fd_sc_hd__nand2_1
X_10410_ _10415_/A _10410_/B _10410_/C vssd1 vssd1 vccd1 vccd1 _10419_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_60_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06714__A _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10341_ hold52/X vssd1 vssd1 vccd1 vccd1 _10342_/B sky130_fd_sc_hd__inv_2
X_10272_ _10272_/A _10272_/B _10272_/C vssd1 vssd1 vccd1 vccd1 _10298_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_56_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08095__B _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10608_ _10630_/A hold65/A hold17/X vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_64_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10721__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10539_ _10646_/B _10539_/B vssd1 vssd1 vccd1 vccd1 _10649_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07455__A _08725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07750_ _07946_/B vssd1 vssd1 vccd1 vccd1 _07945_/B sky130_fd_sc_hd__inv_2
X_06701_ _06701_/A _07284_/A _06701_/C vssd1 vssd1 vccd1 vccd1 _10410_/C sky130_fd_sc_hd__nand3_2
X_07681_ _07744_/B _07768_/B _07739_/A vssd1 vssd1 vccd1 vccd1 _07690_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_35_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09420_ _09421_/B _09421_/A vssd1 vssd1 vccd1 vccd1 _09422_/A sky130_fd_sc_hd__or2_1
X_06632_ _06975_/C vssd1 vssd1 vccd1 vccd1 _06977_/B sky130_fd_sc_hd__inv_2
XFILLER_0_59_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09351_ _09351_/A _09351_/B vssd1 vssd1 vccd1 vccd1 _09352_/B sky130_fd_sc_hd__or2_1
X_06563_ _06534_/Y _06664_/A _06562_/Y vssd1 vssd1 vccd1 vccd1 _06573_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_74_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09282_ _09280_/Y _08661_/B _09281_/Y vssd1 vssd1 vccd1 vccd1 _09557_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_47_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08302_ _08302_/A vssd1 vssd1 vccd1 vccd1 _08345_/B sky130_fd_sc_hd__inv_2
X_05514_ _10128_/A _10004_/A vssd1 vssd1 vccd1 vccd1 _05515_/B sky130_fd_sc_hd__nand2_1
X_08233_ _08233_/A _08233_/B vssd1 vssd1 vccd1 vccd1 _08373_/C sky130_fd_sc_hd__nand2_1
X_06494_ _06494_/A vssd1 vssd1 vccd1 vccd1 _06495_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05445_ _07785_/B input5/X vssd1 vssd1 vccd1 vccd1 _05454_/A sky130_fd_sc_hd__nand2_1
X_08164_ _08164_/A vssd1 vssd1 vccd1 vccd1 _08166_/A sky130_fd_sc_hd__inv_2
X_05376_ _05518_/B vssd1 vssd1 vccd1 vccd1 _05377_/B sky130_fd_sc_hd__inv_2
XFILLER_0_42_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08095_ _08112_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _08100_/A sky130_fd_sc_hd__nand2_1
X_07115_ _07115_/A _07115_/B vssd1 vssd1 vccd1 vccd1 _07118_/B sky130_fd_sc_hd__nand2_1
X_07046_ _07046_/A _07046_/B _07046_/C vssd1 vssd1 vccd1 vccd1 _07065_/B sky130_fd_sc_hd__nand3_1
X_08997_ _09003_/B vssd1 vssd1 vccd1 vccd1 _09001_/A sky130_fd_sc_hd__inv_2
X_07948_ _07979_/A _07979_/B _07948_/C vssd1 vssd1 vccd1 vccd1 _08139_/B sky130_fd_sc_hd__nand3_1
X_07879_ _07912_/B vssd1 vssd1 vccd1 vccd1 _07913_/B sky130_fd_sc_hd__inv_2
X_09618_ _09618_/A _09618_/B vssd1 vssd1 vccd1 vccd1 _09668_/B sky130_fd_sc_hd__nand2_1
X_09549_ input52/X vssd1 vssd1 vccd1 vccd1 _10276_/A sky130_fd_sc_hd__inv_2
XANTENNA__05613__A _08725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_171 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06444__A _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10324_ _10324_/A _10324_/B _10324_/C vssd1 vssd1 vccd1 vccd1 _10329_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10255_ _10255_/A _10255_/B vssd1 vssd1 vccd1 vccd1 _10256_/B sky130_fd_sc_hd__nand2_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10186_ _10186_/A vssd1 vssd1 vccd1 vccd1 _10193_/B sky130_fd_sc_hd__inv_2
XANTENNA__05507__B _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08920_ _08920_/A _08920_/B vssd1 vssd1 vccd1 vccd1 _08927_/B sky130_fd_sc_hd__nand2_1
X_08851_ _10211_/A _10275_/B vssd1 vssd1 vccd1 vccd1 _08852_/C sky130_fd_sc_hd__nand2_1
X_07802_ _07951_/A _07951_/B _07950_/B vssd1 vssd1 vccd1 vccd1 _07910_/B sky130_fd_sc_hd__nand3_1
X_08782_ _08782_/A _08782_/B vssd1 vssd1 vccd1 vccd1 _08792_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10042__C _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05994_ _05994_/A vssd1 vssd1 vccd1 vccd1 _05995_/B sky130_fd_sc_hd__inv_2
XFILLER_0_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07733_ _07733_/A _07733_/B _07733_/C vssd1 vssd1 vccd1 vccd1 _07737_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_1_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07664_ _07664_/A _07664_/B _07664_/C vssd1 vssd1 vccd1 vccd1 _07724_/C sky130_fd_sc_hd__nand3_1
XANTENNA__07632__B _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09403_ _09611_/B _09403_/B _09403_/C vssd1 vssd1 vccd1 vccd1 _09611_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_1_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06615_ _06615_/A _06615_/B vssd1 vssd1 vccd1 vccd1 _06617_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05433__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07595_ _07595_/A _07595_/B _07595_/C vssd1 vssd1 vccd1 vccd1 _07596_/C sky130_fd_sc_hd__nand3_1
X_09334_ _09336_/A vssd1 vssd1 vccd1 vccd1 _09335_/B sky130_fd_sc_hd__inv_2
X_06546_ _06548_/B _06546_/B vssd1 vssd1 vccd1 vccd1 _06547_/B sky130_fd_sc_hd__nand2_1
X_09265_ _10210_/A _09840_/B vssd1 vssd1 vccd1 vccd1 _09266_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06477_ _06477_/A _06477_/B _06477_/C vssd1 vssd1 vccd1 vccd1 _06479_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09196_ _09197_/B _09197_/C _09195_/Y vssd1 vssd1 vccd1 vccd1 _09207_/B sky130_fd_sc_hd__a21bo_1
X_08216_ _08245_/A _08245_/B _08216_/C vssd1 vssd1 vccd1 vccd1 _08363_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_28_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05428_ _05430_/B vssd1 vssd1 vccd1 vccd1 _05429_/B sky130_fd_sc_hd__inv_2
XFILLER_0_62_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08147_ _08276_/B _08154_/A vssd1 vssd1 vccd1 vccd1 _08211_/A sky130_fd_sc_hd__nand2_1
X_05359_ input8/X vssd1 vssd1 vccd1 vccd1 _09922_/B sky130_fd_sc_hd__clkbuf_8
X_08078_ _08078_/A _08232_/B vssd1 vssd1 vccd1 vccd1 _08238_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08910__C _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07029_ _07003_/Y _07134_/B _07028_/Y vssd1 vssd1 vccd1 vccd1 _07124_/A sky130_fd_sc_hd__a21oi_2
X_10040_ _10210_/A _10040_/B vssd1 vssd1 vccd1 vccd1 _10041_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05608__A _07756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 hold32/A vssd1 vssd1 vccd1 vccd1 hold32/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 hold65/A vssd1 vssd1 vccd1 vccd1 hold65/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 hold54/A vssd1 vssd1 vccd1 vccd1 hold54/X sky130_fd_sc_hd__buf_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05343__A input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09783__A2 _09782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10307_ _10307_/A _10307_/B vssd1 vssd1 vccd1 vccd1 _10310_/C sky130_fd_sc_hd__nor2_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ _10238_/A _10238_/B _10238_/C vssd1 vssd1 vccd1 vccd1 _10243_/C sky130_fd_sc_hd__nand3_1
X_10169_ _10172_/B _10172_/C vssd1 vssd1 vccd1 vccd1 _10171_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06349__A _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06400_ _09551_/C _10188_/B _06400_/C vssd1 vssd1 vccd1 vccd1 _06579_/B sky130_fd_sc_hd__nor3_2
XFILLER_0_8_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07380_ _09749_/B _10158_/A vssd1 vssd1 vccd1 vccd1 _07384_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_29_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06331_ _06454_/A _06455_/B vssd1 vssd1 vccd1 vccd1 _06331_/Y sky130_fd_sc_hd__nor2_1
X_09050_ _09048_/Y _09071_/B _09049_/Y vssd1 vssd1 vccd1 vccd1 _09053_/A sky130_fd_sc_hd__a21oi_1
X_06262_ _06265_/B vssd1 vssd1 vccd1 vccd1 _06267_/B sky130_fd_sc_hd__inv_2
X_08001_ _09840_/B _08573_/A vssd1 vssd1 vccd1 vccd1 _08006_/A sky130_fd_sc_hd__nand2_1
X_06193_ _06196_/A _06196_/B vssd1 vssd1 vccd1 vccd1 _06369_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_40_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07627__B _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09952_ _09952_/A _09952_/B vssd1 vssd1 vccd1 vccd1 _09961_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_40_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08903_ _08903_/A _08903_/B vssd1 vssd1 vccd1 vccd1 _09101_/A sky130_fd_sc_hd__nand2_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ _09883_/A _09883_/B vssd1 vssd1 vccd1 vccd1 _09884_/B sky130_fd_sc_hd__nand2_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08739__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08834_ _08836_/B _08836_/C vssd1 vssd1 vccd1 vccd1 _08835_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08765_ _08765_/A _08765_/B vssd1 vssd1 vccd1 vccd1 _08777_/A sky130_fd_sc_hd__nand2_1
X_05977_ _05977_/A vssd1 vssd1 vccd1 vccd1 _05978_/B sky130_fd_sc_hd__inv_2
X_07716_ _07718_/B _07718_/C vssd1 vssd1 vccd1 vccd1 _07717_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07362__B _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08696_ _08696_/A vssd1 vssd1 vccd1 vccd1 _08701_/B sky130_fd_sc_hd__inv_2
X_07647_ _07647_/A vssd1 vssd1 vccd1 vccd1 _07875_/A sky130_fd_sc_hd__inv_2
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07578_ _07578_/A _07578_/B vssd1 vssd1 vccd1 vccd1 _07580_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09317_ _09317_/A _09317_/B _09317_/C vssd1 vssd1 vccd1 vccd1 _09321_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_63_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06529_ _07004_/B _07005_/B vssd1 vssd1 vccd1 vccd1 _06530_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_35_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09248_ _09246_/Y _08710_/B _09247_/Y vssd1 vssd1 vccd1 vccd1 _09251_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09179_ _09179_/A _09180_/A vssd1 vssd1 vccd1 vccd1 _09186_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput66 hold50/A vssd1 vssd1 vccd1 vccd1 y_o[0] sky130_fd_sc_hd__buf_12
Xoutput88 hold51/A vssd1 vssd1 vccd1 vccd1 y_o[2] sky130_fd_sc_hd__buf_12
Xoutput77 hold23/A vssd1 vssd1 vccd1 vccd1 y_o[1] sky130_fd_sc_hd__buf_12
X_10023_ _10229_/B _10024_/A vssd1 vssd1 vccd1 vccd1 _10052_/B sky130_fd_sc_hd__nand2_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09199__B _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08256__A2 _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_269 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09646__C _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06351__B input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09943__A _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06880_ _06880_/A _06880_/B vssd1 vssd1 vccd1 vccd1 _08984_/A sky130_fd_sc_hd__nand2_1
X_05900_ _06708_/A vssd1 vssd1 vccd1 vccd1 _05935_/A sky130_fd_sc_hd__inv_2
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05831_ _05831_/A _05831_/B vssd1 vssd1 vccd1 vccd1 _05833_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07463__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05762_ _05761_/B _05793_/B _05762_/C vssd1 vssd1 vccd1 vccd1 _05853_/C sky130_fd_sc_hd__nand3b_1
X_08550_ _08550_/A _08550_/B vssd1 vssd1 vccd1 vccd1 _08562_/A sky130_fd_sc_hd__nand2_1
X_08481_ _10101_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _08488_/B sky130_fd_sc_hd__nand2_1
X_07501_ _07332_/Y _07511_/B _07346_/Y vssd1 vssd1 vccd1 vccd1 _07502_/A sky130_fd_sc_hd__a21o_1
X_05693_ _06268_/C _06268_/B _05692_/Y vssd1 vssd1 vccd1 vccd1 _06259_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_43_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07432_ _07432_/A _07432_/B _07432_/C vssd1 vssd1 vccd1 vccd1 _07442_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_76_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09102_ _09102_/A _09102_/B vssd1 vssd1 vccd1 vccd1 _09104_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07363_ _07365_/B vssd1 vssd1 vccd1 vccd1 _07364_/B sky130_fd_sc_hd__inv_2
XFILLER_0_72_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07294_ _07294_/A _07294_/B _07294_/C vssd1 vssd1 vccd1 vccd1 _07566_/C sky130_fd_sc_hd__nand3_1
X_06314_ _06314_/A _06314_/B vssd1 vssd1 vccd1 vccd1 _06318_/A sky130_fd_sc_hd__nand2_1
X_09033_ _09033_/A _09033_/B vssd1 vssd1 vccd1 vccd1 _09056_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06245_ _06245_/A _06245_/B vssd1 vssd1 vccd1 vccd1 _06248_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09747__A2 _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06176_ _06147_/Y _06236_/B _06175_/Y vssd1 vssd1 vccd1 vccd1 _06299_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_13_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09935_ _09935_/A _10170_/A _10223_/A vssd1 vssd1 vccd1 vccd1 _09938_/C sky130_fd_sc_hd__nand3_1
X_09866_ _09870_/A _09870_/B vssd1 vssd1 vccd1 vccd1 _10305_/B sky130_fd_sc_hd__nand2_1
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08817_ _08817_/A _08817_/B _08817_/C vssd1 vssd1 vccd1 vccd1 _08872_/B sky130_fd_sc_hd__nand3_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08469__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09797_ _09903_/A _10082_/A _09797_/C vssd1 vssd1 vccd1 vccd1 _09804_/C sky130_fd_sc_hd__nand3_1
XANTENNA__10511__B _10511_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08188__B _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08748_ _08748_/A vssd1 vssd1 vccd1 vccd1 _08750_/A sky130_fd_sc_hd__inv_2
X_08679_ _08678_/B _08694_/B _08679_/C vssd1 vssd1 vccd1 vccd1 _08694_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_67_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10710_ _10718_/CLK _10710_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold50/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10641_ _10641_/A _10641_/B vssd1 vssd1 vccd1 vccd1 _10642_/B sky130_fd_sc_hd__nand2_1
X_10572_ _10572_/A _10572_/B vssd1 vssd1 vccd1 vccd1 _10574_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10006_ _10006_/A _10188_/A _10188_/B _10188_/D vssd1 vssd1 vccd1 vccd1 _10184_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_58_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_49 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06627__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07458__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06030_ _08739_/A vssd1 vssd1 vccd1 vccd1 _10247_/B sky130_fd_sc_hd__buf_8
XFILLER_0_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07981_ _08139_/C _08139_/B vssd1 vssd1 vccd1 vccd1 _08026_/B sky130_fd_sc_hd__nand2_1
X_09720_ _09722_/B vssd1 vssd1 vccd1 vccd1 _09721_/B sky130_fd_sc_hd__inv_2
X_06932_ _06932_/A _06932_/B vssd1 vssd1 vccd1 vccd1 _06936_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09362__B1 _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06863_ _09517_/C _09698_/A vssd1 vssd1 vccd1 vccd1 _06866_/A sky130_fd_sc_hd__nand2_1
X_09651_ _09651_/A _09651_/B vssd1 vssd1 vccd1 vccd1 _09652_/B sky130_fd_sc_hd__nand2_1
X_09582_ _09582_/A _09583_/B _09583_/A vssd1 vssd1 vccd1 vccd1 _09588_/A sky130_fd_sc_hd__nand3_1
X_05814_ _05814_/A vssd1 vssd1 vccd1 vccd1 _05816_/B sky130_fd_sc_hd__inv_2
X_06794_ _05978_/B _05978_/C _06796_/B vssd1 vssd1 vccd1 vccd1 _06800_/B sky130_fd_sc_hd__a21boi_1
X_08602_ _08602_/A _08602_/B _09156_/A vssd1 vssd1 vccd1 vccd1 _09185_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_77_401 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08533_ _08533_/A _08533_/B vssd1 vssd1 vccd1 vccd1 _08539_/A sky130_fd_sc_hd__nand2_1
X_05745_ _05745_/A _05745_/B vssd1 vssd1 vccd1 vccd1 _06230_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08736__B _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08464_ _08450_/B _08449_/A _08872_/A vssd1 vssd1 vccd1 vccd1 _08465_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__06537__A _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05676_ _05676_/A _05676_/B _05676_/C vssd1 vssd1 vccd1 vccd1 _06240_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_70_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08395_ _08395_/A _08395_/B vssd1 vssd1 vccd1 vccd1 _08396_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_9_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07415_ _07415_/A _07415_/B vssd1 vssd1 vccd1 vccd1 _07418_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07346_ _07509_/A _07508_/A vssd1 vssd1 vccd1 vccd1 _07346_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_72_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09016_ _09313_/A _09016_/B _09016_/C vssd1 vssd1 vccd1 vccd1 _09021_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_60_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07277_ _07277_/A _07277_/B vssd1 vssd1 vccd1 vccd1 _07279_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08471__B _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06228_ _06228_/A _06228_/B vssd1 vssd1 vccd1 vccd1 _06230_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07087__B _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06159_ _06161_/A _06159_/B vssd1 vssd1 vccd1 vccd1 _06160_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09918_ _09918_/A _09918_/B vssd1 vssd1 vccd1 vccd1 _09919_/A sky130_fd_sc_hd__nand2_1
X_09849_ _09853_/B vssd1 vssd1 vccd1 vccd1 _09854_/C sky130_fd_sc_hd__inv_2
XANTENNA__06447__A _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05351__A _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10624_ _10624_/A hold1/X vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09477__B _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10555_ _10555_/A _10684_/A vssd1 vssd1 vccd1 vccd1 _10556_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_59_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10486_ _10525_/A _10486_/B vssd1 vssd1 vccd1 vccd1 _10487_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08919__B1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__C _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10151__B _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08259__D _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05530_ _05530_/A _05530_/B _05530_/C vssd1 vssd1 vccd1 vccd1 _05631_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05461_ _05634_/A _05636_/B vssd1 vssd1 vccd1 vccd1 _05461_/Y sky130_fd_sc_hd__nor2_1
X_07200_ _07297_/A _07298_/A vssd1 vssd1 vccd1 vccd1 _07200_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_6_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08180_ _08180_/A _08180_/B vssd1 vssd1 vccd1 vccd1 _08181_/A sky130_fd_sc_hd__nand2_1
X_05392_ _05392_/A vssd1 vssd1 vccd1 vccd1 _05395_/A sky130_fd_sc_hd__inv_2
X_07131_ _07303_/B _07131_/B vssd1 vssd1 vccd1 vccd1 _07132_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08572__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07062_ _07062_/A _07062_/B vssd1 vssd1 vccd1 vccd1 _07203_/C sky130_fd_sc_hd__nand2_1
X_06013_ _06013_/A _06013_/B _06013_/C vssd1 vssd1 vccd1 vccd1 _06015_/B sky130_fd_sc_hd__nand3_1
X_07964_ _07964_/A vssd1 vssd1 vccd1 vccd1 _07965_/A sky130_fd_sc_hd__inv_2
XANTENNA__07635__B _07897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09703_ _09703_/A _09703_/B vssd1 vssd1 vccd1 vccd1 _09708_/C sky130_fd_sc_hd__nand2_1
X_06915_ _06915_/A _06915_/B vssd1 vssd1 vccd1 vccd1 _06916_/B sky130_fd_sc_hd__nand2_1
X_07895_ _07895_/A _07895_/B vssd1 vssd1 vccd1 vccd1 _07900_/B sky130_fd_sc_hd__nand2_1
X_06846_ _06846_/A _06846_/B vssd1 vssd1 vccd1 vccd1 _06846_/Y sky130_fd_sc_hd__nor2_1
X_09634_ _10103_/A input22/X _10103_/B input18/X vssd1 vssd1 vccd1 vccd1 _09635_/B
+ sky130_fd_sc_hd__a22o_1
X_09565_ _09565_/A _09565_/B vssd1 vssd1 vccd1 vccd1 _09816_/A sky130_fd_sc_hd__nand2_1
X_06777_ _06777_/A _06777_/B vssd1 vssd1 vccd1 vccd1 _06781_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09496_ _09497_/A _09497_/B _09497_/C vssd1 vssd1 vccd1 vccd1 _09502_/A sky130_fd_sc_hd__a21o_1
X_05728_ _07675_/A input37/X vssd1 vssd1 vccd1 vccd1 _05731_/A sky130_fd_sc_hd__nand2_1
X_08516_ _08517_/A _08516_/B vssd1 vssd1 vccd1 vccd1 _08518_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_77_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08447_ _08447_/A _08447_/B vssd1 vssd1 vccd1 vccd1 _08450_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_18_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05659_ _07785_/B input4/X vssd1 vssd1 vccd1 vccd1 _05664_/A sky130_fd_sc_hd__nand2_1
X_08378_ _10485_/A _08378_/B vssd1 vssd1 vccd1 vccd1 _08379_/B sky130_fd_sc_hd__nor2_1
XANTENNA__08482__A _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06714__B _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07329_ _07518_/C vssd1 vssd1 vccd1 vccd1 _07520_/B sky130_fd_sc_hd__inv_2
X_10340_ _10343_/A _10343_/C vssd1 vssd1 vccd1 vccd1 _10342_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10271_ _10271_/A _10271_/B vssd1 vssd1 vccd1 vccd1 _10298_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06730__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09488__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08392__A _09201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10607_ _10618_/B _10619_/B vssd1 vssd1 vccd1 vccd1 _10611_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_24_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10538_ _10538_/A _10539_/B _10538_/C vssd1 vssd1 vccd1 vccd1 _10646_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_10_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10469_ _10479_/A _10472_/C vssd1 vssd1 vccd1 vccd1 _10471_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07455__B _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06700_ _06700_/A vssd1 vssd1 vccd1 vccd1 _06701_/C sky130_fd_sc_hd__inv_2
X_07680_ _07741_/A _07742_/A vssd1 vssd1 vccd1 vccd1 _07739_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08286__B _08366_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06631_ _10115_/A _10004_/A vssd1 vssd1 vccd1 vccd1 _06975_/C sky130_fd_sc_hd__nand2_1
X_09350_ _10364_/B _09350_/B vssd1 vssd1 vccd1 vccd1 _09352_/A sky130_fd_sc_hd__nand2_1
X_06562_ _06659_/A _06661_/A vssd1 vssd1 vccd1 vccd1 _06562_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_35_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09281_ _09281_/A _09281_/B vssd1 vssd1 vccd1 vccd1 _09281_/Y sky130_fd_sc_hd__nor2_1
X_08301_ _08301_/A _08301_/B vssd1 vssd1 vccd1 vccd1 _08302_/A sky130_fd_sc_hd__xor2_1
X_05513_ input5/X vssd1 vssd1 vccd1 vccd1 _10004_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08232_ _08232_/A _08232_/B _08232_/C vssd1 vssd1 vccd1 vccd1 _08373_/B sky130_fd_sc_hd__nand3_1
X_06493_ _06494_/A _06493_/B _06493_/C vssd1 vssd1 vccd1 vccd1 _06498_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05444_ _05458_/B _05458_/C vssd1 vssd1 vccd1 vccd1 _05457_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08163_ _08254_/B _08255_/A _08162_/Y vssd1 vssd1 vccd1 vccd1 _08181_/B sky130_fd_sc_hd__a21o_1
X_05375_ _08337_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _05518_/B sky130_fd_sc_hd__nand2_1
X_08094_ _08153_/A _08153_/B vssd1 vssd1 vccd1 vccd1 _08151_/A sky130_fd_sc_hd__nand2_1
X_07114_ _07122_/C _07122_/B _07071_/Y vssd1 vssd1 vccd1 vccd1 _07115_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_70_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07045_ _07045_/A _07045_/B vssd1 vssd1 vccd1 vccd1 _07046_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07646__A _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08996_ _08994_/Y _08987_/B _08995_/Y vssd1 vssd1 vccd1 vccd1 _09003_/B sky130_fd_sc_hd__a21oi_1
X_07947_ _07930_/C _07947_/B _07947_/C vssd1 vssd1 vccd1 vccd1 _07979_/A sky130_fd_sc_hd__nand3b_2
X_07878_ _09517_/D _08101_/B vssd1 vssd1 vccd1 vccd1 _07912_/B sky130_fd_sc_hd__nand2_1
X_06829_ _06830_/A _06830_/B vssd1 vssd1 vccd1 vccd1 _08772_/B sky130_fd_sc_hd__or2_1
X_09617_ _09612_/Y _09617_/B _09617_/C vssd1 vssd1 vccd1 vccd1 _09618_/B sky130_fd_sc_hd__nand3b_1
X_09548_ _09555_/A _09555_/B vssd1 vssd1 vccd1 vccd1 _09553_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05613__B input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09479_ _10212_/B _09477_/C _10211_/B _09698_/A vssd1 vssd1 vccd1 vccd1 _09480_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06725__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10247__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10323_ _10323_/A _10323_/B vssd1 vssd1 vccd1 vccd1 _10329_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10254_ _10257_/B _10257_/C vssd1 vssd1 vccd1 vccd1 _10256_/A sky130_fd_sc_hd__nand2_1
X_10185_ _09925_/X _09927_/A _09926_/A vssd1 vssd1 vccd1 vccd1 _10186_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10157__A _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08850__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08850_ _09517_/D vssd1 vssd1 vccd1 vccd1 _10276_/D sky130_fd_sc_hd__inv_2
X_07801_ _07801_/A _07801_/B vssd1 vssd1 vccd1 vccd1 _07804_/A sky130_fd_sc_hd__nand2_1
X_08781_ _08722_/Y _08781_/B _08781_/C vssd1 vssd1 vccd1 vccd1 _08782_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__10042__D _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05993_ _05993_/A _05994_/A vssd1 vssd1 vccd1 vccd1 _05996_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07732_ _07734_/A _07735_/B vssd1 vssd1 vccd1 vccd1 _07733_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07663_ _07663_/A _07663_/B vssd1 vssd1 vccd1 vccd1 _07724_/B sky130_fd_sc_hd__nand2_1
X_09402_ _09402_/A vssd1 vssd1 vccd1 vccd1 _09403_/B sky130_fd_sc_hd__inv_2
XFILLER_0_1_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06614_ _06954_/B _06954_/C vssd1 vssd1 vccd1 vccd1 _06953_/A sky130_fd_sc_hd__nand2_1
X_09333_ _09339_/A _09339_/B _09332_/Y vssd1 vssd1 vccd1 vccd1 _09354_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_47_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07594_ _07594_/A _07594_/B vssd1 vssd1 vccd1 vccd1 _07596_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_62_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06545_ _06545_/A vssd1 vssd1 vccd1 vccd1 _06548_/B sky130_fd_sc_hd__inv_2
X_09264_ _09264_/A _09264_/B vssd1 vssd1 vccd1 vccd1 _09274_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06476_ _06476_/A _06476_/B vssd1 vssd1 vccd1 vccd1 _06479_/B sky130_fd_sc_hd__nand2_1
X_09195_ _08639_/C _08639_/B _08633_/Y vssd1 vssd1 vccd1 vccd1 _09195_/Y sky130_fd_sc_hd__a21oi_1
X_08215_ _08287_/B vssd1 vssd1 vccd1 vccd1 _08216_/C sky130_fd_sc_hd__inv_2
X_05427_ _07785_/B input6/X vssd1 vssd1 vccd1 vccd1 _05430_/B sky130_fd_sc_hd__nand2_1
X_08146_ _08154_/A _08154_/B _08146_/C vssd1 vssd1 vccd1 vccd1 _08276_/B sky130_fd_sc_hd__nand3_1
X_05358_ _08573_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _05392_/A sky130_fd_sc_hd__nand2_1
X_08077_ _08080_/B _08087_/B vssd1 vssd1 vccd1 vccd1 _08078_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08910__D input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07028_ _07127_/A _07132_/A vssd1 vssd1 vccd1 vccd1 _07028_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_30_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05608__B _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09591__A _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08979_ _08995_/A _08980_/A _08980_/B vssd1 vssd1 vccd1 vccd1 _08988_/A sky130_fd_sc_hd__nand3_1
Xhold55 hold55/A vssd1 vssd1 vccd1 vccd1 hold55/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10306_ _10306_/A vssd1 vssd1 vccd1 vccd1 _10307_/B sky130_fd_sc_hd__inv_2
X_10237_ _10237_/A _10237_/B vssd1 vssd1 vccd1 vccd1 _10243_/B sky130_fd_sc_hd__nand2_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10168_ _10166_/Y _10168_/B _10168_/C vssd1 vssd1 vccd1 vccd1 _10172_/C sky130_fd_sc_hd__nand3b_1
X_10099_ _10317_/A vssd1 vssd1 vccd1 vccd1 _10316_/A sky130_fd_sc_hd__inv_2
XANTENNA__06349__B input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06330_ _06456_/C vssd1 vssd1 vccd1 vccd1 _06458_/B sky130_fd_sc_hd__inv_2
X_06261_ _06425_/B _06425_/C vssd1 vssd1 vccd1 vccd1 _06424_/A sky130_fd_sc_hd__nand2_1
X_08000_ _08010_/C _08010_/B vssd1 vssd1 vccd1 vccd1 _08008_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06192_ _08739_/A _10151_/A vssd1 vssd1 vccd1 vccd1 _06196_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09951_ _09952_/B _09952_/A vssd1 vssd1 vccd1 vccd1 _10100_/B sky130_fd_sc_hd__or2_1
X_08902_ _08903_/B _08903_/A vssd1 vssd1 vccd1 vccd1 _08908_/B sky130_fd_sc_hd__or2_1
XANTENNA__10334__B _10334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09882_ _09882_/A vssd1 vssd1 vccd1 vccd1 _09884_/A sky130_fd_sc_hd__inv_2
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _08833_/A _08833_/B _08833_/C vssd1 vssd1 vccd1 vccd1 _08836_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_57_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07924__A _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08764_ _08764_/A vssd1 vssd1 vccd1 vccd1 _08765_/B sky130_fd_sc_hd__inv_2
X_05976_ _05976_/A _05977_/A vssd1 vssd1 vccd1 vccd1 _05980_/A sky130_fd_sc_hd__nand2_1
X_07715_ _07715_/A _07715_/B vssd1 vssd1 vccd1 vccd1 _07718_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_73_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08695_ _10211_/B _10187_/B vssd1 vssd1 vccd1 vccd1 _08696_/A sky130_fd_sc_hd__nand2_1
X_07646_ _09778_/D input1/X _10158_/A _07646_/D vssd1 vssd1 vccd1 vccd1 _07647_/A
+ sky130_fd_sc_hd__and4_1
X_07577_ _07577_/A _07577_/B vssd1 vssd1 vccd1 vccd1 _07584_/A sky130_fd_sc_hd__nor2_1
X_09316_ _09316_/A _09316_/B vssd1 vssd1 vccd1 vccd1 _09587_/A sky130_fd_sc_hd__nand2_2
X_06528_ _07006_/C vssd1 vssd1 vccd1 vccd1 _06530_/B sky130_fd_sc_hd__inv_2
X_09247_ _09247_/A _09247_/B vssd1 vssd1 vccd1 vccd1 _09247_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06459_ _06459_/A _06459_/B vssd1 vssd1 vccd1 vccd1 _06617_/C sky130_fd_sc_hd__nand2_1
X_09178_ _09178_/A _09436_/A vssd1 vssd1 vccd1 vccd1 _09180_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08129_ _08129_/A _08129_/B vssd1 vssd1 vccd1 vccd1 _08133_/B sky130_fd_sc_hd__nand2_1
Xoutput67 hold25/A vssd1 vssd1 vccd1 vccd1 y_o[10] sky130_fd_sc_hd__buf_12
Xoutput89 hold10/A vssd1 vssd1 vccd1 vccd1 y_o[30] sky130_fd_sc_hd__buf_12
Xoutput78 hold64/A vssd1 vssd1 vccd1 vccd1 y_o[20] sky130_fd_sc_hd__buf_12
X_10022_ _10022_/A _10022_/B vssd1 vssd1 vccd1 vccd1 _10024_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09150__A1 _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05830_ input46/X _08897_/B vssd1 vssd1 vccd1 vccd1 _05831_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07463__B _07891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05761_ _05761_/A _05761_/B vssd1 vssd1 vccd1 vccd1 _05853_/A sky130_fd_sc_hd__nand2_1
X_07500_ _07500_/A _07500_/B _07500_/C vssd1 vssd1 vccd1 vccd1 _07505_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_49_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08480_ _08480_/A _08480_/B vssd1 vssd1 vccd1 vccd1 _08549_/A sky130_fd_sc_hd__nand2_1
X_05692_ _06264_/A _06265_/B vssd1 vssd1 vccd1 vccd1 _05692_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_76_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07431_ _07431_/A _07572_/A _07572_/B vssd1 vssd1 vccd1 vccd1 _07848_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_57_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07362_ _09710_/B _10130_/A vssd1 vssd1 vccd1 vccd1 _07365_/B sky130_fd_sc_hd__nand2_1
X_09101_ _09101_/A vssd1 vssd1 vccd1 vccd1 _09102_/B sky130_fd_sc_hd__inv_2
XFILLER_0_72_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06313_ _06315_/A vssd1 vssd1 vccd1 vccd1 _06314_/B sky130_fd_sc_hd__inv_2
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07293_ _07430_/C _07293_/B vssd1 vssd1 vccd1 vccd1 _07294_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_17_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09032_ _09034_/A _09034_/B vssd1 vssd1 vccd1 vccd1 _09033_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06244_ _06425_/B _06244_/B vssd1 vssd1 vccd1 vccd1 _06245_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06175_ _06234_/A _06233_/A vssd1 vssd1 vccd1 vccd1 _06175_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09934_ _09934_/A vssd1 vssd1 vccd1 vccd1 _10223_/A sky130_fd_sc_hd__inv_2
X_09865_ _09861_/B _09865_/B _09865_/C vssd1 vssd1 vccd1 vccd1 _09870_/B sky130_fd_sc_hd__nand3b_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08816_ _08827_/B _08827_/C vssd1 vssd1 vccd1 vccd1 _08894_/B sky130_fd_sc_hd__nand2_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09796_ _10082_/B _09796_/B vssd1 vssd1 vccd1 vccd1 _09804_/A sky130_fd_sc_hd__nand2_1
X_08747_ _08748_/A _08735_/Y _08749_/A vssd1 vssd1 vccd1 vccd1 _08751_/A sky130_fd_sc_hd__o21ai_1
X_05959_ _05961_/C vssd1 vssd1 vccd1 vccd1 _05960_/B sky130_fd_sc_hd__inv_2
X_08678_ _08678_/A _08678_/B vssd1 vssd1 vccd1 vccd1 _08692_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07629_ _07629_/A _07629_/B vssd1 vssd1 vccd1 vccd1 _07684_/A sky130_fd_sc_hd__nor2_1
X_10640_ _10640_/A vssd1 vssd1 vccd1 vccd1 _10710_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10571_ hold64/X vssd1 vssd1 vccd1 vccd1 _10572_/B sky130_fd_sc_hd__inv_2
XFILLER_0_31_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10005_ _10005_/A vssd1 vssd1 vccd1 vccd1 _10188_/D sky130_fd_sc_hd__inv_2
XFILLER_0_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10715__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06627__B _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07458__B _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09954__A _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07980_ _07980_/A _07980_/B vssd1 vssd1 vccd1 vccd1 _08139_/C sky130_fd_sc_hd__nand2_1
X_06931_ _06704_/Y _06310_/B _06705_/Y vssd1 vssd1 vccd1 vccd1 _06932_/B sky130_fd_sc_hd__a21oi_1
X_09650_ _09651_/B _09651_/A vssd1 vssd1 vccd1 vccd1 _09982_/A sky130_fd_sc_hd__or2_1
XANTENNA__09362__A1 _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06862_ _09749_/B _10201_/B vssd1 vssd1 vccd1 vccd1 _06870_/B sky130_fd_sc_hd__nand2_1
X_08601_ _08601_/A _08601_/B vssd1 vssd1 vccd1 vccd1 _08602_/A sky130_fd_sc_hd__nand2_1
X_09581_ _09583_/B _09581_/B _09581_/C vssd1 vssd1 vccd1 vccd1 _09583_/A sky130_fd_sc_hd__nand3_1
X_05813_ input12/X _10201_/B vssd1 vssd1 vccd1 vccd1 _05814_/A sky130_fd_sc_hd__nand2_1
X_06793_ _06800_/A _08442_/A vssd1 vssd1 vccd1 vccd1 _06799_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08532_ _10128_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _08533_/B sky130_fd_sc_hd__nand2_1
X_05744_ _05743_/B _05744_/B _05744_/C vssd1 vssd1 vccd1 vccd1 _05745_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08463_ _08463_/A _08463_/B vssd1 vssd1 vccd1 vccd1 _08872_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07414_ _07414_/A _07414_/B vssd1 vssd1 vccd1 vccd1 _07415_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06537__B _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05675_ _05675_/A _05675_/B vssd1 vssd1 vccd1 vccd1 _06240_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_70_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08394_ _08394_/A vssd1 vssd1 vccd1 vccd1 _08395_/B sky130_fd_sc_hd__inv_2
XFILLER_0_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07345_ _07512_/C vssd1 vssd1 vccd1 vccd1 _07511_/B sky130_fd_sc_hd__inv_2
X_07276_ _07859_/B vssd1 vssd1 vccd1 vccd1 _07276_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09015_ _09313_/B _09015_/B vssd1 vssd1 vccd1 vccd1 _09021_/A sky130_fd_sc_hd__nand2_1
X_06227_ _06227_/A _06227_/B _06227_/C vssd1 vssd1 vccd1 vccd1 _06315_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_13_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06158_ _06158_/A vssd1 vssd1 vccd1 vccd1 _06161_/A sky130_fd_sc_hd__inv_2
X_06089_ _06089_/A _06089_/B _06089_/C vssd1 vssd1 vccd1 vccd1 _06103_/C sky130_fd_sc_hd__nand3_1
X_09917_ _10155_/A _09917_/B vssd1 vssd1 vccd1 vccd1 _09921_/B sky130_fd_sc_hd__nand2_1
X_09848_ _09713_/X _09715_/A _09714_/A vssd1 vssd1 vccd1 vccd1 _09853_/B sky130_fd_sc_hd__a21oi_2
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09779_ _09779_/A vssd1 vssd1 vccd1 vccd1 _09873_/B sky130_fd_sc_hd__inv_2
XFILLER_0_68_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09656__A2 _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06447__B _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05351__B _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10623_ _10623_/A vssd1 vssd1 vccd1 vccd1 _10738_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10554_ _10678_/B _10681_/A _10681_/B vssd1 vssd1 vccd1 vccd1 _10684_/A sky130_fd_sc_hd__nand3_1
XANTENNA__09477__C _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08919__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10485_ _10485_/A vssd1 vssd1 vccd1 vccd1 _10486_/B sky130_fd_sc_hd__inv_2
XANTENNA__08919__B2 _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09924__D _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05542__A _07756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05460_ _05639_/C vssd1 vssd1 vccd1 vccd1 _05638_/B sky130_fd_sc_hd__inv_2
XFILLER_0_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05391_ _05395_/B _05392_/A vssd1 vssd1 vccd1 vccd1 _05394_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07130_ _07131_/B _07130_/B _07130_/C vssd1 vssd1 vccd1 vccd1 _07303_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07061_ _07061_/A _07061_/B vssd1 vssd1 vccd1 vccd1 _07062_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06012_ _06012_/A _06012_/B vssd1 vssd1 vccd1 vccd1 _06015_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07963_ _07964_/A _07963_/B _07963_/C vssd1 vssd1 vccd1 vccd1 _07968_/B sky130_fd_sc_hd__nand3_1
X_09702_ _09703_/B _09703_/A vssd1 vssd1 vccd1 vccd1 _10035_/A sky130_fd_sc_hd__or2_1
XFILLER_0_65_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06914_ _09331_/C vssd1 vssd1 vccd1 vccd1 _09330_/B sky130_fd_sc_hd__inv_2
X_07894_ _07896_/B vssd1 vssd1 vccd1 vccd1 _07895_/B sky130_fd_sc_hd__inv_2
XFILLER_0_4_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06845_ _06846_/B _06846_/A vssd1 vssd1 vccd1 vccd1 _06845_/Y sky130_fd_sc_hd__nand2_1
X_09633_ _09633_/A vssd1 vssd1 vccd1 vccd1 _09635_/A sky130_fd_sc_hd__inv_2
X_09564_ _09564_/A _09564_/B vssd1 vssd1 vccd1 vccd1 _09565_/B sky130_fd_sc_hd__nand2_1
X_06776_ _06777_/A _06777_/B vssd1 vssd1 vccd1 vccd1 _08769_/B sky130_fd_sc_hd__or2_1
X_08515_ _08517_/B vssd1 vssd1 vccd1 vccd1 _08516_/B sky130_fd_sc_hd__inv_2
XANTENNA__05452__A _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09495_ _09495_/A _09744_/A vssd1 vssd1 vccd1 vccd1 _09497_/C sky130_fd_sc_hd__nand2_1
X_05727_ _06121_/B _06121_/A _06120_/B vssd1 vssd1 vccd1 vccd1 _05742_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_81_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08446_ _08447_/A _08402_/Y vssd1 vssd1 vccd1 vccd1 _08450_/A sky130_fd_sc_hd__or2b_1
X_05658_ _08672_/A _07897_/B vssd1 vssd1 vccd1 vccd1 _06125_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_37_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08377_ _10534_/B _10532_/B _10522_/B vssd1 vssd1 vccd1 vccd1 _10485_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05589_ _10158_/A input4/X vssd1 vssd1 vccd1 vccd1 _05592_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07379__A _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07328_ _08672_/A _08114_/B vssd1 vssd1 vccd1 vccd1 _07518_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_33_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08482__B _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07259_ _07579_/A _07579_/B _07578_/B vssd1 vssd1 vccd1 vccd1 _07260_/B sky130_fd_sc_hd__nand3_1
X_10270_ _10272_/C vssd1 vssd1 vccd1 vccd1 _10271_/B sky130_fd_sc_hd__inv_2
XANTENNA__06730__B _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05362__A _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08673__A _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09488__B _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10606_ _10606_/A _10606_/B vssd1 vssd1 vccd1 vccd1 _10619_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_51_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10537_ _10537_/A _10537_/B vssd1 vssd1 vccd1 vccd1 _10538_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_24_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10468_ _10479_/A _10479_/B hold33/X vssd1 vssd1 vccd1 vccd1 _10660_/B sky130_fd_sc_hd__nand3_1
X_10399_ _10399_/A vssd1 vssd1 vccd1 vccd1 _10687_/B sky130_fd_sc_hd__inv_2
XFILLER_0_19_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10730__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ _08114_/B vssd1 vssd1 vccd1 vccd1 _10115_/A sky130_fd_sc_hd__buf_6
XFILLER_0_59_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06561_ _06553_/A _06552_/A _07036_/A vssd1 vssd1 vccd1 vccd1 _06664_/A sky130_fd_sc_hd__o21ai_2
X_09280_ _09281_/B _09281_/A vssd1 vssd1 vccd1 vccd1 _09280_/Y sky130_fd_sc_hd__nand2_1
X_08300_ _08266_/Y _08300_/B vssd1 vssd1 vccd1 vccd1 _08301_/B sky130_fd_sc_hd__nand2b_1
X_05512_ _07897_/B vssd1 vssd1 vccd1 vccd1 _10128_/A sky130_fd_sc_hd__clkbuf_8
X_06492_ _06697_/B vssd1 vssd1 vccd1 vccd1 _06499_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08231_ _08233_/B vssd1 vssd1 vccd1 vccd1 _08232_/A sky130_fd_sc_hd__inv_2
X_05443_ _05443_/A _05583_/A _05524_/A vssd1 vssd1 vccd1 vccd1 _05458_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10337__B _10338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08162_ _08162_/A _08162_/B vssd1 vssd1 vccd1 vccd1 _08162_/Y sky130_fd_sc_hd__nor2_1
X_05374_ input13/X vssd1 vssd1 vccd1 vccd1 _10156_/B sky130_fd_sc_hd__buf_6
XFILLER_0_70_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08093_ _08093_/A _08093_/B vssd1 vssd1 vccd1 vccd1 _08153_/A sky130_fd_sc_hd__nand2_1
X_07113_ _07113_/A _07113_/B _07113_/C vssd1 vssd1 vccd1 vccd1 _07118_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_70_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07044_ _07044_/A _07044_/B _07044_/C vssd1 vssd1 vccd1 vccd1 _07065_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07646__B input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ _08995_/A _08995_/B vssd1 vssd1 vccd1 vccd1 _08995_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__05447__A _07891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07946_ _07946_/A _07946_/B vssd1 vssd1 vccd1 vccd1 _07947_/C sky130_fd_sc_hd__nand2_1
X_07877_ _07889_/A _07889_/C vssd1 vssd1 vccd1 vccd1 _07902_/B sky130_fd_sc_hd__nand2_1
X_06828_ _10210_/B _09678_/C vssd1 vssd1 vccd1 vccd1 _06830_/B sky130_fd_sc_hd__nand2_1
X_09616_ _09612_/Y _09614_/Y _09617_/B vssd1 vssd1 vccd1 vccd1 _09618_/A sky130_fd_sc_hd__o21bai_1
X_09547_ _09547_/A _09547_/B _09799_/A vssd1 vssd1 vccd1 vccd1 _09555_/B sky130_fd_sc_hd__nand3_1
X_06759_ _06763_/A _08819_/B vssd1 vssd1 vccd1 vccd1 _06762_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09478_ _09478_/A vssd1 vssd1 vccd1 vccd1 _09705_/B sky130_fd_sc_hd__inv_2
XFILLER_0_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08429_ _08430_/B _08430_/A vssd1 vssd1 vccd1 vccd1 _08556_/B sky130_fd_sc_hd__or2_1
XANTENNA__06725__B _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10247__B _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10322_ _10324_/C vssd1 vssd1 vccd1 vccd1 _10323_/B sky130_fd_sc_hd__inv_2
XFILLER_0_61_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10253_ _10253_/A _10253_/B vssd1 vssd1 vccd1 vccd1 _10257_/C sky130_fd_sc_hd__nand2_1
X_10184_ _10184_/A _10184_/B vssd1 vssd1 vccd1 vccd1 _10196_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05820__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10157__B _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07747__A _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08780_ _08722_/Y _08779_/Y _08721_/A vssd1 vssd1 vccd1 vccd1 _08782_/A sky130_fd_sc_hd__o21ai_1
X_07800_ _07800_/A _07800_/B _07800_/C vssd1 vssd1 vccd1 vccd1 _07801_/B sky130_fd_sc_hd__nand3_1
X_05992_ _08724_/A _10148_/A vssd1 vssd1 vccd1 vccd1 _05994_/A sky130_fd_sc_hd__nand2_1
X_07731_ _07775_/B _07800_/B vssd1 vssd1 vccd1 vccd1 _07735_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07662_ _07664_/A _07664_/B vssd1 vssd1 vccd1 vccd1 _07663_/A sky130_fd_sc_hd__nand2_1
X_09401_ _09401_/A _09402_/A vssd1 vssd1 vccd1 vccd1 _09404_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07593_ _07848_/A _07593_/B vssd1 vssd1 vccd1 vccd1 _07596_/A sky130_fd_sc_hd__nor2_1
X_06613_ _06613_/A _06613_/B _06613_/C vssd1 vssd1 vccd1 vccd1 _06954_/C sky130_fd_sc_hd__nand3_2
X_09332_ _09340_/C _09340_/B vssd1 vssd1 vccd1 vccd1 _09332_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06544_ _06548_/A _06545_/A vssd1 vssd1 vccd1 vccd1 _06547_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09263_ _09264_/B _09264_/A vssd1 vssd1 vccd1 vccd1 _09534_/B sky130_fd_sc_hd__or2_1
XFILLER_0_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06475_ _06333_/Y _06468_/B _06344_/Y vssd1 vssd1 vccd1 vccd1 _06476_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09194_ _09194_/A _09194_/B vssd1 vssd1 vccd1 vccd1 _09197_/C sky130_fd_sc_hd__nand2_1
X_05426_ input61/X vssd1 vssd1 vccd1 vccd1 _07785_/B sky130_fd_sc_hd__buf_6
X_08214_ _08214_/A _08280_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08287_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_398 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08145_ _08145_/A _08145_/B _08145_/C vssd1 vssd1 vccd1 vccd1 _08154_/B sky130_fd_sc_hd__nand3_1
X_05357_ _05368_/B _05368_/C vssd1 vssd1 vccd1 vccd1 _05501_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_70_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08076_ _08076_/A _08076_/B vssd1 vssd1 vccd1 vccd1 _08080_/B sky130_fd_sc_hd__nand2_1
X_07027_ _07135_/C vssd1 vssd1 vccd1 vccd1 _07134_/B sky130_fd_sc_hd__inv_2
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09591__B _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _08978_/A _08978_/B _08978_/C vssd1 vssd1 vccd1 vccd1 _08980_/B sky130_fd_sc_hd__nand3_1
Xhold56 hold56/A vssd1 vssd1 vccd1 vccd1 hold56/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _07999_/B _07999_/C _07928_/Y vssd1 vssd1 vccd1 vccd1 _07930_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10305_ _10305_/A _10305_/B vssd1 vssd1 vccd1 vccd1 _10307_/A sky130_fd_sc_hd__nor2_1
X_10236_ _10238_/A vssd1 vssd1 vccd1 vccd1 _10237_/B sky130_fd_sc_hd__inv_2
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08398__A _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ _10168_/B _10168_/C _10166_/Y vssd1 vssd1 vccd1 vccd1 _10172_/B sky130_fd_sc_hd__a21bo_1
X_10098_ _10074_/A _10075_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10317_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_16_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06260_ _06260_/A _06260_/B _06260_/C vssd1 vssd1 vccd1 vccd1 _06425_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_32_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06191_ _09517_/C input37/X vssd1 vssd1 vccd1 vccd1 _06196_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09950_ _09950_/A vssd1 vssd1 vccd1 vccd1 _09952_/A sky130_fd_sc_hd__inv_2
X_08901_ _09100_/C _08901_/B vssd1 vssd1 vccd1 vccd1 _08903_/A sky130_fd_sc_hd__xor2_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _09883_/B _09883_/A vssd1 vssd1 vccd1 vccd1 _09882_/A sky130_fd_sc_hd__nor2_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _08832_/A _08832_/B vssd1 vssd1 vccd1 vccd1 _08836_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_57_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07924__B _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ _08763_/A _08763_/B vssd1 vssd1 vccd1 vccd1 _08765_/A sky130_fd_sc_hd__nand2_1
X_05975_ _10201_/A _10156_/A vssd1 vssd1 vccd1 vccd1 _05977_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08101__A _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07714_ _07714_/A _07714_/B vssd1 vssd1 vccd1 vccd1 _07715_/A sky130_fd_sc_hd__nand2_1
X_08694_ _08694_/A _08694_/B vssd1 vssd1 vccd1 vccd1 _08710_/B sky130_fd_sc_hd__nand2_1
X_07645_ _07653_/A _07710_/B vssd1 vssd1 vccd1 vccd1 _07652_/A sky130_fd_sc_hd__nand2_1
X_07576_ _07851_/B vssd1 vssd1 vccd1 vccd1 _07587_/A sky130_fd_sc_hd__inv_2
XFILLER_0_75_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09315_ _09317_/B vssd1 vssd1 vccd1 vccd1 _09316_/B sky130_fd_sc_hd__inv_2
X_06527_ _10040_/B _10128_/A vssd1 vssd1 vccd1 vccd1 _07006_/C sky130_fd_sc_hd__nand2_1
X_09246_ _09247_/B _09247_/A vssd1 vssd1 vccd1 vccd1 _09246_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_35_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06458_ _06458_/A _06458_/B _06458_/C vssd1 vssd1 vccd1 vccd1 _06459_/B sky130_fd_sc_hd__nand3_1
X_05409_ _08337_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _05439_/B sky130_fd_sc_hd__nand2_1
X_09177_ _09176_/B _09177_/B _09436_/B vssd1 vssd1 vccd1 vccd1 _09436_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_16_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06389_ _09517_/D input37/X vssd1 vssd1 vccd1 vccd1 _06394_/A sky130_fd_sc_hd__nand2_1
X_08128_ _09551_/C _09971_/A _08021_/C vssd1 vssd1 vccd1 vccd1 _08129_/B sky130_fd_sc_hd__o21ai_1
X_08059_ _08059_/A _08059_/B vssd1 vssd1 vccd1 vccd1 _08061_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10021_ _10025_/A _10183_/A vssd1 vssd1 vccd1 vccd1 _10229_/B sky130_fd_sc_hd__nand2_1
Xoutput79 hold52/A vssd1 vssd1 vccd1 vccd1 y_o[21] sky130_fd_sc_hd__buf_12
XFILLER_0_11_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput68 hold63/A vssd1 vssd1 vccd1 vccd1 y_o[11] sky130_fd_sc_hd__buf_12
XANTENNA__09150__A2 _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10219_ _10219_/A _10219_/B vssd1 vssd1 vccd1 vccd1 _10227_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05545__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05760_ _09517_/D _10187_/B vssd1 vssd1 vccd1 vccd1 _05761_/B sky130_fd_sc_hd__nand2_1
X_05691_ _06266_/C vssd1 vssd1 vccd1 vccd1 _06268_/B sky130_fd_sc_hd__inv_2
XFILLER_0_76_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07430_ _07430_/A _07430_/B _07430_/C vssd1 vssd1 vccd1 vccd1 _07572_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_43_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07361_ _07365_/A vssd1 vssd1 vccd1 vccd1 _07364_/A sky130_fd_sc_hd__inv_2
X_09100_ _10248_/A _09875_/D _09100_/C vssd1 vssd1 vccd1 vccd1 _09102_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_72_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06312_ _06502_/A _06502_/B vssd1 vssd1 vccd1 vccd1 _06500_/A sky130_fd_sc_hd__nand2_1
X_09031_ _09031_/A _09031_/B _09031_/C vssd1 vssd1 vccd1 vccd1 _09034_/B sky130_fd_sc_hd__nand3_1
X_07292_ _07429_/B vssd1 vssd1 vccd1 vccd1 _07430_/C sky130_fd_sc_hd__inv_2
X_06243_ _06244_/B _06243_/B _06243_/C vssd1 vssd1 vccd1 vccd1 _06425_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06174_ _06166_/A _06165_/A _06477_/B vssd1 vssd1 vccd1 vccd1 _06236_/B sky130_fd_sc_hd__o21ai_2
X_09933_ _10223_/B _09934_/A vssd1 vssd1 vccd1 vccd1 _09938_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09864_ _09864_/A _09864_/B vssd1 vssd1 vccd1 vccd1 _09865_/C sky130_fd_sc_hd__nand2_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08815_ _08815_/A _08815_/B _08815_/C vssd1 vssd1 vccd1 vccd1 _08827_/C sky130_fd_sc_hd__nand3_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _10082_/A vssd1 vssd1 vccd1 vccd1 _09796_/B sky130_fd_sc_hd__inv_2
X_08746_ _08746_/A _08746_/B vssd1 vssd1 vccd1 vccd1 _08749_/A sky130_fd_sc_hd__nand2_1
X_05958_ _05958_/A _05958_/B vssd1 vssd1 vccd1 vccd1 _05961_/C sky130_fd_sc_hd__nand2_1
X_08677_ _10210_/B _10187_/B vssd1 vssd1 vccd1 vccd1 _08678_/B sky130_fd_sc_hd__nand2_1
X_05889_ _06111_/C vssd1 vssd1 vccd1 vccd1 _06110_/B sky130_fd_sc_hd__inv_2
X_07628_ _07687_/B vssd1 vssd1 vccd1 vccd1 _07686_/B sky130_fd_sc_hd__inv_2
XFILLER_0_63_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07559_ _07555_/Y _07717_/B _07558_/Y vssd1 vssd1 vccd1 vccd1 _07604_/A sky130_fd_sc_hd__a21oi_2
X_10570_ _10573_/A _10573_/B vssd1 vssd1 vccd1 vccd1 _10572_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09229_ _09229_/A vssd1 vssd1 vccd1 vccd1 _09243_/B sky130_fd_sc_hd__inv_2
XFILLER_0_63_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10004_ _10004_/A _10187_/B vssd1 vssd1 vccd1 vccd1 _10010_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10699_ _10566_/B _10693_/A _10383_/A vssd1 vssd1 vccd1 vccd1 _10701_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_1_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09954__B _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06930_ _09325_/A _06930_/B vssd1 vssd1 vccd1 vccd1 _06932_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09970__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06861_ _08935_/A _06861_/B vssd1 vssd1 vccd1 vccd1 _06877_/B sky130_fd_sc_hd__nand2_1
X_08600_ _08600_/A _08600_/B vssd1 vssd1 vccd1 vccd1 _08623_/A sky130_fd_sc_hd__nand2_1
X_09580_ _09584_/A _09821_/A vssd1 vssd1 vccd1 vccd1 _09582_/A sky130_fd_sc_hd__nand2_1
X_05812_ input45/X vssd1 vssd1 vccd1 vccd1 _10201_/B sky130_fd_sc_hd__buf_4
X_06792_ _08442_/B _06792_/B _06792_/C vssd1 vssd1 vccd1 vccd1 _08442_/A sky130_fd_sc_hd__nand3_2
XANTENNA__08586__A _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08531_ _08604_/B _08534_/C vssd1 vssd1 vccd1 vccd1 _08533_/A sky130_fd_sc_hd__nand2_1
X_05743_ _05743_/A _05743_/B vssd1 vssd1 vccd1 vccd1 _05745_/A sky130_fd_sc_hd__nand2_1
X_08462_ _08817_/A vssd1 vssd1 vccd1 vccd1 _08463_/B sky130_fd_sc_hd__inv_2
XFILLER_0_49_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05674_ _05676_/A _05676_/B vssd1 vssd1 vccd1 vccd1 _05675_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07413_ _07437_/B _07432_/A vssd1 vssd1 vccd1 vccd1 _07413_/Y sky130_fd_sc_hd__nand2_1
X_08393_ _09201_/A _10202_/B _08392_/C vssd1 vssd1 vccd1 vccd1 _08394_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07344_ _07344_/A _07344_/B vssd1 vssd1 vccd1 vccd1 _07512_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07275_ _07277_/A _07277_/B _07856_/B vssd1 vssd1 vccd1 vccd1 _07859_/B sky130_fd_sc_hd__nand3_1
X_09014_ _09313_/A vssd1 vssd1 vccd1 vccd1 _09015_/B sky130_fd_sc_hd__inv_2
XFILLER_0_60_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06226_ _06228_/A _06229_/A vssd1 vssd1 vccd1 vccd1 _06227_/A sky130_fd_sc_hd__nand2_1
X_06157_ _06161_/B _06158_/A vssd1 vssd1 vccd1 vccd1 _06160_/A sky130_fd_sc_hd__nand2_1
X_06088_ _06088_/A _06088_/B vssd1 vssd1 vccd1 vccd1 _06103_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10091__A _10334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09916_ _09916_/A _09916_/B vssd1 vssd1 vccd1 vccd1 _09917_/B sky130_fd_sc_hd__nand2_1
X_09847_ _10255_/A _09854_/B vssd1 vssd1 vccd1 vccd1 _09853_/A sky130_fd_sc_hd__nand2_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ input52/X input53/X _10275_/B _09778_/D vssd1 vssd1 vccd1 vccd1 _09779_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__08496__A _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08729_ _09710_/B _10201_/B vssd1 vssd1 vccd1 vccd1 _08729_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__09656__A3 _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10622_ hold40/X _10624_/A vssd1 vssd1 vccd1 vccd1 _10623_/A sky130_fd_sc_hd__nor2b_1
XFILLER_0_63_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06744__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ _10553_/A vssd1 vssd1 vccd1 vccd1 _10678_/B sky130_fd_sc_hd__inv_2
XANTENNA__09477__D _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ _10484_/A _10484_/B _10657_/B vssd1 vssd1 vccd1 vccd1 _10510_/A sky130_fd_sc_hd__nand3_1
XANTENNA__08919__A2 _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05542__B _07646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05390_ _05393_/B vssd1 vssd1 vccd1 vccd1 _05395_/B sky130_fd_sc_hd__inv_2
XFILLER_0_27_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07060_ _07060_/A _07060_/B vssd1 vssd1 vccd1 vccd1 _07061_/A sky130_fd_sc_hd__nand2_1
X_06011_ _06013_/C vssd1 vssd1 vccd1 vccd1 _06012_/B sky130_fd_sc_hd__inv_2
XFILLER_0_50_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07485__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09701_ _10035_/B _09701_/B vssd1 vssd1 vccd1 vccd1 _09703_/A sky130_fd_sc_hd__nand2_1
X_07962_ _08058_/C _08058_/B _07961_/Y vssd1 vssd1 vccd1 vccd1 _08069_/A sky130_fd_sc_hd__a21oi_1
X_06913_ _06915_/B _06915_/A vssd1 vssd1 vccd1 vccd1 _09331_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_4_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07893_ _08112_/A _10130_/A vssd1 vssd1 vccd1 vccd1 _07896_/B sky130_fd_sc_hd__nand2_1
X_06844_ _06850_/A _06850_/B vssd1 vssd1 vccd1 vccd1 _08983_/B sky130_fd_sc_hd__nand2_1
X_09632_ _10103_/A _10103_/B input18/X input22/X vssd1 vssd1 vccd1 vccd1 _09633_/A
+ sky130_fd_sc_hd__and4_1
X_09563_ _09566_/B _09566_/C vssd1 vssd1 vccd1 vccd1 _09565_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06775_ _10201_/A _10151_/A vssd1 vssd1 vccd1 vccd1 _06777_/B sky130_fd_sc_hd__nand2_1
X_08514_ _10101_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _08517_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05452__B _07897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09494_ _09744_/B _09494_/B _09494_/C vssd1 vssd1 vccd1 vccd1 _09744_/A sky130_fd_sc_hd__nand3_1
X_05726_ _06121_/C vssd1 vssd1 vccd1 vccd1 _06120_/B sky130_fd_sc_hd__inv_2
XFILLER_0_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08445_ _08445_/A _08445_/B vssd1 vssd1 vccd1 vccd1 _08447_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05657_ _05668_/B _05668_/C vssd1 vssd1 vccd1 vccd1 _05667_/A sky130_fd_sc_hd__nand2_1
X_08376_ _08376_/A _08376_/B vssd1 vssd1 vccd1 vccd1 _10522_/B sky130_fd_sc_hd__nand2_1
X_05588_ input64/X vssd1 vssd1 vccd1 vccd1 _10158_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_73_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07327_ _07516_/A _07517_/B vssd1 vssd1 vccd1 vccd1 _07520_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07379__B _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07258_ _07579_/C vssd1 vssd1 vccd1 vccd1 _07578_/B sky130_fd_sc_hd__inv_2
X_07189_ _07201_/B _07193_/A vssd1 vssd1 vccd1 vccd1 _07192_/B sky130_fd_sc_hd__nand2_1
X_06209_ _06209_/A _06209_/B vssd1 vssd1 vccd1 vccd1 _06386_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05908__A _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05643__A _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05362__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08673__B _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09488__C _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10605_ _10605_/A _10605_/B vssd1 vssd1 vccd1 vccd1 _10606_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_36_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10536_ _10537_/B _10537_/A vssd1 vssd1 vccd1 vccd1 _10539_/B sky130_fd_sc_hd__or2_1
XFILLER_0_3_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10467_ _10467_/A _10467_/B _10467_/C vssd1 vssd1 vccd1 vccd1 _10479_/B sky130_fd_sc_hd__nand3_1
XANTENNA__05818__A input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10398_ _10398_/A _10690_/B vssd1 vssd1 vccd1 vccd1 _10399_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06560_ _06560_/A _06560_/B vssd1 vssd1 vccd1 vccd1 _07036_/A sky130_fd_sc_hd__nand2_1
X_06491_ _06488_/Y _06692_/B _06490_/Y vssd1 vssd1 vccd1 vccd1 _06697_/B sky130_fd_sc_hd__a21oi_1
X_05511_ _05954_/B _05516_/C vssd1 vssd1 vccd1 vccd1 _05515_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08230_ _08376_/B _08376_/A vssd1 vssd1 vccd1 vccd1 _08375_/A sky130_fd_sc_hd__nor2_1
X_05442_ _05583_/B _05442_/B vssd1 vssd1 vccd1 vccd1 _05458_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08161_ _08161_/A vssd1 vssd1 vccd1 vccd1 _08255_/A sky130_fd_sc_hd__inv_2
X_05373_ input33/X vssd1 vssd1 vccd1 vccd1 _08337_/A sky130_fd_sc_hd__buf_8
XFILLER_0_70_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08092_ _08092_/A vssd1 vssd1 vccd1 vccd1 _08093_/B sky130_fd_sc_hd__inv_2
XFILLER_0_15_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07112_ _07595_/B _07595_/C vssd1 vssd1 vccd1 vccd1 _07594_/A sky130_fd_sc_hd__nand2_1
X_07043_ _07045_/B _07043_/B vssd1 vssd1 vccd1 vccd1 _07044_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05728__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07646__C _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08994_ _08995_/B _08995_/A vssd1 vssd1 vccd1 vccd1 _08994_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__05447__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07945_ _07945_/A _07945_/B vssd1 vssd1 vccd1 vccd1 _07947_/B sky130_fd_sc_hd__nand2_1
X_09615_ _09615_/A _09615_/B vssd1 vssd1 vccd1 vccd1 _09617_/B sky130_fd_sc_hd__nand2_1
X_07876_ _07794_/B _07793_/C _07793_/B vssd1 vssd1 vccd1 vccd1 _07889_/A sky130_fd_sc_hd__a21o_1
XANTENNA__05463__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06827_ _10040_/B _10005_/A vssd1 vssd1 vccd1 vccd1 _06830_/A sky130_fd_sc_hd__nand2_1
X_09546_ _09546_/A vssd1 vssd1 vccd1 vccd1 _09799_/A sky130_fd_sc_hd__inv_2
X_06758_ _06758_/A _06758_/B _08435_/A vssd1 vssd1 vccd1 vccd1 _08819_/B sky130_fd_sc_hd__nand3_1
X_09477_ _10212_/B _10211_/B _09477_/C _09698_/A vssd1 vssd1 vccd1 vccd1 _09478_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_65_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05709_ _05709_/A _05709_/B _05709_/C vssd1 vssd1 vccd1 vccd1 _05712_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_38_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08428_ _08541_/B _08428_/B vssd1 vssd1 vccd1 vccd1 _08430_/A sky130_fd_sc_hd__nand2_1
X_06689_ _06689_/A vssd1 vssd1 vccd1 vccd1 _06690_/A sky130_fd_sc_hd__inv_2
XFILLER_0_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08359_ _08359_/A _08359_/B vssd1 vssd1 vccd1 vccd1 _08360_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_33_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10321_ _10321_/A _10321_/B vssd1 vssd1 vccd1 vccd1 _10324_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10252_ _10253_/B _10253_/A vssd1 vssd1 vccd1 vccd1 _10257_/B sky130_fd_sc_hd__or2_1
X_10183_ _10183_/A _10183_/B vssd1 vssd1 vccd1 vccd1 _10199_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08684__A _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05820__B _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10519_ _10642_/A vssd1 vssd1 vccd1 vccd1 _10519_/Y sky130_fd_sc_hd__inv_2
XANTENNA__07747__B _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05991_ _05995_/A _05995_/C vssd1 vssd1 vccd1 vccd1 _05993_/A sky130_fd_sc_hd__nand2_1
X_07730_ _07800_/B _07800_/C _07799_/B vssd1 vssd1 vccd1 vccd1 _07775_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_46_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07661_ _07661_/A _07661_/B vssd1 vssd1 vccd1 vccd1 _07664_/B sky130_fd_sc_hd__nand2_1
X_09400_ _09400_/A _09400_/B vssd1 vssd1 vccd1 vccd1 _09402_/A sky130_fd_sc_hd__nor2_1
X_07592_ _10453_/B _07590_/X _07591_/X vssd1 vssd1 vccd1 vccd1 _07855_/A sky130_fd_sc_hd__o21ai_1
X_06612_ _06612_/A _06612_/B vssd1 vssd1 vccd1 vccd1 _06954_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09331_ _09331_/A _09331_/B _09331_/C vssd1 vssd1 vccd1 vccd1 _09340_/B sky130_fd_sc_hd__nand3_1
X_06543_ _06546_/B vssd1 vssd1 vccd1 vccd1 _06548_/A sky130_fd_sc_hd__inv_2
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09262_ _09262_/A vssd1 vssd1 vccd1 vccd1 _09264_/A sky130_fd_sc_hd__inv_2
X_06474_ _06601_/A _06602_/A vssd1 vssd1 vccd1 vccd1 _06600_/C sky130_fd_sc_hd__nand2_1
X_09193_ _09194_/B _09194_/A vssd1 vssd1 vccd1 vccd1 _09197_/B sky130_fd_sc_hd__or2_1
X_08213_ _08213_/A _08213_/B vssd1 vssd1 vccd1 vccd1 _08280_/B sky130_fd_sc_hd__nand2_1
X_05425_ _05430_/A vssd1 vssd1 vccd1 vccd1 _05429_/A sky130_fd_sc_hd__inv_2
X_08144_ _08144_/A _08144_/B vssd1 vssd1 vccd1 vccd1 _08154_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05356_ _05356_/A _05356_/B _05356_/C vssd1 vssd1 vccd1 vccd1 _05368_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08075_ _08075_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08076_/A sky130_fd_sc_hd__nand2_1
X_07026_ _07026_/A _07026_/B vssd1 vssd1 vccd1 vccd1 _07135_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09872__B _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _08981_/B vssd1 vssd1 vccd1 vccd1 _08995_/A sky130_fd_sc_hd__inv_2
XANTENNA__09591__C _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 hold35/A vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 hold57/A vssd1 vssd1 vccd1 vccd1 hold57/X sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _07994_/A _07995_/A vssd1 vssd1 vccd1 vccd1 _07928_/Y sky130_fd_sc_hd__nor2_1
X_07859_ _07859_/A _07859_/B vssd1 vssd1 vccd1 vccd1 _10431_/B sky130_fd_sc_hd__nand2_1
X_09529_ _09094_/A _09094_/B _09539_/B vssd1 vssd1 vccd1 vccd1 _09530_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_78_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05921__A _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10304_ _10310_/A _10310_/B vssd1 vssd1 vccd1 vccd1 _10309_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09782__B _09782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10235_ _10235_/A _10235_/B vssd1 vssd1 vccd1 vccd1 _10238_/A sky130_fd_sc_hd__nand2_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10166_ _10166_/A _10166_/B vssd1 vssd1 vccd1 vccd1 _10166_/Y sky130_fd_sc_hd__nand2_1
X_10097_ _10573_/A _10339_/C vssd1 vssd1 vccd1 vccd1 _10337_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_325 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06190_ _06217_/B _06217_/C vssd1 vssd1 vccd1 vccd1 _06216_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08900_ input49/X _10275_/B vssd1 vssd1 vccd1 vccd1 _08901_/B sky130_fd_sc_hd__nand2_1
X_09880_ _10280_/A _09880_/B vssd1 vssd1 vccd1 vccd1 _09883_/A sky130_fd_sc_hd__nand2_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _08829_/Y _06842_/B _08830_/Y vssd1 vssd1 vccd1 vccd1 _08840_/C sky130_fd_sc_hd__a21oi_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ _08809_/B _08809_/C vssd1 vssd1 vccd1 vccd1 _08808_/A sky130_fd_sc_hd__nand2_1
X_05974_ _06796_/B _05978_/C vssd1 vssd1 vccd1 vccd1 _05976_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08101__B _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08693_ _08763_/A _08764_/A _08763_/B vssd1 vssd1 vccd1 vccd1 _09287_/B sky130_fd_sc_hd__a21boi_1
X_07713_ _07713_/A _07713_/B _07713_/C vssd1 vssd1 vccd1 vccd1 _07718_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_79_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07644_ _07644_/A _07644_/B _07644_/C vssd1 vssd1 vccd1 vccd1 _07710_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07575_ _07848_/A _07847_/B _07848_/C vssd1 vssd1 vccd1 vccd1 _07851_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_75_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09314_ _09312_/Y _09021_/C _09313_/Y vssd1 vssd1 vccd1 vccd1 _09317_/B sky130_fd_sc_hd__a21oi_1
X_06526_ _07005_/A _07004_/A vssd1 vssd1 vccd1 vccd1 _06531_/B sky130_fd_sc_hd__nand2_1
X_09245_ _09471_/A _09251_/C vssd1 vssd1 vccd1 vccd1 _09250_/A sky130_fd_sc_hd__nand2_1
X_06457_ _06457_/A _06457_/B vssd1 vssd1 vccd1 vccd1 _06458_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05408_ _05439_/A vssd1 vssd1 vccd1 vccd1 _05411_/A sky130_fd_sc_hd__inv_2
XFILLER_0_50_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09176_ _09176_/A _09176_/B vssd1 vssd1 vccd1 vccd1 _09178_/A sky130_fd_sc_hd__nand2_1
X_06388_ _06388_/A _06388_/B vssd1 vssd1 vccd1 vccd1 _06401_/B sky130_fd_sc_hd__nand2_1
X_08127_ _08135_/B _08135_/A vssd1 vssd1 vccd1 vccd1 _08204_/B sky130_fd_sc_hd__nand2_1
X_05339_ input58/X vssd1 vssd1 vccd1 vccd1 _08574_/A sky130_fd_sc_hd__buf_6
XFILLER_0_31_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08058_ _08058_/A _08058_/B _08058_/C vssd1 vssd1 vccd1 vccd1 _08217_/A sky130_fd_sc_hd__nand3_1
X_07009_ _06998_/C _06998_/B _07008_/Y vssd1 vssd1 vccd1 vccd1 _07032_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10020_ _10020_/A _10020_/B _10183_/B vssd1 vssd1 vccd1 vccd1 _10183_/A sky130_fd_sc_hd__nand3_1
Xoutput69 hold36/A vssd1 vssd1 vccd1 vccd1 y_o[12] sky130_fd_sc_hd__buf_12
XANTENNA__06747__A _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10218_ _10220_/B vssd1 vssd1 vccd1 vccd1 _10219_/B sky130_fd_sc_hd__inv_2
X_10149_ _10149_/A vssd1 vssd1 vccd1 vccd1 _10153_/A sky130_fd_sc_hd__inv_2
XANTENNA__05545__B input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05690_ _08114_/B input8/X vssd1 vssd1 vccd1 vccd1 _06266_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_69_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07360_ _10247_/B _10129_/A vssd1 vssd1 vccd1 vccd1 _07365_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09968__A _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06311_ _06310_/B _06311_/B _06311_/C vssd1 vssd1 vccd1 vccd1 _06502_/B sky130_fd_sc_hd__nand3b_2
XFILLER_0_17_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09030_ _09030_/A _09030_/B vssd1 vssd1 vccd1 vccd1 _09034_/A sky130_fd_sc_hd__nand2_1
X_07291_ _07291_/A _07291_/B vssd1 vssd1 vccd1 vccd1 _07566_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_72_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06392__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06242_ _06258_/B _06259_/C _06259_/B vssd1 vssd1 vccd1 vccd1 _06244_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_4_166 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06173_ _06173_/A _06173_/B vssd1 vssd1 vccd1 vccd1 _06477_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09932_ _09932_/A _09932_/B vssd1 vssd1 vccd1 vccd1 _09934_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09863_ _09863_/A vssd1 vssd1 vccd1 vccd1 _09864_/A sky130_fd_sc_hd__inv_2
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08112__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08814_ _08891_/B _09133_/A vssd1 vssd1 vccd1 vccd1 _09082_/B sky130_fd_sc_hd__nand2_1
X_09794_ _09792_/Y _09505_/B _09793_/Y vssd1 vssd1 vccd1 vccd1 _10082_/A sky130_fd_sc_hd__a21oi_2
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08745_ _08745_/A _08745_/B vssd1 vssd1 vccd1 vccd1 _08746_/B sky130_fd_sc_hd__nand2_1
X_05957_ _05957_/A _05957_/B _05957_/C vssd1 vssd1 vccd1 vccd1 _05958_/B sky130_fd_sc_hd__nand3_1
X_08676_ _08694_/B _08679_/C vssd1 vssd1 vccd1 vccd1 _08678_/A sky130_fd_sc_hd__nand2_1
X_05888_ _05888_/A _05888_/B vssd1 vssd1 vccd1 vccd1 _06111_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08340__A1 _09782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07627_ _08739_/A _08101_/B vssd1 vssd1 vccd1 vccd1 _07687_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07558_ _07713_/A _07715_/B vssd1 vssd1 vccd1 vccd1 _07558_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_48_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06509_ _06652_/C _06652_/B vssd1 vssd1 vccd1 vccd1 _06649_/A sky130_fd_sc_hd__nand2_1
X_07489_ _07489_/A _07489_/B vssd1 vssd1 vccd1 vccd1 _07648_/A sky130_fd_sc_hd__nor2_1
X_09228_ _10027_/A _10188_/B _09228_/C vssd1 vssd1 vccd1 vccd1 _09243_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_23_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09159_ _09159_/A _09159_/B _09381_/A vssd1 vssd1 vccd1 vccd1 _09409_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10003_ _10003_/A _10003_/B vssd1 vssd1 vccd1 vccd1 _10020_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05381__A _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10698_ _10698_/A _10698_/B vssd1 vssd1 vccd1 vccd1 hold32/A sky130_fd_sc_hd__xor2_1
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10724__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05556__A input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06860_ _06860_/A _06860_/B vssd1 vssd1 vccd1 vccd1 _06861_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05811_ _05811_/A _05811_/B vssd1 vssd1 vccd1 vccd1 _05816_/C sky130_fd_sc_hd__nand2_1
X_06791_ _08442_/B _06792_/C _06792_/B vssd1 vssd1 vccd1 vccd1 _06800_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08586__B _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08530_ _09971_/A _08529_/B _08529_/C vssd1 vssd1 vccd1 vccd1 _08534_/C sky130_fd_sc_hd__o21ai_1
X_05742_ _06234_/B _05742_/B vssd1 vssd1 vccd1 vccd1 _05743_/B sky130_fd_sc_hd__nand2_1
X_08461_ _08461_/A _08681_/A vssd1 vssd1 vccd1 vccd1 _08817_/A sky130_fd_sc_hd__nand2_1
X_05673_ _05673_/A _05673_/B _05673_/C vssd1 vssd1 vccd1 vccd1 _05676_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09698__A _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07412_ _07435_/C _07435_/B _07411_/Y vssd1 vssd1 vccd1 vccd1 _07432_/A sky130_fd_sc_hd__a21oi_1
X_08392_ _09201_/A _10202_/B _08392_/C vssd1 vssd1 vccd1 vccd1 _08395_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_9_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07343_ _07343_/A _07343_/B _07343_/C vssd1 vssd1 vccd1 vccd1 _07344_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_45_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07274_ _07274_/A _07274_/B _07274_/C vssd1 vssd1 vccd1 vccd1 _07277_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_72_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09013_ _08993_/Y _09027_/B _09012_/Y vssd1 vssd1 vccd1 vccd1 _09313_/A sky130_fd_sc_hd__a21oi_2
X_06225_ _06228_/B vssd1 vssd1 vccd1 vccd1 _06229_/A sky130_fd_sc_hd__inv_2
XFILLER_0_60_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_1__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06156_ _06159_/B vssd1 vssd1 vccd1 vccd1 _06161_/B sky130_fd_sc_hd__inv_2
X_06087_ _06089_/C vssd1 vssd1 vccd1 vccd1 _06088_/B sky130_fd_sc_hd__inv_2
X_09915_ _09916_/B _09916_/A vssd1 vssd1 vccd1 vccd1 _10155_/A sky130_fd_sc_hd__or2_1
XANTENNA__10091__B _10093_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ _09846_/A _09846_/B vssd1 vssd1 vccd1 vccd1 _09854_/B sky130_fd_sc_hd__nand2_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ input54/X vssd1 vssd1 vccd1 vccd1 _09782_/A sky130_fd_sc_hd__inv_2
X_06989_ _10212_/B _08171_/B vssd1 vssd1 vccd1 vccd1 _07008_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08496__B _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08728_ _08726_/A _10202_/C _08726_/C vssd1 vssd1 vccd1 vccd1 _08731_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08659_ _08662_/B _08662_/C vssd1 vssd1 vccd1 vccd1 _08661_/A sky130_fd_sc_hd__nand2_1
X_10621_ _10632_/A hold39/X vssd1 vssd1 vccd1 vccd1 _10624_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06744__B _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10552_ _10552_/A _10682_/B vssd1 vssd1 vccd1 vccd1 _10553_/A sky130_fd_sc_hd__nand2_1
X_10483_ _10483_/A vssd1 vssd1 vccd1 vccd1 _10657_/B sky130_fd_sc_hd__inv_2
XFILLER_0_59_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06010_ _06010_/A _06010_/B vssd1 vssd1 vccd1 vccd1 _06013_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07485__B input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07961_ _08059_/B _08060_/B vssd1 vssd1 vccd1 vccd1 _07961_/Y sky130_fd_sc_hd__nor2_1
X_09700_ _10212_/B _09698_/A _10201_/A _09477_/C vssd1 vssd1 vccd1 vccd1 _09701_/B
+ sky130_fd_sc_hd__a22o_1
X_06912_ _06081_/A _06082_/A _06086_/B vssd1 vssd1 vccd1 vccd1 _06915_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_4_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07892_ _07896_/A vssd1 vssd1 vccd1 vccd1 _07895_/A sky130_fd_sc_hd__inv_2
XFILLER_0_4_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06843_ _06842_/B _06843_/B _06843_/C vssd1 vssd1 vccd1 vccd1 _06850_/B sky130_fd_sc_hd__nand3b_1
X_09631_ _10101_/A input17/X vssd1 vssd1 vccd1 vccd1 _09636_/A sky130_fd_sc_hd__nand2_1
X_09562_ _09800_/A _09562_/B _09815_/A vssd1 vssd1 vccd1 vccd1 _09566_/C sky130_fd_sc_hd__nand3_1
X_06774_ _10212_/B _10150_/A vssd1 vssd1 vccd1 vccd1 _06777_/A sky130_fd_sc_hd__nand2_1
X_05725_ _06120_/A _06121_/C vssd1 vssd1 vccd1 vccd1 _05741_/A sky130_fd_sc_hd__nand2_1
X_08513_ _08513_/A _08513_/B vssd1 vssd1 vccd1 vccd1 _08517_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09493_ _09744_/B _09494_/C _09494_/B vssd1 vssd1 vccd1 vccd1 _09495_/A sky130_fd_sc_hd__a21o_1
X_08444_ _08444_/A vssd1 vssd1 vccd1 vccd1 _08445_/A sky130_fd_sc_hd__inv_2
X_05656_ _05706_/B _05656_/B vssd1 vssd1 vccd1 vccd1 _05668_/C sky130_fd_sc_hd__nand2_1
X_05587_ _05592_/A vssd1 vssd1 vccd1 vccd1 _05591_/A sky130_fd_sc_hd__inv_2
X_08375_ _08375_/A vssd1 vssd1 vccd1 vccd1 _10532_/B sky130_fd_sc_hd__inv_2
XFILLER_0_45_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07326_ _08724_/A input58/X vssd1 vssd1 vccd1 vccd1 _07517_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_73_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07257_ _07578_/A _07579_/C vssd1 vssd1 vccd1 vccd1 _07260_/A sky130_fd_sc_hd__nand2_1
X_07188_ _07167_/C _07167_/B _07187_/Y vssd1 vssd1 vccd1 vccd1 _07193_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07676__A _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06208_ _06210_/B vssd1 vssd1 vccd1 vccd1 _06209_/B sky130_fd_sc_hd__inv_2
XANTENNA__05908__B _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06139_ _06323_/A _06322_/A vssd1 vssd1 vccd1 vccd1 _06253_/B sky130_fd_sc_hd__nand2_1
X_09829_ _10348_/C _10353_/B vssd1 vssd1 vccd1 vccd1 _09830_/B sky130_fd_sc_hd__nor2_1
XANTENNA__05643__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09488__D _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10604_ _10604_/A _10604_/B vssd1 vssd1 vccd1 vccd1 _10606_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_24_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10535_ _10535_/A _10535_/B vssd1 vssd1 vccd1 vccd1 _10537_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10466_ _10466_/A _10466_/B vssd1 vssd1 vccd1 vccd1 _10479_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10397_ _10390_/B _10387_/C hold28/X vssd1 vssd1 vccd1 vccd1 _10398_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_19_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06490_ _06689_/A _06690_/B vssd1 vssd1 vccd1 vccd1 _06490_/Y sky130_fd_sc_hd__nor2_1
X_05510_ _05510_/A _05510_/B vssd1 vssd1 vccd1 vccd1 _05516_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_74_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05441_ _05583_/A vssd1 vssd1 vccd1 vccd1 _05442_/B sky130_fd_sc_hd__inv_2
XANTENNA__10187__A _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08160_ _09749_/B _10115_/A vssd1 vssd1 vccd1 vccd1 _08161_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07111_ _07267_/A _07111_/B _07111_/C vssd1 vssd1 vccd1 vccd1 _07595_/C sky130_fd_sc_hd__nand3_1
X_05372_ _05518_/A vssd1 vssd1 vccd1 vccd1 _05377_/A sky130_fd_sc_hd__inv_2
XFILLER_0_70_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08091_ _08091_/A _08091_/B vssd1 vssd1 vccd1 vccd1 _08093_/A sky130_fd_sc_hd__nand2_1
X_07042_ _07042_/A vssd1 vssd1 vccd1 vccd1 _07045_/B sky130_fd_sc_hd__inv_2
XFILLER_0_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05728__B input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07646__D _07646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ _09024_/A _09025_/A vssd1 vssd1 vccd1 vccd1 _08993_/Y sky130_fd_sc_hd__nand2_1
X_07944_ _07944_/A _07956_/A _07956_/B vssd1 vssd1 vccd1 vccd1 _08041_/A sky130_fd_sc_hd__nand3_2
XANTENNA__09713__B1 _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ _07875_/A _07875_/B vssd1 vssd1 vccd1 vccd1 _07905_/B sky130_fd_sc_hd__nand2_1
X_09614_ _09617_/C vssd1 vssd1 vccd1 vccd1 _09614_/Y sky130_fd_sc_hd__inv_2
X_06826_ _06899_/A _06899_/B vssd1 vssd1 vccd1 vccd1 _06898_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05463__B _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09545_ _09799_/B _09546_/A vssd1 vssd1 vccd1 vccd1 _09555_/A sky130_fd_sc_hd__nand2_1
X_06757_ _06757_/A _06757_/B vssd1 vssd1 vccd1 vccd1 _06763_/A sky130_fd_sc_hd__nand2_1
X_09476_ _10210_/B _10201_/B vssd1 vssd1 vccd1 vccd1 _09482_/B sky130_fd_sc_hd__nand2_1
X_05708_ _05839_/A vssd1 vssd1 vccd1 vccd1 _05711_/A sky130_fd_sc_hd__inv_2
X_06688_ _06689_/A _06688_/B _06688_/C vssd1 vssd1 vccd1 vccd1 _06693_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08427_ _08427_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08428_/B sky130_fd_sc_hd__nand2_1
X_05639_ _05639_/A _05639_/B _05639_/C vssd1 vssd1 vccd1 vccd1 _05640_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_18_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08358_ _08358_/A _08358_/B vssd1 vssd1 vccd1 vccd1 _08359_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_73_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07309_ _07445_/B _07445_/C vssd1 vssd1 vccd1 vccd1 _07444_/A sky130_fd_sc_hd__nand2_1
X_08289_ _08289_/A _08289_/B _08289_/C vssd1 vssd1 vccd1 vccd1 _08325_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10320_ _10320_/A vssd1 vssd1 vccd1 vccd1 _10321_/B sky130_fd_sc_hd__inv_2
XANTENNA__05919__A _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10251_ _10251_/A _10251_/B vssd1 vssd1 vccd1 vccd1 _10253_/A sky130_fd_sc_hd__xnor2_1
X_10182_ _10238_/B _10238_/C vssd1 vssd1 vccd1 vccd1 _10237_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08684__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05829__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10518_ _10638_/B _10638_/A vssd1 vssd1 vccd1 vccd1 _10642_/A sky130_fd_sc_hd__or2_1
XFILLER_0_24_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10449_ _10449_/A _10449_/B vssd1 vssd1 vccd1 vccd1 _10542_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05990_ _05990_/A _05990_/B vssd1 vssd1 vccd1 vccd1 _05995_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_79_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07660_ _07669_/A _07660_/B vssd1 vssd1 vccd1 vccd1 _07661_/B sky130_fd_sc_hd__nand2_1
X_07591_ _07599_/B _07591_/B vssd1 vssd1 vccd1 vccd1 _07591_/X sky130_fd_sc_hd__or2_1
X_06611_ _06613_/A _06613_/B vssd1 vssd1 vccd1 vccd1 _06612_/A sky130_fd_sc_hd__nand2_1
X_09330_ _09330_/A _09330_/B vssd1 vssd1 vccd1 vccd1 _09340_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_1_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06542_ _07046_/C _07046_/B _06541_/Y vssd1 vssd1 vccd1 vccd1 _06553_/A sky130_fd_sc_hd__a21oi_2
X_09261_ _09261_/A _09261_/B vssd1 vssd1 vccd1 vccd1 _09262_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08212_ _08212_/A _08212_/B vssd1 vssd1 vccd1 vccd1 _08213_/B sky130_fd_sc_hd__nand2_1
X_06473_ _06463_/Y _06612_/B _06472_/Y vssd1 vssd1 vccd1 vccd1 _06602_/A sky130_fd_sc_hd__a21oi_1
X_09192_ _09192_/A _09192_/B vssd1 vssd1 vccd1 vccd1 _09194_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_43_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05424_ _07891_/B input5/X vssd1 vssd1 vccd1 vccd1 _05430_/A sky130_fd_sc_hd__nand2_1
X_08143_ _08145_/C _08145_/B vssd1 vssd1 vccd1 vccd1 _08144_/B sky130_fd_sc_hd__nand2_1
X_05355_ _05476_/A _05476_/B vssd1 vssd1 vccd1 vccd1 _05356_/C sky130_fd_sc_hd__nand2_1
X_08074_ _08233_/B _08233_/A vssd1 vssd1 vccd1 vccd1 _08081_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_15_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07025_ _07024_/B _07025_/B _07025_/C vssd1 vssd1 vccd1 vccd1 _07026_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_30_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _08976_/A _08976_/B vssd1 vssd1 vccd1 vccd1 _08981_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09591__D _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold47 hold47/A vssd1 vssd1 vccd1 vccd1 hold47/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 hold36/A vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 hold58/A vssd1 vssd1 vccd1 vccd1 hold58/X sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _07998_/B vssd1 vssd1 vccd1 vccd1 _07999_/C sky130_fd_sc_hd__inv_2
XANTENNA__08785__A _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ _10431_/C _07858_/B vssd1 vssd1 vccd1 vccd1 _10426_/B sky130_fd_sc_hd__nand2_1
X_06809_ _06812_/B _06812_/C vssd1 vssd1 vccd1 vccd1 _06811_/A sky130_fd_sc_hd__nand2_1
X_07789_ _07789_/A _07789_/B vssd1 vssd1 vccd1 vccd1 _07794_/B sky130_fd_sc_hd__nand2_1
X_09528_ _09528_/A _09528_/B vssd1 vssd1 vccd1 vccd1 _09532_/C sky130_fd_sc_hd__nand2_1
XANTENNA__05921__B _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09459_ _09459_/A vssd1 vssd1 vccd1 vccd1 _09459_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_207 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10303_ _10303_/A _10303_/B _10303_/C vssd1 vssd1 vccd1 vccd1 _10310_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10234_ _10234_/A _10234_/B _10234_/C vssd1 vssd1 vccd1 vccd1 _10235_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09925__B1 _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10165_ _10165_/A _10165_/B vssd1 vssd1 vccd1 vccd1 _10168_/C sky130_fd_sc_hd__nand2_1
X_10096_ _10096_/A _10096_/B vssd1 vssd1 vccd1 vccd1 _10573_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08695__A _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _08830_/A _08830_/B vssd1 vssd1 vccd1 vccd1 _08830_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_57_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ _09085_/A _09288_/A _08761_/C vssd1 vssd1 vccd1 vccd1 _08809_/C sky130_fd_sc_hd__nand3_1
X_05973_ _05973_/A _05973_/B vssd1 vssd1 vccd1 vccd1 _05978_/C sky130_fd_sc_hd__nand2_1
X_08692_ _08692_/A _08694_/A _08692_/C vssd1 vssd1 vccd1 vccd1 _08763_/B sky130_fd_sc_hd__nand3_2
X_07712_ _07821_/C _07824_/A _07711_/Y vssd1 vssd1 vccd1 vccd1 _07719_/A sky130_fd_sc_hd__a21o_1
X_07643_ _07643_/A vssd1 vssd1 vccd1 vccd1 _07644_/A sky130_fd_sc_hd__inv_2
X_09313_ _09313_/A _09313_/B vssd1 vssd1 vccd1 vccd1 _09313_/Y sky130_fd_sc_hd__nor2_1
X_07574_ _07577_/B _07577_/A vssd1 vssd1 vccd1 vccd1 _07848_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07014__A _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06525_ _07005_/B vssd1 vssd1 vccd1 vccd1 _07004_/A sky130_fd_sc_hd__inv_2
XANTENNA__06853__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09244_ _09244_/A _09244_/B _09244_/C vssd1 vssd1 vccd1 vccd1 _09251_/C sky130_fd_sc_hd__nand3_1
X_06456_ _06456_/A _06456_/B _06456_/C vssd1 vssd1 vccd1 vccd1 _06459_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09175_ _08609_/A _08609_/B _08616_/B vssd1 vssd1 vccd1 vccd1 _09176_/B sky130_fd_sc_hd__o21a_1
X_05407_ _08171_/B _09602_/B vssd1 vssd1 vccd1 vccd1 _05439_/A sky130_fd_sc_hd__nand2_1
X_08126_ _08126_/A _08138_/A vssd1 vssd1 vccd1 vccd1 _08135_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06387_ _06387_/A _06387_/B vssd1 vssd1 vccd1 vccd1 _06388_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05469__A _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08057_ _08059_/A _08060_/A vssd1 vssd1 vccd1 vccd1 _08058_/A sky130_fd_sc_hd__nand2_1
X_07008_ _07008_/A _07008_/B vssd1 vssd1 vccd1 vccd1 _07008_/Y sky130_fd_sc_hd__nor2_1
X_08959_ _08959_/A _08959_/B _08959_/C vssd1 vssd1 vccd1 vccd1 _09016_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_78_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10217_ _10217_/A _10217_/B vssd1 vssd1 vccd1 vccd1 _10220_/B sky130_fd_sc_hd__nand2_1
X_10148_ _10148_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _10149_/A sky130_fd_sc_hd__nand2_1
X_10079_ _10079_/A vssd1 vssd1 vccd1 vccd1 _10087_/A sky130_fd_sc_hd__inv_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09968__B _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07290_ _07294_/A _07294_/B vssd1 vssd1 vccd1 vccd1 _07291_/A sky130_fd_sc_hd__nand2_1
X_06310_ _06310_/A _06310_/B vssd1 vssd1 vccd1 vccd1 _06502_/A sky130_fd_sc_hd__nand2_1
X_06241_ _06259_/A vssd1 vssd1 vccd1 vccd1 _06258_/B sky130_fd_sc_hd__inv_2
XFILLER_0_72_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06392__B _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06172_ _06320_/C vssd1 vssd1 vccd1 vccd1 _06173_/B sky130_fd_sc_hd__inv_2
XFILLER_0_4_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09931_ _09935_/A _10170_/A vssd1 vssd1 vccd1 vccd1 _10223_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09862_ _09863_/A _09862_/B _10265_/A vssd1 vssd1 vccd1 vccd1 _09865_/B sky130_fd_sc_hd__nand3_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08112__B _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08813_ _09133_/B _08813_/B _08813_/C vssd1 vssd1 vccd1 vccd1 _09133_/A sky130_fd_sc_hd__nand3_2
X_09793_ _09793_/A _09793_/B vssd1 vssd1 vccd1 vccd1 _09793_/Y sky130_fd_sc_hd__nor2_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08744_ _08745_/B _08745_/A vssd1 vssd1 vccd1 vccd1 _08746_/A sky130_fd_sc_hd__or2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05956_ _05956_/A vssd1 vssd1 vccd1 vccd1 _05957_/C sky130_fd_sc_hd__inv_2
X_08675_ _09699_/A _10188_/B _08674_/C vssd1 vssd1 vccd1 vccd1 _08679_/C sky130_fd_sc_hd__o21ai_1
X_05887_ _05887_/A _05887_/B _05887_/C vssd1 vssd1 vccd1 vccd1 _05888_/B sky130_fd_sc_hd__nand3_1
X_07626_ _07629_/A _07629_/B vssd1 vssd1 vccd1 vccd1 _07687_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07557_ _07561_/A _07561_/B vssd1 vssd1 vccd1 vccd1 _07717_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_75_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06508_ _06508_/A _06508_/B _06508_/C vssd1 vssd1 vccd1 vccd1 _06652_/C sky130_fd_sc_hd__nand3_1
X_07488_ _07649_/A vssd1 vssd1 vccd1 vccd1 _07488_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06583__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09227_ _10201_/A vssd1 vssd1 vccd1 vccd1 _10027_/A sky130_fd_sc_hd__inv_2
XFILLER_0_51_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06439_ _06439_/A _06439_/B vssd1 vssd1 vccd1 vccd1 _06440_/A sky130_fd_sc_hd__nand2_1
X_09158_ _09158_/A _09158_/B vssd1 vssd1 vccd1 vccd1 _09181_/A sky130_fd_sc_hd__nand2_1
X_09089_ _09109_/B vssd1 vssd1 vccd1 vccd1 _09107_/A sky130_fd_sc_hd__inv_2
XFILLER_0_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08109_ _08107_/A _08109_/B vssd1 vssd1 vccd1 vccd1 _08120_/A sky130_fd_sc_hd__and2b_1
XFILLER_0_31_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10002_ _10068_/A _10068_/C vssd1 vssd1 vccd1 vccd1 _10066_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10697_ _10697_/A _10697_/B vssd1 vssd1 vccd1 vccd1 _10698_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05810_ _05810_/A _05810_/B vssd1 vssd1 vccd1 vccd1 _06057_/B sky130_fd_sc_hd__nand2_1
X_06790_ _06790_/A vssd1 vssd1 vccd1 vccd1 _06792_/B sky130_fd_sc_hd__inv_2
X_05741_ _05741_/A _05742_/B _05741_/C vssd1 vssd1 vccd1 vccd1 _06234_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08460_ _08459_/Y _08460_/B _08460_/C vssd1 vssd1 vccd1 vccd1 _08681_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_54_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05672_ _05672_/A _05672_/B vssd1 vssd1 vccd1 vccd1 _05676_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08391_ _09677_/A _10150_/A vssd1 vssd1 vccd1 vccd1 _08392_/C sky130_fd_sc_hd__nand2_1
X_07411_ _07445_/A _07444_/A vssd1 vssd1 vccd1 vccd1 _07411_/Y sky130_fd_sc_hd__nor2_1
X_07342_ _07342_/A vssd1 vssd1 vccd1 vccd1 _07343_/B sky130_fd_sc_hd__inv_2
XFILLER_0_45_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07273_ _07273_/A _07273_/B vssd1 vssd1 vccd1 vccd1 _07277_/A sky130_fd_sc_hd__nand2_1
X_09012_ _09025_/A _09024_/A vssd1 vssd1 vccd1 vccd1 _09012_/Y sky130_fd_sc_hd__nor2_1
X_06224_ _06229_/B vssd1 vssd1 vccd1 vccd1 _06228_/A sky130_fd_sc_hd__inv_2
XFILLER_0_5_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06155_ _06361_/C _06361_/B _06154_/Y vssd1 vssd1 vccd1 vccd1 _06166_/A sky130_fd_sc_hd__a21oi_2
X_06086_ _06086_/A _06086_/B vssd1 vssd1 vccd1 vccd1 _06089_/C sky130_fd_sc_hd__nand2_1
XANTENNA__05747__A _06228_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09914_ _10155_/B _09914_/B vssd1 vssd1 vccd1 vccd1 _09916_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09845_ _09846_/B _09846_/A vssd1 vssd1 vccd1 vccd1 _10255_/A sky130_fd_sc_hd__or2_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _09790_/A _09790_/B vssd1 vssd1 vccd1 vccd1 _09789_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05482__A _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06988_ _07008_/B vssd1 vssd1 vccd1 vccd1 _06995_/B sky130_fd_sc_hd__inv_2
X_08727_ _08727_/A vssd1 vssd1 vccd1 vccd1 _09261_/B sky130_fd_sc_hd__inv_2
X_05939_ _07785_/B vssd1 vssd1 vccd1 vccd1 _10130_/A sky130_fd_sc_hd__clkbuf_8
X_08658_ _08658_/A _09281_/A vssd1 vssd1 vccd1 vccd1 _08662_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08793__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07609_ _07721_/B _07721_/C vssd1 vssd1 vccd1 vccd1 _07842_/B sky130_fd_sc_hd__nand2_1
X_08589_ _08593_/C vssd1 vssd1 vccd1 vccd1 _08589_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_36_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10620_ hold39/X _10632_/A vssd1 vssd1 vccd1 vccd1 hold40/A sky130_fd_sc_hd__nor2_1
XFILLER_0_63_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10551_ _10415_/A _10415_/B hold36/X vssd1 vssd1 vccd1 vccd1 _10552_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10482_ _10482_/A _10660_/B vssd1 vssd1 vccd1 vccd1 _10483_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05567__A _08725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07960_ _08061_/B vssd1 vssd1 vccd1 vccd1 _08058_/B sky130_fd_sc_hd__inv_2
X_06911_ _09040_/B _06911_/B vssd1 vssd1 vccd1 vccd1 _06915_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07891_ _09778_/D _07891_/B vssd1 vssd1 vccd1 vccd1 _07896_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06842_ _06842_/A _06842_/B vssd1 vssd1 vccd1 vccd1 _06850_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06398__A _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09630_ _09638_/B _09963_/B vssd1 vssd1 vccd1 vccd1 _09637_/A sky130_fd_sc_hd__nand2_1
X_09561_ _09815_/B _09561_/B vssd1 vssd1 vccd1 vccd1 _09566_/B sky130_fd_sc_hd__nand2_1
X_06773_ _06816_/A _06817_/A vssd1 vssd1 vccd1 vccd1 _06815_/B sky130_fd_sc_hd__nand2_1
X_08512_ _09393_/A _08510_/B _08510_/C vssd1 vssd1 vccd1 vccd1 _08513_/B sky130_fd_sc_hd__o21ai_1
X_05724_ _06162_/C _06162_/B _05723_/Y vssd1 vssd1 vccd1 vccd1 _06121_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_81_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09492_ _09492_/A vssd1 vssd1 vccd1 vccd1 _09494_/B sky130_fd_sc_hd__inv_2
XFILLER_0_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08443_ _08449_/B vssd1 vssd1 vccd1 vccd1 _08450_/B sky130_fd_sc_hd__inv_2
X_05655_ _05697_/B _05695_/A vssd1 vssd1 vccd1 vccd1 _05656_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_73_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05586_ _10201_/A _07646_/D vssd1 vssd1 vccd1 vccd1 _05592_/A sky130_fd_sc_hd__nand2_1
X_08374_ _08374_/A _08374_/B vssd1 vssd1 vccd1 vccd1 _10534_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_73_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07325_ _07756_/A input55/X vssd1 vssd1 vccd1 vccd1 _07516_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07256_ _07579_/A _07579_/B vssd1 vssd1 vccd1 vccd1 _07578_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06207_ _08112_/A _09678_/C vssd1 vssd1 vccd1 vccd1 _06210_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07187_ _07187_/A _07187_/B vssd1 vssd1 vccd1 vccd1 _07187_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07676__B input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06138_ _06323_/B vssd1 vssd1 vccd1 vccd1 _06322_/A sky130_fd_sc_hd__inv_2
X_06069_ _06071_/C vssd1 vssd1 vccd1 vccd1 _06070_/B sky130_fd_sc_hd__inv_2
X_09828_ _09828_/A _09828_/B vssd1 vssd1 vccd1 vccd1 _10353_/B sky130_fd_sc_hd__nand2_2
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09759_ _09759_/A _09759_/B vssd1 vssd1 vccd1 vccd1 _09761_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05940__A _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10603_ _10603_/A _10707_/A _10603_/C vssd1 vssd1 vccd1 vccd1 _10604_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10534_ _10534_/A _10534_/B vssd1 vssd1 vccd1 vccd1 _10535_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10465_ _10467_/C vssd1 vssd1 vccd1 vccd1 _10466_/B sky130_fd_sc_hd__inv_2
X_10396_ _10690_/B _10691_/A _10400_/C vssd1 vssd1 vccd1 vccd1 _10423_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__08698__A _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05440_ _05417_/C _05417_/B _05439_/Y vssd1 vssd1 vccd1 vccd1 _05583_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__10187__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05371_ _08171_/B input8/X vssd1 vssd1 vccd1 vccd1 _05518_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07110_ _07267_/B _07110_/B vssd1 vssd1 vccd1 vccd1 _07595_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08090_ _10493_/B _08086_/Y _10490_/A vssd1 vssd1 vccd1 vccd1 _08244_/A sky130_fd_sc_hd__o21ai_1
X_07041_ _07045_/A _07042_/A vssd1 vssd1 vccd1 vccd1 _07044_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08992_ _08974_/Y _09033_/B _08991_/Y vssd1 vssd1 vccd1 vccd1 _09025_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__08401__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07943_ _07943_/A _07943_/B _07943_/C vssd1 vssd1 vccd1 vccd1 _07956_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09713__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09713__B2 _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ _10284_/B _10158_/A _08897_/B _10157_/A vssd1 vssd1 vccd1 vccd1 _07875_/B
+ sky130_fd_sc_hd__a22o_1
X_09613_ _09613_/A _09613_/B vssd1 vssd1 vccd1 vccd1 _09617_/C sky130_fd_sc_hd__nand2_1
X_06825_ _06825_/A _09036_/B _09036_/C vssd1 vssd1 vccd1 vccd1 _06899_/B sky130_fd_sc_hd__nand3_1
X_09544_ _09544_/A _09544_/B vssd1 vssd1 vccd1 vccd1 _09546_/A sky130_fd_sc_hd__nand2_1
X_06756_ _06758_/A vssd1 vssd1 vccd1 vccd1 _06757_/B sky130_fd_sc_hd__inv_2
X_09475_ _09257_/A _09257_/B _09260_/B vssd1 vssd1 vccd1 vccd1 _09486_/B sky130_fd_sc_hd__o21a_1
XANTENNA__09232__A _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05760__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06687_ _07111_/B _06687_/B vssd1 vssd1 vccd1 vccd1 _07264_/A sky130_fd_sc_hd__nand2_1
X_05707_ _05705_/Y _05667_/B _05706_/Y vssd1 vssd1 vccd1 vccd1 _05839_/A sky130_fd_sc_hd__a21oi_4
X_08426_ _08427_/A _08427_/B vssd1 vssd1 vccd1 vccd1 _08541_/B sky130_fd_sc_hd__or2_1
X_05638_ _05638_/A _05638_/B vssd1 vssd1 vccd1 vccd1 _05640_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05569_ _05571_/A _05571_/B vssd1 vssd1 vccd1 vccd1 _05570_/A sky130_fd_sc_hd__nor2_1
X_08357_ _08357_/A _08357_/B vssd1 vssd1 vccd1 vccd1 _08358_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07308_ _07308_/A _07308_/B _07308_/C vssd1 vssd1 vccd1 vccd1 _07445_/C sky130_fd_sc_hd__nand3_1
X_08288_ _08324_/B vssd1 vssd1 vccd1 vccd1 _08289_/A sky130_fd_sc_hd__inv_2
XANTENNA__05919__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07239_ _07298_/A _07297_/A vssd1 vssd1 vccd1 vccd1 _07239_/Y sky130_fd_sc_hd__nor2_1
X_10250_ _10250_/A _10250_/B vssd1 vssd1 vccd1 vccd1 _10251_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10181_ _10181_/A _10181_/B _10181_/C vssd1 vssd1 vccd1 vccd1 _10238_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_29_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10517_ _10517_/A _10517_/B vssd1 vssd1 vccd1 vccd1 _10638_/A sky130_fd_sc_hd__nand2_2
X_10448_ _10457_/B vssd1 vssd1 vccd1 vccd1 _10449_/B sky130_fd_sc_hd__inv_2
X_10379_ _10379_/A _10705_/B vssd1 vssd1 vccd1 vccd1 _10380_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05845__A _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07590_ _07591_/B _07599_/B vssd1 vssd1 vccd1 vccd1 _07590_/X sky130_fd_sc_hd__and2_1
X_06610_ _06610_/A _06610_/B vssd1 vssd1 vccd1 vccd1 _06613_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06541_ _07043_/B _07042_/A vssd1 vssd1 vccd1 vccd1 _06541_/Y sky130_fd_sc_hd__nor2_1
X_09260_ _09260_/A _09260_/B vssd1 vssd1 vccd1 vccd1 _09264_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06472_ _06605_/A _06610_/A vssd1 vssd1 vccd1 vccd1 _06472_/Y sky130_fd_sc_hd__nor2_1
X_05423_ input62/X vssd1 vssd1 vccd1 vccd1 _07891_/B sky130_fd_sc_hd__clkbuf_8
X_08211_ _08211_/A vssd1 vssd1 vccd1 vccd1 _08213_/A sky130_fd_sc_hd__inv_2
XFILLER_0_55_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09191_ _10158_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _09192_/B sky130_fd_sc_hd__nand2_1
X_08142_ _08141_/B _08142_/B _08142_/C vssd1 vssd1 vccd1 vccd1 _08145_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05354_ _05354_/A vssd1 vssd1 vccd1 vccd1 _05356_/B sky130_fd_sc_hd__inv_2
X_08073_ _08232_/C _08232_/B vssd1 vssd1 vccd1 vccd1 _08233_/A sky130_fd_sc_hd__nand2_1
X_07024_ _07024_/A _07024_/B vssd1 vssd1 vccd1 vccd1 _07026_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06748__A1 _09971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09227__A _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ _08975_/A _08975_/B vssd1 vssd1 vccd1 vccd1 _08976_/B sky130_fd_sc_hd__or2_1
XFILLER_0_11_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _09710_/B _08114_/B vssd1 vssd1 vccd1 vccd1 _07998_/B sky130_fd_sc_hd__nand2_1
Xhold26 hold26/A vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 hold48/A vssd1 vssd1 vccd1 vccd1 hold48/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 hold59/A vssd1 vssd1 vccd1 vccd1 hold59/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08785__B _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07857_ _07857_/A _07857_/B vssd1 vssd1 vccd1 vccd1 _07858_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06586__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06808_ _08975_/A _08822_/A _06808_/C vssd1 vssd1 vccd1 vccd1 _06812_/C sky130_fd_sc_hd__nand3_1
X_07788_ _07792_/B vssd1 vssd1 vccd1 vccd1 _07789_/B sky130_fd_sc_hd__inv_2
X_09527_ _09528_/B _09528_/A vssd1 vssd1 vccd1 vccd1 _09766_/B sky130_fd_sc_hd__or2_1
X_06739_ _06739_/A _08552_/B vssd1 vssd1 vccd1 vccd1 _06740_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05490__A _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09458_ _09458_/A _09458_/B vssd1 vssd1 vccd1 vccd1 _09463_/B sky130_fd_sc_hd__nand2_1
X_08409_ _08413_/C vssd1 vssd1 vccd1 vccd1 _08409_/Y sky130_fd_sc_hd__inv_2
X_09389_ _09390_/B _09390_/A vssd1 vssd1 vccd1 vccd1 _09391_/A sky130_fd_sc_hd__or2_1
X_10302_ _10302_/A vssd1 vssd1 vccd1 vccd1 _10303_/A sky130_fd_sc_hd__inv_2
XFILLER_0_14_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10233_ _10233_/A _10233_/B vssd1 vssd1 vccd1 vccd1 _10235_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09925__A1 _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09925__B2 _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10164_ _10165_/B _10165_/A vssd1 vssd1 vccd1 vccd1 _10168_/B sky130_fd_sc_hd__or2_1
X_10095_ _10569_/C vssd1 vssd1 vccd1 vccd1 _10096_/B sky130_fd_sc_hd__inv_2
XANTENNA__07880__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08695__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10718__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ _09085_/B _08760_/B vssd1 vssd1 vccd1 vccd1 _08809_/B sky130_fd_sc_hd__nand2_1
X_05972_ _05972_/A _05972_/B vssd1 vssd1 vccd1 vccd1 _06796_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07790__A _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08691_ _08833_/B _08691_/B vssd1 vssd1 vccd1 vccd1 _08764_/A sky130_fd_sc_hd__nand2_1
X_07711_ _07822_/B _07823_/B vssd1 vssd1 vccd1 vccd1 _07711_/Y sky130_fd_sc_hd__nor2_1
X_07642_ _07642_/A _07643_/A vssd1 vssd1 vccd1 vccd1 _07653_/A sky130_fd_sc_hd__nand2_1
X_09312_ _09313_/B _09313_/A vssd1 vssd1 vccd1 vccd1 _09312_/Y sky130_fd_sc_hd__nand2_1
X_07573_ _07422_/Y _07835_/C _07423_/Y vssd1 vssd1 vccd1 vccd1 _07577_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__07014__B _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06524_ _10210_/B _10129_/A vssd1 vssd1 vccd1 vccd1 _07005_/B sky130_fd_sc_hd__nand2_1
X_09243_ _09243_/A _09243_/B vssd1 vssd1 vccd1 vccd1 _09244_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_7_132 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06455_ _06457_/A _06455_/B vssd1 vssd1 vccd1 vccd1 _06456_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06853__B _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09174_ _09177_/B _09436_/B vssd1 vssd1 vccd1 vccd1 _09176_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05406_ _05672_/A _05673_/A vssd1 vssd1 vccd1 vccd1 _05406_/Y sky130_fd_sc_hd__nand2_1
X_06386_ _06386_/A _06386_/B vssd1 vssd1 vccd1 vccd1 _06387_/A sky130_fd_sc_hd__nand2_1
X_08125_ _08199_/A _08198_/B _08199_/B vssd1 vssd1 vccd1 vccd1 _08138_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05469__B _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08056_ _08059_/B vssd1 vssd1 vccd1 vccd1 _08060_/A sky130_fd_sc_hd__inv_2
X_07007_ _07012_/B _07012_/C vssd1 vssd1 vccd1 vccd1 _07032_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05485__A _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08958_ _08958_/A _08958_/B vssd1 vssd1 vccd1 vccd1 _09016_/B sky130_fd_sc_hd__nand2_1
X_08889_ _09082_/A vssd1 vssd1 vccd1 vccd1 _08890_/B sky130_fd_sc_hd__inv_2
X_07909_ _07950_/A _07951_/C vssd1 vssd1 vccd1 vccd1 _07910_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09843__B1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10216_ _10208_/A _10216_/B _10216_/C vssd1 vssd1 vccd1 vccd1 _10217_/B sky130_fd_sc_hd__nand3b_1
X_10147_ _10176_/A _10176_/C vssd1 vssd1 vccd1 vccd1 _10175_/A sky130_fd_sc_hd__nand2_1
X_10078_ _10080_/B _10080_/A vssd1 vssd1 vccd1 vccd1 _10079_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06240_ _06240_/A _06240_/B _06240_/C vssd1 vssd1 vccd1 vccd1 _06248_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_80_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06171_ _06171_/A _06171_/B vssd1 vssd1 vccd1 vccd1 _06320_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07785__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09930_ _10170_/B _09930_/B _09930_/C vssd1 vssd1 vccd1 vccd1 _10170_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_68_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09861_ _09861_/A _09861_/B _09861_/C vssd1 vssd1 vccd1 vccd1 _09870_/A sky130_fd_sc_hd__nand3_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09792_ _09793_/B _09793_/A vssd1 vssd1 vccd1 vccd1 _09792_/Y sky130_fd_sc_hd__nand2_1
X_08812_ _08812_/A vssd1 vssd1 vccd1 vccd1 _08813_/B sky130_fd_sc_hd__inv_2
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _08743_/A _08742_/Y vssd1 vssd1 vccd1 vccd1 _08745_/A sky130_fd_sc_hd__nor2b_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05955_ _05955_/A _05956_/A vssd1 vssd1 vccd1 vccd1 _05958_/A sky130_fd_sc_hd__nand2_1
X_08674_ _09699_/A _10188_/B _08674_/C vssd1 vssd1 vccd1 vccd1 _08694_/B sky130_fd_sc_hd__or3_1
X_05886_ _05886_/A _05886_/B vssd1 vssd1 vccd1 vccd1 _05888_/A sky130_fd_sc_hd__nand2_1
X_07625_ _08672_/A _08337_/A vssd1 vssd1 vccd1 vccd1 _07629_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06864__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07556_ _07476_/A _07477_/A _07498_/A vssd1 vssd1 vccd1 vccd1 _07561_/B sky130_fd_sc_hd__o21a_1
XANTENNA__09878__C _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06507_ _06507_/A _06507_/B vssd1 vssd1 vccd1 vccd1 _06508_/B sky130_fd_sc_hd__nand2_1
X_09226_ _09512_/B _09295_/C vssd1 vssd1 vccd1 vccd1 _09294_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07487_ _08897_/B _10156_/A vssd1 vssd1 vccd1 vccd1 _07649_/A sky130_fd_sc_hd__nand2_1
X_06438_ _06438_/A _06438_/B _06438_/C vssd1 vssd1 vccd1 vccd1 _06616_/B sky130_fd_sc_hd__nand3_1
X_09157_ _09159_/A vssd1 vssd1 vccd1 vccd1 _09158_/B sky130_fd_sc_hd__inv_2
X_06369_ _06196_/Y _06369_/B _06369_/C vssd1 vssd1 vccd1 vccd1 _06370_/B sky130_fd_sc_hd__nand3b_1
X_09088_ _08750_/B _08750_/C _08748_/A vssd1 vssd1 vccd1 vccd1 _09109_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_71_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08108_ _08119_/A _08120_/B vssd1 vssd1 vccd1 vccd1 _08118_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08039_ _08041_/A _08041_/B vssd1 vssd1 vccd1 vccd1 _08040_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10001_ _10001_/A _10001_/B _10001_/C vssd1 vssd1 vccd1 vccd1 _10068_/C sky130_fd_sc_hd__nand3_1
XANTENNA__06774__A _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_369 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10696_ hold56/X vssd1 vssd1 vccd1 vccd1 _10726_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10733__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05740_ _06122_/C vssd1 vssd1 vccd1 vccd1 _05741_/C sky130_fd_sc_hd__inv_2
X_05671_ _05673_/A vssd1 vssd1 vccd1 vccd1 _05672_/B sky130_fd_sc_hd__inv_2
XFILLER_0_70_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08390_ input5/X vssd1 vssd1 vccd1 vccd1 _10202_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07410_ _07446_/C vssd1 vssd1 vccd1 vccd1 _07435_/B sky130_fd_sc_hd__inv_2
X_07341_ _07341_/A _07342_/A vssd1 vssd1 vccd1 vccd1 _07344_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07272_ _07274_/A _07274_/B vssd1 vssd1 vccd1 vccd1 _07273_/A sky130_fd_sc_hd__nand2_1
X_09011_ _09028_/C vssd1 vssd1 vccd1 vccd1 _09027_/B sky130_fd_sc_hd__inv_2
X_06223_ _06318_/C vssd1 vssd1 vccd1 vccd1 _06317_/B sky130_fd_sc_hd__inv_2
XFILLER_0_79_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06154_ _06357_/A _06358_/B vssd1 vssd1 vccd1 vccd1 _06154_/Y sky130_fd_sc_hd__nor2_1
X_06085_ _06085_/A _06085_/B vssd1 vssd1 vccd1 vccd1 _06086_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05747__B _06229_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09913_ _09912_/A _09912_/B _09912_/C vssd1 vssd1 vccd1 vccd1 _09914_/B sky130_fd_sc_hd__o21ai_1
X_09844_ _10255_/B _09844_/B vssd1 vssd1 vccd1 vccd1 _09846_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06859__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ _09775_/A _09775_/B _09902_/A vssd1 vssd1 vccd1 vccd1 _09790_/B sky130_fd_sc_hd__nand3_1
X_06987_ _08337_/A _10187_/A vssd1 vssd1 vccd1 vccd1 _07008_/B sky130_fd_sc_hd__nand2_1
X_08726_ _08726_/A _10202_/C _08726_/C vssd1 vssd1 vccd1 vccd1 _08727_/A sky130_fd_sc_hd__nor3_1
X_05938_ _07891_/B _09602_/B vssd1 vssd1 vccd1 vccd1 _05942_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05482__B _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08657_ _09216_/A _08657_/B vssd1 vssd1 vccd1 vccd1 _09281_/A sky130_fd_sc_hd__nand2_1
X_05869_ _06170_/C _06170_/B _05868_/Y vssd1 vssd1 vccd1 vccd1 _06186_/C sky130_fd_sc_hd__a21oi_2
XANTENNA__08793__B _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07608_ _07608_/A _07608_/B _07608_/C vssd1 vssd1 vccd1 vccd1 _07721_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_48_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08588_ _09393_/A _08587_/B _08587_/C vssd1 vssd1 vccd1 vccd1 _08593_/C sky130_fd_sc_hd__o21ai_2
X_07539_ _07659_/B _07659_/C _07538_/Y vssd1 vssd1 vccd1 vccd1 _07656_/A sky130_fd_sc_hd__a21oi_2
X_10550_ _10550_/A _10550_/B vssd1 vssd1 vccd1 vccd1 _10678_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09209_ _09210_/B _09210_/A vssd1 vssd1 vccd1 vccd1 _09209_/Y sky130_fd_sc_hd__nand2_1
X_10481_ _10481_/A _10481_/B vssd1 vssd1 vccd1 vccd1 _10482_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05938__A _07891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10679_ _10679_/A _10682_/A vssd1 vssd1 vccd1 vccd1 _10680_/A sky130_fd_sc_hd__and2_1
XFILLER_0_2_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08224__A _08245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05567__B input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06910_ _06910_/A _06910_/B vssd1 vssd1 vccd1 vccd1 _06911_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07890_ _07975_/A _07975_/B vssd1 vssd1 vccd1 vccd1 _07935_/A sky130_fd_sc_hd__nand2_1
X_06841_ _06841_/A _06841_/B vssd1 vssd1 vccd1 vccd1 _06842_/B sky130_fd_sc_hd__nand2_1
X_09560_ _09815_/A vssd1 vssd1 vccd1 vccd1 _09561_/B sky130_fd_sc_hd__inv_2
X_06772_ _05960_/B _06707_/Y _06708_/Y vssd1 vssd1 vccd1 vccd1 _06817_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09491_ _09491_/A _09491_/B vssd1 vssd1 vccd1 vccd1 _09492_/A sky130_fd_sc_hd__xor2_1
X_08511_ _08511_/A vssd1 vssd1 vccd1 vccd1 _08513_/A sky130_fd_sc_hd__inv_2
X_05723_ _06158_/A _06159_/B vssd1 vssd1 vccd1 vccd1 _05723_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_81_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08442_ _08442_/A _08442_/B vssd1 vssd1 vccd1 vccd1 _08449_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05654_ _05695_/A _05654_/B _05695_/B vssd1 vssd1 vccd1 vccd1 _05697_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_58_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05585_ _06078_/A vssd1 vssd1 vccd1 vccd1 _05622_/A sky130_fd_sc_hd__inv_2
XFILLER_0_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08373_ _08373_/A _08373_/B _08373_/C vssd1 vssd1 vccd1 vccd1 _08374_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_45_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07324_ _07509_/B _07509_/C vssd1 vssd1 vccd1 vccd1 _07508_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07255_ _07255_/A _07255_/B _07255_/C vssd1 vssd1 vccd1 vccd1 _07579_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_33_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09875__D _09875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06206_ _06210_/A vssd1 vssd1 vccd1 vccd1 _06209_/A sky130_fd_sc_hd__inv_2
XFILLER_0_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07186_ _07193_/C _07193_/B vssd1 vssd1 vccd1 vccd1 _07201_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06137_ _08453_/A _07785_/B vssd1 vssd1 vccd1 vccd1 _06323_/B sky130_fd_sc_hd__nand2_1
X_06068_ _06910_/B _06068_/B vssd1 vssd1 vccd1 vccd1 _06071_/C sky130_fd_sc_hd__nand2_1
X_09827_ _09831_/A _09827_/B _10092_/B vssd1 vssd1 vccd1 vccd1 _09828_/B sky130_fd_sc_hd__nand3b_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09758_ _09758_/A _09758_/B vssd1 vssd1 vccd1 vccd1 _09761_/C sky130_fd_sc_hd__nand2_1
X_08709_ _08709_/A _08709_/B vssd1 vssd1 vccd1 vccd1 _08710_/A sky130_fd_sc_hd__nand2_1
X_09689_ _10022_/B _09690_/C _09690_/B vssd1 vssd1 vccd1 vccd1 _09691_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_68_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05940__B _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10602_ hold65/X hold17/X vssd1 vssd1 vccd1 vccd1 _10618_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_36_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10533_ _10534_/B _10534_/A vssd1 vssd1 vccd1 vccd1 _10535_/A sky130_fd_sc_hd__or2_1
XFILLER_0_24_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10464_ _10464_/A _10464_/B vssd1 vssd1 vccd1 vccd1 _10550_/A sky130_fd_sc_hd__nor2_1
X_10395_ _10400_/B _10400_/C vssd1 vssd1 vccd1 vccd1 _10691_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08698__B _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09603__A _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05370_ input59/X vssd1 vssd1 vccd1 vccd1 _08171_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_55_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07040_ _07043_/B vssd1 vssd1 vccd1 vccd1 _07045_/A sky130_fd_sc_hd__inv_2
X_08991_ _09031_/A _09030_/A vssd1 vssd1 vccd1 vccd1 _08991_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08401__B _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07942_ _07942_/A vssd1 vssd1 vccd1 vccd1 _07943_/A sky130_fd_sc_hd__inv_2
XANTENNA__09713__A2 _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07873_ _07873_/A _07873_/B vssd1 vssd1 vccd1 vccd1 _08060_/B sky130_fd_sc_hd__nand2_2
X_09612_ _09613_/B _09613_/A vssd1 vssd1 vccd1 vccd1 _09612_/Y sky130_fd_sc_hd__nor2_1
X_06824_ _06820_/Y _06012_/B _06821_/Y vssd1 vssd1 vccd1 vccd1 _06825_/A sky130_fd_sc_hd__a21oi_1
X_09543_ _09547_/A _09547_/B vssd1 vssd1 vccd1 vccd1 _09799_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06755_ _06755_/A _06755_/B vssd1 vssd1 vccd1 vccd1 _06758_/A sky130_fd_sc_hd__nand2_1
X_09474_ _09474_/A _09692_/A _09474_/C vssd1 vssd1 vccd1 vccd1 _09497_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09232__B _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05760__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06686_ _06687_/B _06686_/B _06940_/A vssd1 vssd1 vccd1 vccd1 _07111_/B sky130_fd_sc_hd__nand3_1
X_05706_ _05706_/A _05706_/B vssd1 vssd1 vccd1 vccd1 _05706_/Y sky130_fd_sc_hd__nor2_1
X_08425_ _10130_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _08427_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05637_ _05639_/A _05639_/B vssd1 vssd1 vccd1 vccd1 _05638_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08356_ _08356_/A _08356_/B _08356_/C _08356_/D vssd1 vssd1 vccd1 vccd1 _08358_/A
+ sky130_fd_sc_hd__and4_1
X_05568_ _08724_/A input36/X vssd1 vssd1 vccd1 vccd1 _05571_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07307_ _07307_/A _07307_/B vssd1 vssd1 vccd1 vccd1 _07445_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05499_ _05894_/B vssd1 vssd1 vccd1 vccd1 _05531_/A sky130_fd_sc_hd__inv_2
X_08287_ _08287_/A _08287_/B vssd1 vssd1 vccd1 vccd1 _08290_/A sky130_fd_sc_hd__nand2_1
X_07238_ _07301_/C vssd1 vssd1 vccd1 vccd1 _07300_/B sky130_fd_sc_hd__inv_2
XFILLER_0_33_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07169_ _07315_/C vssd1 vssd1 vccd1 vccd1 _07314_/B sky130_fd_sc_hd__inv_2
X_10180_ _10180_/A _10180_/B vssd1 vssd1 vccd1 vccd1 _10238_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07878__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10516_ _08360_/A _08361_/B _08360_/C vssd1 vssd1 vccd1 vccd1 _10517_/A sky130_fd_sc_hd__a21o_1
XANTENNA__05398__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10447_ _10453_/B _10447_/B vssd1 vssd1 vccd1 vccd1 _10457_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10378_ _10378_/A _10378_/B vssd1 vssd1 vccd1 vccd1 _10379_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05845__B input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08221__B _08245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06540_ _07044_/C vssd1 vssd1 vccd1 vccd1 _07046_/B sky130_fd_sc_hd__inv_2
X_06471_ _06613_/C vssd1 vssd1 vccd1 vccd1 _06612_/B sky130_fd_sc_hd__inv_2
X_08210_ _08277_/B _08277_/A vssd1 vssd1 vccd1 vccd1 _08214_/A sky130_fd_sc_hd__nor2_1
X_05422_ _05636_/B _05634_/A vssd1 vssd1 vccd1 vccd1 _05422_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_62_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09190_ _10157_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _09192_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_423 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08141_ _08141_/A _08141_/B vssd1 vssd1 vccd1 vccd1 _08145_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05353_ _05353_/A _05353_/B vssd1 vssd1 vccd1 vccd1 _05356_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08072_ _08072_/A _08076_/B _08072_/C vssd1 vssd1 vccd1 vccd1 _08232_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_15_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07023_ _07193_/B _07023_/B vssd1 vssd1 vccd1 vccd1 _07024_/B sky130_fd_sc_hd__nand2_1
X_08974_ _09030_/A _09031_/A vssd1 vssd1 vccd1 vccd1 _08974_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ _07994_/A _07995_/A vssd1 vssd1 vccd1 vccd1 _07999_/B sky130_fd_sc_hd__nand2_1
Xhold27 hold27/A vssd1 vssd1 vccd1 vccd1 hold27/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 hold38/A vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 hold65/A vssd1 vssd1 vccd1 vccd1 hold49/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__05771__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ _07856_/A _07856_/B vssd1 vssd1 vccd1 vccd1 _07857_/A sky130_fd_sc_hd__nand2_1
X_06807_ _08975_/B _06807_/B vssd1 vssd1 vccd1 vccd1 _06812_/B sky130_fd_sc_hd__nand2_1
X_07787_ _08112_/A _07891_/B vssd1 vssd1 vccd1 vccd1 _07792_/B sky130_fd_sc_hd__nand2_1
X_09526_ _09759_/A _09526_/B vssd1 vssd1 vccd1 vccd1 _09528_/A sky130_fd_sc_hd__nand2_1
X_06738_ _06740_/B _06739_/A _08552_/B vssd1 vssd1 vccd1 vccd1 _08552_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__05490__B _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09457_ _09458_/B _09458_/A vssd1 vssd1 vccd1 vccd1 _09463_/A sky130_fd_sc_hd__or2_1
X_08408_ _09912_/A _10188_/C _08407_/C vssd1 vssd1 vccd1 vccd1 _08413_/C sky130_fd_sc_hd__o21ai_2
XFILLER_0_19_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06669_ _06952_/C _06952_/B _06668_/Y vssd1 vssd1 vccd1 vccd1 _06943_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09388_ _09386_/X _09388_/B vssd1 vssd1 vccd1 vccd1 _09390_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_46_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08339_ _10108_/B vssd1 vssd1 vccd1 vccd1 _10113_/A sky130_fd_sc_hd__inv_2
XFILLER_0_34_434 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10301_ _10301_/A _10302_/A vssd1 vssd1 vccd1 vccd1 _10310_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10232_ _10234_/C vssd1 vssd1 vccd1 vccd1 _10233_/B sky130_fd_sc_hd__inv_2
XANTENNA__09925__A2 _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10163_ _10163_/A _10163_/B vssd1 vssd1 vccd1 vccd1 _10165_/A sky130_fd_sc_hd__nand2_1
X_10094_ _10094_/A _10339_/C vssd1 vssd1 vccd1 vccd1 _10569_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08216__B _08245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05971_ _05973_/B vssd1 vssd1 vccd1 vccd1 _05972_/B sky130_fd_sc_hd__inv_2
X_07710_ _07710_/A _07710_/B vssd1 vssd1 vccd1 vccd1 _07824_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_79_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08690_ _08767_/B _08767_/A vssd1 vssd1 vccd1 vccd1 _08833_/B sky130_fd_sc_hd__or2_1
XANTENNA__07790__B _07897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ _07631_/Y _07699_/B _07640_/Y vssd1 vssd1 vccd1 vccd1 _07643_/A sky130_fd_sc_hd__a21oi_2
X_07572_ _07572_/A _07572_/B vssd1 vssd1 vccd1 vccd1 _07577_/B sky130_fd_sc_hd__nand2_1
X_09311_ _09317_/A _09317_/C vssd1 vssd1 vccd1 vccd1 _09316_/A sky130_fd_sc_hd__nand2_1
X_06523_ _07891_/B vssd1 vssd1 vccd1 vccd1 _10129_/A sky130_fd_sc_hd__buf_6
XFILLER_0_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09242_ _09243_/A _09243_/B _09241_/Y vssd1 vssd1 vccd1 vccd1 _09471_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_28_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06454_ _06454_/A vssd1 vssd1 vccd1 vccd1 _06457_/A sky130_fd_sc_hd__inv_2
X_09173_ _09172_/B _09173_/B _09399_/A vssd1 vssd1 vccd1 vccd1 _09436_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_7_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05405_ _05684_/C _05684_/B _05404_/Y vssd1 vssd1 vccd1 vccd1 _05673_/A sky130_fd_sc_hd__a21oi_2
X_06385_ _06567_/B _06567_/C vssd1 vssd1 vccd1 vccd1 _06566_/A sky130_fd_sc_hd__nand2_1
X_08124_ _08198_/A _08199_/C vssd1 vssd1 vccd1 vccd1 _08126_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08055_ _08060_/B vssd1 vssd1 vccd1 vccd1 _08059_/A sky130_fd_sc_hd__inv_2
X_07006_ _07006_/A _07006_/B _07006_/C vssd1 vssd1 vccd1 vccd1 _07012_/B sky130_fd_sc_hd__nand3_1
XANTENNA__05485__B _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08957_ _08959_/C vssd1 vssd1 vccd1 vccd1 _08958_/B sky130_fd_sc_hd__inv_2
X_08888_ _08966_/B _08886_/Y _08887_/Y vssd1 vssd1 vccd1 vccd1 _09082_/A sky130_fd_sc_hd__a21oi_2
X_07908_ _07951_/A _07951_/B vssd1 vssd1 vccd1 vccd1 _07950_/A sky130_fd_sc_hd__nand2_1
X_07839_ _07839_/A _07839_/B vssd1 vssd1 vccd1 vccd1 _07843_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_66_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09843__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09843__B2 _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09509_ _09509_/A vssd1 vssd1 vccd1 vccd1 _09510_/A sky130_fd_sc_hd__inv_2
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09148__A _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10215_ _10208_/Y _10216_/C _10216_/B vssd1 vssd1 vccd1 vccd1 _10217_/A sky130_fd_sc_hd__a21o_1
XANTENNA__07891__A _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ _10146_/A _10146_/B _10146_/C vssd1 vssd1 vccd1 vccd1 _10176_/C sky130_fd_sc_hd__nand3_1
X_10077_ _10077_/A _10077_/B vssd1 vssd1 vccd1 vccd1 _10080_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06170_ _05868_/Y _06170_/B _06170_/C vssd1 vssd1 vccd1 vccd1 _06171_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__07785__B _07785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05586__A _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09860_ _09864_/B _09863_/A vssd1 vssd1 vccd1 vccd1 _09861_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_68_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08897__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _09903_/A _09797_/C vssd1 vssd1 vccd1 vccd1 _10082_/B sky130_fd_sc_hd__nand2_1
X_08811_ _08811_/A _08812_/A vssd1 vssd1 vccd1 vccd1 _08891_/B sky130_fd_sc_hd__nand2_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08742_ _09268_/A _09842_/D _08741_/C vssd1 vssd1 vccd1 vccd1 _08742_/Y sky130_fd_sc_hd__o21ai_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05954_ _05954_/A _05954_/B vssd1 vssd1 vccd1 vccd1 _05956_/A sky130_fd_sc_hd__nand2_1
X_08673_ _10211_/B _10005_/A vssd1 vssd1 vccd1 vccd1 _08674_/C sky130_fd_sc_hd__nand2_1
X_05885_ _05887_/C vssd1 vssd1 vccd1 vccd1 _05886_/B sky130_fd_sc_hd__inv_2
X_07624_ _07675_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _07629_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07555_ _07715_/B _07713_/A vssd1 vssd1 vccd1 vccd1 _07555_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__06864__B _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07486_ _07489_/A _07489_/B vssd1 vssd1 vccd1 vccd1 _07486_/Y sky130_fd_sc_hd__nand2_1
X_06506_ _06506_/A _06506_/B vssd1 vssd1 vccd1 vccd1 _06508_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09225_ _09225_/A _09225_/B vssd1 vssd1 vccd1 vccd1 _09295_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06437_ _06439_/A _06437_/B vssd1 vssd1 vccd1 vccd1 _06438_/B sky130_fd_sc_hd__nand2_1
X_09156_ _09156_/A _09156_/B vssd1 vssd1 vccd1 vccd1 _09159_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06368_ _06196_/Y _06367_/Y _06195_/A vssd1 vssd1 vccd1 vccd1 _06370_/A sky130_fd_sc_hd__o21ai_1
X_09087_ _09126_/A vssd1 vssd1 vccd1 vccd1 _09125_/A sky130_fd_sc_hd__inv_2
X_06299_ _06299_/A _06299_/B vssd1 vssd1 vccd1 vccd1 _06300_/B sky130_fd_sc_hd__or2_1
X_08107_ _08107_/A _08109_/B vssd1 vssd1 vccd1 vccd1 _08119_/A sky130_fd_sc_hd__or2b_1
X_08038_ _08148_/B _08049_/C _08037_/Y vssd1 vssd1 vccd1 vccd1 _08042_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10000_ _10000_/A _10000_/B vssd1 vssd1 vccd1 vccd1 _10068_/A sky130_fd_sc_hd__nand2_1
X_09989_ _09993_/A _09993_/C vssd1 vssd1 vccd1 vccd1 _09992_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06774__B _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10695_ hold55/X _10697_/A vssd1 vssd1 vccd1 vccd1 hold56/A sky130_fd_sc_hd__and2_1
XFILLER_0_81_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10129_ _10129_/A input17/X vssd1 vssd1 vccd1 vccd1 _10131_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06030__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10114__A1 _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05670_ _06248_/C vssd1 vssd1 vccd1 vccd1 _06247_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07340_ _10040_/B _10101_/A vssd1 vssd1 vccd1 vccd1 _07342_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09010_ _09010_/A _09018_/A vssd1 vssd1 vccd1 vccd1 _09028_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_5_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07271_ _07857_/B _07856_/A _07856_/B vssd1 vssd1 vccd1 vccd1 _10431_/C sky130_fd_sc_hd__nand3b_2
XFILLER_0_60_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06222_ _06300_/A _06222_/B vssd1 vssd1 vccd1 vccd1 _06318_/C sky130_fd_sc_hd__nand2_1
X_06153_ _06359_/C vssd1 vssd1 vccd1 vccd1 _06361_/B sky130_fd_sc_hd__inv_2
XFILLER_0_79_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06084_ _06084_/A _06084_/B vssd1 vssd1 vccd1 vccd1 _06085_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06205__A _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09912_ _09912_/A _09912_/B _09912_/C vssd1 vssd1 vccd1 vccd1 _10155_/B sky130_fd_sc_hd__or3_1
X_09843_ input49/X _09710_/B input50/X _10247_/B vssd1 vssd1 vccd1 vccd1 _09844_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06859__B _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _09902_/B _09774_/B vssd1 vssd1 vccd1 vccd1 _09790_/A sky130_fd_sc_hd__nand2_1
X_06986_ _07137_/A _07138_/A vssd1 vssd1 vccd1 vccd1 _07130_/B sky130_fd_sc_hd__nand2_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08725_ _08725_/A _09698_/A vssd1 vssd1 vccd1 vccd1 _08726_/C sky130_fd_sc_hd__nand2_1
X_05937_ _05961_/A _05961_/B vssd1 vssd1 vccd1 vccd1 _05960_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08656_ _09281_/B vssd1 vssd1 vccd1 vccd1 _08658_/A sky130_fd_sc_hd__inv_2
X_05868_ _05868_/A _05868_/B vssd1 vssd1 vccd1 vccd1 _05868_/Y sky130_fd_sc_hd__nor2_1
X_07607_ _07607_/A vssd1 vssd1 vccd1 vccd1 _07608_/C sky130_fd_sc_hd__inv_2
X_08587_ _09393_/A _08587_/B _08587_/C vssd1 vssd1 vccd1 vccd1 _08587_/Y sky130_fd_sc_hd__nor3_1
X_05799_ _05800_/A _05801_/A _05801_/B vssd1 vssd1 vccd1 vccd1 _05836_/A sky130_fd_sc_hd__nand3_1
X_07538_ _07667_/A _07666_/A vssd1 vssd1 vccd1 vccd1 _07538_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_63_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07469_ _07622_/C vssd1 vssd1 vccd1 vccd1 _07471_/B sky130_fd_sc_hd__inv_2
X_09208_ _09214_/A _09441_/A vssd1 vssd1 vccd1 vccd1 _09213_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_294 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10480_ hold33/X vssd1 vssd1 vccd1 vccd1 _10481_/B sky130_fd_sc_hd__inv_2
XANTENNA__05938__B _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ _10112_/A input17/X vssd1 vssd1 vccd1 vccd1 _09140_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09426__A _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__A _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__A _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_0__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _10724_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10678_ _10678_/A _10678_/B vssd1 vssd1 vccd1 vccd1 _10682_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06025__A _08725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05864__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06840_ _06843_/B _06843_/C vssd1 vssd1 vccd1 vccd1 _06842_/A sky130_fd_sc_hd__nand2_1
X_06771_ _08881_/A _06817_/C vssd1 vssd1 vccd1 vccd1 _06816_/A sky130_fd_sc_hd__nand2_1
X_09490_ _09488_/X _09490_/B vssd1 vssd1 vccd1 vccd1 _09491_/B sky130_fd_sc_hd__and2b_1
X_08510_ _09393_/A _08510_/B _08510_/C vssd1 vssd1 vccd1 vccd1 _08511_/A sky130_fd_sc_hd__nor3_1
X_05722_ _06160_/C vssd1 vssd1 vccd1 vccd1 _06162_/B sky130_fd_sc_hd__inv_2
XFILLER_0_81_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08441_ _08466_/B _08466_/C vssd1 vssd1 vccd1 vccd1 _08465_/A sky130_fd_sc_hd__nand2_1
X_05653_ _05653_/A _05653_/B vssd1 vssd1 vccd1 vccd1 _05706_/B sky130_fd_sc_hd__nand2_1
X_08372_ _08372_/A _08372_/B vssd1 vssd1 vccd1 vccd1 _08374_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05584_ _05582_/Y _05457_/B _05583_/Y vssd1 vssd1 vccd1 vccd1 _06078_/A sky130_fd_sc_hd__a21oi_4
X_07323_ _07323_/A _07323_/B _07323_/C vssd1 vssd1 vccd1 vccd1 _07509_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_5_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07254_ _07254_/A _07254_/B vssd1 vssd1 vccd1 vccd1 _07579_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06205_ _09778_/D _10005_/A vssd1 vssd1 vccd1 vccd1 _06210_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07185_ _07185_/A _07185_/B _07185_/C vssd1 vssd1 vccd1 vccd1 _07193_/C sky130_fd_sc_hd__nand3_1
X_06136_ _06322_/B vssd1 vssd1 vccd1 vccd1 _06323_/A sky130_fd_sc_hd__inv_2
X_06067_ _06067_/A _06067_/B vssd1 vssd1 vccd1 vccd1 _06068_/B sky130_fd_sc_hd__nand2_1
X_09826_ _09831_/B _09831_/A vssd1 vssd1 vccd1 vccd1 _09828_/A sky130_fd_sc_hd__nand2_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09757_ _09757_/A vssd1 vssd1 vccd1 vccd1 _09859_/B sky130_fd_sc_hd__inv_2
X_06969_ _06969_/A _06969_/B _06969_/C vssd1 vssd1 vccd1 vccd1 _07127_/C sky130_fd_sc_hd__nand3_1
X_08708_ _08710_/B _08709_/A _08709_/B vssd1 vssd1 vccd1 vccd1 _08714_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_68_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09688_ _09456_/B _10201_/A _10187_/B _09454_/X vssd1 vssd1 vccd1 vccd1 _09690_/B
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08639_ _08633_/Y _08639_/B _08639_/C vssd1 vssd1 vccd1 vccd1 _08643_/C sky130_fd_sc_hd__nand3b_1
XANTENNA__08309__B _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10601_ _10601_/A vssd1 vssd1 vccd1 vccd1 _10734_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10532_ _10532_/A _10532_/B vssd1 vssd1 vccd1 vccd1 _10534_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10463_ _10548_/A _10463_/B vssd1 vssd1 vccd1 vccd1 _10464_/B sky130_fd_sc_hd__nor2_1
X_10394_ _10394_/A _10394_/B _10725_/Q vssd1 vssd1 vccd1 vccd1 _10400_/C sky130_fd_sc_hd__nand3_1
XANTENNA__09603__B _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08990_ _09034_/C vssd1 vssd1 vccd1 vccd1 _09033_/B sky130_fd_sc_hd__inv_2
XANTENNA__05594__A _08672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07941_ _07941_/A _07942_/A vssd1 vssd1 vccd1 vccd1 _07956_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10005__A _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ _07872_/A _07872_/B _07872_/C vssd1 vssd1 vccd1 vccd1 _07873_/B sky130_fd_sc_hd__nand3_1
X_06823_ _06823_/A _09036_/A vssd1 vssd1 vccd1 vccd1 _06899_/A sky130_fd_sc_hd__nand2_1
X_09611_ _09611_/A _09611_/B vssd1 vssd1 vccd1 vccd1 _09613_/A sky130_fd_sc_hd__and2_1
X_09542_ _09541_/B _09542_/B _09542_/C vssd1 vssd1 vccd1 vccd1 _09547_/B sky130_fd_sc_hd__nand3b_1
X_06754_ _06758_/B _08435_/A vssd1 vssd1 vccd1 vccd1 _06757_/A sky130_fd_sc_hd__nand2_1
X_05705_ _05706_/B _05706_/A vssd1 vssd1 vccd1 vccd1 _05705_/Y sky130_fd_sc_hd__nand2_1
X_09473_ _09473_/A vssd1 vssd1 vccd1 vccd1 _09474_/C sky130_fd_sc_hd__inv_2
X_06685_ _06685_/A _06685_/B vssd1 vssd1 vccd1 vccd1 _06940_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08424_ _10129_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _08427_/A sky130_fd_sc_hd__nand2_1
X_05636_ _05636_/A _05636_/B vssd1 vssd1 vccd1 vccd1 _05639_/B sky130_fd_sc_hd__nand2_1
X_05567_ _08725_/A input37/X vssd1 vssd1 vccd1 vccd1 _05571_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08355_ _08355_/A _08355_/B vssd1 vssd1 vccd1 vccd1 _08356_/D sky130_fd_sc_hd__nand2_1
XFILLER_0_18_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05769__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07306_ _07308_/A _07308_/B vssd1 vssd1 vccd1 vccd1 _07307_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05498_ _05498_/A _05498_/B vssd1 vssd1 vccd1 vccd1 _05894_/B sky130_fd_sc_hd__nand2_1
X_08286_ _08330_/B _08366_/B vssd1 vssd1 vccd1 vccd1 _08329_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07237_ _07237_/A _07237_/B vssd1 vssd1 vccd1 vccd1 _07301_/C sky130_fd_sc_hd__nand2_1
X_07168_ _07168_/A _07168_/B vssd1 vssd1 vccd1 vccd1 _07315_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06119_ _06179_/B _06179_/C vssd1 vssd1 vccd1 vccd1 _06299_/B sky130_fd_sc_hd__nand2_1
X_07099_ _07099_/A _07243_/A vssd1 vssd1 vccd1 vccd1 _07101_/A sky130_fd_sc_hd__nand2_1
X_09809_ _09813_/B _09836_/A vssd1 vssd1 vccd1 vccd1 _09812_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07878__B _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10515_ hold50/X vssd1 vssd1 vccd1 vccd1 _10638_/B sky130_fd_sc_hd__inv_2
XFILLER_0_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05398__B _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10446_ _10446_/A _10446_/B vssd1 vssd1 vccd1 vccd1 _10449_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10377_ hold61/X vssd1 vssd1 vccd1 vccd1 _10378_/B sky130_fd_sc_hd__inv_2
XANTENNA__05845__C _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06470_ _06470_/A _06470_/B vssd1 vssd1 vccd1 vccd1 _06613_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_7_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05421_ _05406_/Y _05675_/B _05420_/Y vssd1 vssd1 vccd1 vccd1 _05634_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__05589__A _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08140_ _08142_/B _08142_/C vssd1 vssd1 vccd1 vccd1 _08141_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05352_ _05352_/A _05352_/B _05354_/A vssd1 vssd1 vccd1 vccd1 _05368_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_43_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08071_ _08079_/B _08079_/A vssd1 vssd1 vccd1 vccd1 _08232_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_70_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07022_ _07023_/B _07022_/B _07022_/C vssd1 vssd1 vccd1 vccd1 _07193_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_11_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08973_ _09030_/B vssd1 vssd1 vccd1 vccd1 _09031_/A sky130_fd_sc_hd__inv_2
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _09840_/B _08574_/A vssd1 vssd1 vccd1 vccd1 _07995_/A sky130_fd_sc_hd__nand2_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_07855_ _07855_/A _07855_/B vssd1 vssd1 vccd1 vccd1 _10426_/C sky130_fd_sc_hd__nor2_1
X_06806_ _08975_/A vssd1 vssd1 vccd1 vccd1 _06807_/B sky130_fd_sc_hd__inv_2
XANTENNA__05771__B _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07786_ _07792_/A vssd1 vssd1 vccd1 vccd1 _07789_/A sky130_fd_sc_hd__inv_2
X_09525_ _09525_/A _09525_/B vssd1 vssd1 vccd1 vccd1 _09526_/B sky130_fd_sc_hd__nand2_1
X_06737_ _06737_/A _06737_/B _08478_/A vssd1 vssd1 vccd1 vccd1 _08552_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_78_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09456_ _09454_/X _09456_/B vssd1 vssd1 vccd1 vccd1 _09458_/A sky130_fd_sc_hd__nand2b_1
X_06668_ _06954_/A _06953_/A vssd1 vssd1 vccd1 vccd1 _06668_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_38_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08407_ _09912_/A _10188_/C _08407_/C vssd1 vssd1 vccd1 vccd1 _08407_/Y sky130_fd_sc_hd__nor3_1
X_05619_ _05619_/A _05619_/B vssd1 vssd1 vccd1 vccd1 _05623_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_81_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09387_ _10130_/A _10158_/B _10129_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _09388_/B
+ sky130_fd_sc_hd__a22o_1
X_06599_ _06601_/B _06602_/B _06602_/C vssd1 vssd1 vccd1 vccd1 _06600_/A sky130_fd_sc_hd__nand3_1
X_08338_ _08897_/B vssd1 vssd1 vccd1 vccd1 _09782_/B sky130_fd_sc_hd__inv_2
XFILLER_0_61_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08269_ _08269_/A _08269_/B vssd1 vssd1 vccd1 vccd1 _08269_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_34_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10300_ _10300_/A _10300_/B vssd1 vssd1 vccd1 vccd1 _10302_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10231_ _10231_/A _10231_/B vssd1 vssd1 vccd1 vccd1 _10234_/C sky130_fd_sc_hd__nor2_1
X_10162_ _10162_/A _10161_/A vssd1 vssd1 vccd1 vccd1 _10163_/B sky130_fd_sc_hd__or2b_1
X_10093_ _10092_/B _10334_/B _10093_/C vssd1 vssd1 vccd1 vccd1 _10339_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_69_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10727__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10429_ _10431_/B vssd1 vssd1 vccd1 vccd1 _10430_/B sky130_fd_sc_hd__inv_2
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05970_ _10158_/A _10004_/A vssd1 vssd1 vccd1 vccd1 _05973_/B sky130_fd_sc_hd__nand2_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05872__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07640_ _07697_/A _07696_/A vssd1 vssd1 vccd1 vccd1 _07640_/Y sky130_fd_sc_hd__nor2_1
X_07571_ _07839_/B _07839_/A vssd1 vssd1 vccd1 vccd1 _07847_/B sky130_fd_sc_hd__nor2_1
X_09310_ _09310_/A _09310_/B _09581_/C vssd1 vssd1 vccd1 vccd1 _09317_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_75_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06522_ _07004_/B vssd1 vssd1 vccd1 vccd1 _07005_/A sky130_fd_sc_hd__inv_2
XFILLER_0_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09241_ _09244_/A _09244_/C vssd1 vssd1 vccd1 vccd1 _09241_/Y sky130_fd_sc_hd__nand2_1
X_06453_ _06457_/B _06454_/A vssd1 vssd1 vccd1 vccd1 _06456_/A sky130_fd_sc_hd__nand2_1
X_09172_ _09172_/A _09172_/B vssd1 vssd1 vccd1 vccd1 _09177_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_16_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05404_ _05680_/A _05681_/B vssd1 vssd1 vccd1 vccd1 _05404_/Y sky130_fd_sc_hd__nor2_1
X_06384_ _06384_/A _06384_/B vssd1 vssd1 vccd1 vccd1 _06567_/B sky130_fd_sc_hd__nand2_1
X_08123_ _08199_/A _08199_/B vssd1 vssd1 vccd1 vccd1 _08198_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08054_ _08153_/B _08091_/B vssd1 vssd1 vccd1 vccd1 _08218_/A sky130_fd_sc_hd__nand2_2
XANTENNA__08423__A _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07005_ _07005_/A _07005_/B vssd1 vssd1 vccd1 vccd1 _07006_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_24_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08956_ _08956_/A _09080_/A vssd1 vssd1 vccd1 vccd1 _08959_/C sky130_fd_sc_hd__nand2_1
X_08887_ _08964_/A _08963_/A vssd1 vssd1 vccd1 vccd1 _08887_/Y sky130_fd_sc_hd__nor2_1
X_07907_ _08041_/C vssd1 vssd1 vccd1 vccd1 _08040_/B sky130_fd_sc_hd__inv_2
X_07838_ _07838_/A _07838_/B vssd1 vssd1 vccd1 vccd1 _07850_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09508_ _09508_/A _09509_/A vssd1 vssd1 vccd1 vccd1 _09514_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07769_ _07769_/A _07769_/B vssd1 vssd1 vccd1 vccd1 _07770_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09843__A2 _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _09439_/A _09615_/A _09725_/A vssd1 vssd1 vccd1 vccd1 _09443_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_54_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09429__A _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10214_ _10214_/A _10214_/B vssd1 vssd1 vccd1 vccd1 _10216_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07891__B _07891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ _10145_/A _10145_/B vssd1 vssd1 vccd1 vccd1 _10176_/A sky130_fd_sc_hd__nand2_1
X_10076_ _10076_/A _10076_/B vssd1 vssd1 vccd1 vccd1 _10077_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09164__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10103__A _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05586__B _07646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08897__B _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08810_ _08810_/A _08810_/B vssd1 vssd1 vccd1 vccd1 _08812_/A sky130_fd_sc_hd__nand2_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09790_ _09790_/A _09790_/B _09790_/C vssd1 vssd1 vccd1 vccd1 _09797_/C sky130_fd_sc_hd__nand3_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08741_ _09268_/A _09842_/D _08741_/C vssd1 vssd1 vccd1 vccd1 _08743_/A sky130_fd_sc_hd__nor3_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05953_ _05957_/A _05957_/B vssd1 vssd1 vccd1 vccd1 _05955_/A sky130_fd_sc_hd__nand2_1
X_08672_ _08672_/A vssd1 vssd1 vccd1 vccd1 _09699_/A sky130_fd_sc_hd__inv_2
X_05884_ _06117_/B _05882_/Y _05883_/Y vssd1 vssd1 vccd1 vccd1 _05887_/C sky130_fd_sc_hd__a21oi_1
X_07623_ _07697_/B _07697_/C vssd1 vssd1 vccd1 vccd1 _07696_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07554_ _07612_/B _07612_/C _07553_/Y vssd1 vssd1 vccd1 vccd1 _07713_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_75_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07485_ _08112_/A input64/X vssd1 vssd1 vccd1 vccd1 _07489_/B sky130_fd_sc_hd__nand2_1
X_06505_ _06659_/B _06659_/C vssd1 vssd1 vccd1 vccd1 _06661_/A sky130_fd_sc_hd__nand2_1
X_09224_ _08666_/B _08666_/C _09134_/B vssd1 vssd1 vccd1 vccd1 _09225_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_8_443 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06436_ _06436_/A vssd1 vssd1 vccd1 vccd1 _06439_/A sky130_fd_sc_hd__inv_2
XFILLER_0_8_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09155_ _09159_/B _09381_/A vssd1 vssd1 vccd1 vccd1 _09158_/A sky130_fd_sc_hd__nand2_1
X_06367_ _06369_/C vssd1 vssd1 vccd1 vccd1 _06367_/Y sky130_fd_sc_hd__inv_2
X_09086_ _09084_/Y _08808_/B _09085_/Y vssd1 vssd1 vccd1 vccd1 _09126_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08106_ _08184_/B vssd1 vssd1 vccd1 vccd1 _08185_/C sky130_fd_sc_hd__inv_2
XFILLER_0_16_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06298_ _06495_/B _06494_/A vssd1 vssd1 vccd1 vccd1 _06298_/Y sky130_fd_sc_hd__nand2_1
X_08037_ _08037_/A _08037_/B vssd1 vssd1 vccd1 vccd1 _08037_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09988_ _09988_/A _09988_/B _09988_/C vssd1 vssd1 vccd1 vccd1 _09993_/C sky130_fd_sc_hd__nand3_1
X_08939_ _08998_/B _08939_/B vssd1 vssd1 vccd1 vccd1 _08942_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09712__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10694_ _10694_/A _10694_/B vssd1 vssd1 vccd1 vccd1 _10697_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05687__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10128_ _10128_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _10132_/A sky130_fd_sc_hd__nand2_1
X_10059_ _10059_/A _10059_/B vssd1 vssd1 vccd1 vccd1 _10061_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09622__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07270_ _07270_/A _07274_/C _07270_/C vssd1 vssd1 vccd1 vccd1 _07856_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_72_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06221_ _06220_/B _06221_/B _06221_/C vssd1 vssd1 vccd1 vccd1 _06222_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_5_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06152_ _07675_/A input35/X vssd1 vssd1 vccd1 vccd1 _06359_/C sky130_fd_sc_hd__nand2_1
X_06083_ _06085_/B _06084_/A _06084_/B vssd1 vssd1 vccd1 vccd1 _06086_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_13_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09911_ _10157_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _09912_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06205__B _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09842_ _10248_/A _10248_/C _10248_/D _09842_/D vssd1 vssd1 vccd1 vccd1 _10255_/B
+ sky130_fd_sc_hd__or4_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _09902_/A vssd1 vssd1 vccd1 vccd1 _09774_/B sky130_fd_sc_hd__inv_2
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08724_ _08724_/A vssd1 vssd1 vccd1 vccd1 _08726_/A sky130_fd_sc_hd__inv_2
X_06985_ _07147_/C _07147_/B _06984_/Y vssd1 vssd1 vccd1 vccd1 _07138_/A sky130_fd_sc_hd__a21oi_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05936_ _06708_/A _05936_/B _05936_/C vssd1 vssd1 vccd1 vccd1 _05961_/B sky130_fd_sc_hd__nand3_1
X_08655_ _09281_/B _08657_/B _09216_/A vssd1 vssd1 vccd1 vccd1 _08662_/B sky130_fd_sc_hd__nand3_1
X_05867_ _05867_/A vssd1 vssd1 vccd1 vccd1 _06170_/B sky130_fd_sc_hd__inv_2
X_07606_ _07606_/A _07607_/A vssd1 vssd1 vccd1 vccd1 _07721_/B sky130_fd_sc_hd__nand2_1
X_08586_ _10103_/B _10158_/B vssd1 vssd1 vccd1 vccd1 _08587_/C sky130_fd_sc_hd__nand2_1
X_05798_ _05798_/A _05798_/B _05798_/C vssd1 vssd1 vccd1 vccd1 _05801_/B sky130_fd_sc_hd__nand3_1
X_07537_ _07668_/C vssd1 vssd1 vccd1 vccd1 _07659_/C sky130_fd_sc_hd__inv_2
XANTENNA__07052__A _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07468_ _09517_/D _07897_/B vssd1 vssd1 vccd1 vccd1 _07622_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_29_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_338 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09207_ _09206_/B _09207_/B _09441_/B vssd1 vssd1 vccd1 vccd1 _09441_/A sky130_fd_sc_hd__nand3b_1
X_07399_ _07405_/B _07405_/C vssd1 vssd1 vccd1 vccd1 _07403_/A sky130_fd_sc_hd__nand2_1
X_06419_ _06676_/B _06676_/C vssd1 vssd1 vccd1 vccd1 _06675_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09138_ _10108_/B input18/X vssd1 vssd1 vccd1 vccd1 _09140_/A sky130_fd_sc_hd__nand2_1
X_09069_ _09069_/A _09069_/B _09069_/C vssd1 vssd1 vccd1 vccd1 _09072_/C sky130_fd_sc_hd__nand3_1
XANTENNA__09426__B _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05970__A _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__B _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09161__B _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07897__A _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10677_ _10678_/B _10678_/A vssd1 vssd1 vccd1 vccd1 _10679_/A sky130_fd_sc_hd__or2_1
XANTENNA__09973__A1 _09971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06025__B _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05864__B _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09489__B1 _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ _06816_/B _08881_/A _06817_/C vssd1 vssd1 vccd1 vccd1 _08972_/B sky130_fd_sc_hd__nand3_1
X_05721_ _08725_/A input35/X vssd1 vssd1 vccd1 vccd1 _06160_/C sky130_fd_sc_hd__nand2_1
X_08440_ _08660_/A _08440_/B _08757_/A vssd1 vssd1 vccd1 vccd1 _08466_/C sky130_fd_sc_hd__nand3_1
X_05652_ _05706_/A _05653_/B _05653_/A vssd1 vssd1 vccd1 vccd1 _05668_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_73_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08371_ _08373_/A vssd1 vssd1 vccd1 vccd1 _08372_/B sky130_fd_sc_hd__inv_2
XFILLER_0_18_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05583_ _05583_/A _05583_/B vssd1 vssd1 vccd1 vccd1 _05583_/Y sky130_fd_sc_hd__nor2_1
X_07322_ _07322_/A _07322_/B vssd1 vssd1 vccd1 vccd1 _07323_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07253_ _07255_/A vssd1 vssd1 vccd1 vccd1 _07254_/B sky130_fd_sc_hd__inv_2
X_07184_ _07184_/A _07184_/B vssd1 vssd1 vccd1 vccd1 _07185_/B sky130_fd_sc_hd__nand2_1
X_06204_ input1/X _10187_/B vssd1 vssd1 vccd1 vccd1 _06387_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_53_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06135_ _08672_/A _07891_/B vssd1 vssd1 vccd1 vccd1 _06322_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06066_ _06066_/A vssd1 vssd1 vccd1 vccd1 _06910_/B sky130_fd_sc_hd__inv_2
XFILLER_0_41_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09825_ _09827_/B _10092_/B vssd1 vssd1 vccd1 vccd1 _09831_/B sky130_fd_sc_hd__nand2_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09756_ _09758_/B _09758_/A vssd1 vssd1 vccd1 vccd1 _09757_/A sky130_fd_sc_hd__nor2_1
X_06968_ _06968_/A _06968_/B _06968_/C vssd1 vssd1 vccd1 vccd1 _06969_/B sky130_fd_sc_hd__nand3_1
X_08707_ _08707_/A _09229_/A _09247_/A vssd1 vssd1 vccd1 vccd1 _08709_/B sky130_fd_sc_hd__nand3_1
X_09687_ _09687_/A _09687_/B vssd1 vssd1 vccd1 vccd1 _09690_/C sky130_fd_sc_hd__nand2_1
X_05919_ _08171_/B _10150_/B vssd1 vssd1 vccd1 vccd1 _05924_/A sky130_fd_sc_hd__nand2_1
X_08638_ _08638_/A vssd1 vssd1 vccd1 vccd1 _08639_/B sky130_fd_sc_hd__inv_2
X_06899_ _06899_/A _06899_/B _06899_/C vssd1 vssd1 vccd1 vccd1 _06906_/C sky130_fd_sc_hd__nand3_1
XANTENNA__10201__A _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08309__C _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08569_ _08964_/C _08868_/B vssd1 vssd1 vccd1 vccd1 _08667_/A sky130_fd_sc_hd__nand2_1
X_10600_ _10600_/A _10600_/B vssd1 vssd1 vccd1 vccd1 _10601_/A sky130_fd_sc_hd__and2_1
X_10531_ hold58/X vssd1 vssd1 vccd1 vccd1 _10537_/B sky130_fd_sc_hd__inv_2
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10462_ _10667_/A _10459_/Y _10461_/Y vssd1 vssd1 vccd1 vccd1 _10463_/B sky130_fd_sc_hd__a21oi_1
X_10393_ _10393_/A _10393_/B vssd1 vssd1 vccd1 vccd1 _10400_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09603__C _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10729_ _10733_/CLK hold42/X fanout98/X vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07940_ _07943_/B _07943_/C vssd1 vssd1 vccd1 vccd1 _07941_/A sky130_fd_sc_hd__nand2_1
X_07871_ _07871_/A _07871_/B vssd1 vssd1 vccd1 vccd1 _07872_/A sky130_fd_sc_hd__nand2_1
X_09610_ _09610_/A _09936_/A vssd1 vssd1 vccd1 vccd1 _09613_/B sky130_fd_sc_hd__nand2_1
X_06822_ _06820_/Y _06012_/B _06821_/Y vssd1 vssd1 vccd1 vccd1 _09036_/A sky130_fd_sc_hd__a21o_1
X_09541_ _09541_/A _09541_/B vssd1 vssd1 vccd1 vccd1 _09547_/A sky130_fd_sc_hd__nand2_1
X_06753_ _08435_/B _06753_/B _06753_/C vssd1 vssd1 vccd1 vccd1 _08435_/A sky130_fd_sc_hd__nand3_1
X_05704_ _06229_/B _06228_/B vssd1 vssd1 vccd1 vccd1 _06227_/C sky130_fd_sc_hd__nand2_1
X_09472_ _09472_/A _09473_/A vssd1 vssd1 vccd1 vccd1 _09497_/A sky130_fd_sc_hd__nand2_1
X_06684_ _06939_/A _06938_/A vssd1 vssd1 vccd1 vccd1 _06686_/B sky130_fd_sc_hd__nand2_1
X_08423_ _10128_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _08430_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_46_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05635_ _05406_/Y _05675_/B _05420_/Y vssd1 vssd1 vccd1 vccd1 _05636_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_58_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05566_ input30/X vssd1 vssd1 vccd1 vccd1 _08725_/A sky130_fd_sc_hd__clkbuf_8
X_08354_ _08354_/A _08354_/B vssd1 vssd1 vccd1 vccd1 _08356_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09634__B1 _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05769__B _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07305_ _07305_/A _07305_/B vssd1 vssd1 vccd1 vccd1 _07308_/B sky130_fd_sc_hd__nand2_1
X_05497_ _05497_/A _05497_/B _05497_/C vssd1 vssd1 vccd1 vccd1 _05498_/B sky130_fd_sc_hd__nand3_1
X_08285_ _08285_/A _08285_/B _08363_/B vssd1 vssd1 vccd1 vccd1 _08366_/B sky130_fd_sc_hd__nand3_4
X_07236_ _07235_/B _07236_/B _07236_/C vssd1 vssd1 vccd1 vccd1 _07237_/B sky130_fd_sc_hd__nand3b_1
X_07167_ _07167_/A _07167_/B _07167_/C vssd1 vssd1 vccd1 vccd1 _07168_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06118_ _06118_/A _06118_/B _06118_/C vssd1 vssd1 vccd1 vccd1 _06179_/C sky130_fd_sc_hd__nand3_1
X_07098_ _07415_/A _07242_/A vssd1 vssd1 vccd1 vccd1 _07243_/A sky130_fd_sc_hd__or2_1
X_06049_ _09517_/C vssd1 vssd1 vccd1 vccd1 _10276_/B sky130_fd_sc_hd__inv_2
X_09808_ _09808_/A _09808_/B _09836_/B vssd1 vssd1 vccd1 vccd1 _09836_/A sky130_fd_sc_hd__nand3_1
X_09739_ _09739_/A _09739_/B vssd1 vssd1 vccd1 vccd1 _09742_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08336__A _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10514_ _10514_/A _10514_/B vssd1 vssd1 vccd1 vccd1 _10641_/A sky130_fd_sc_hd__nand2_1
X_10445_ _10466_/A _10445_/B vssd1 vssd1 vccd1 vccd1 _10446_/A sky130_fd_sc_hd__nand2_1
X_10376_ _10376_/A _10376_/B vssd1 vssd1 vccd1 vccd1 _10378_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05845__D _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08364__B1 _08366_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05420_ _05673_/A _05672_/A vssd1 vssd1 vccd1 vccd1 _05420_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07150__A _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05351_ _08114_/B _10151_/B vssd1 vssd1 vccd1 vccd1 _05354_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05589__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08070_ _08072_/A vssd1 vssd1 vccd1 vccd1 _08079_/A sky130_fd_sc_hd__inv_2
XFILLER_0_15_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07021_ _07183_/B _07184_/B vssd1 vssd1 vccd1 vccd1 _07022_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_51_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_355 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08972_ _09036_/B _08972_/B vssd1 vssd1 vccd1 vccd1 _09030_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
X_07923_ _10247_/B _08573_/A vssd1 vssd1 vccd1 vccd1 _07994_/A sky130_fd_sc_hd__nand2_1
X_07854_ _08386_/C _10446_/B vssd1 vssd1 vccd1 vccd1 _07855_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06805_ _06803_/Y _05956_/A _06804_/Y vssd1 vssd1 vccd1 vccd1 _08975_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__07325__A _07756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07785_ _09517_/D _07785_/B vssd1 vssd1 vccd1 vccd1 _07792_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09524_ _09524_/A _09524_/B vssd1 vssd1 vccd1 vccd1 _09759_/A sky130_fd_sc_hd__nand2_1
X_06736_ _06736_/A _06736_/B vssd1 vssd1 vccd1 vccd1 _06739_/A sky130_fd_sc_hd__nand2_1
X_09455_ _09677_/A _10005_/A _10004_/A _09678_/C vssd1 vssd1 vccd1 vccd1 _09456_/B
+ sky130_fd_sc_hd__a22o_1
X_06667_ _06955_/C vssd1 vssd1 vccd1 vccd1 _06952_/B sky130_fd_sc_hd__inv_2
XFILLER_0_38_208 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08406_ _10157_/A _09602_/B vssd1 vssd1 vccd1 vccd1 _08407_/C sky130_fd_sc_hd__nand2_1
X_05618_ _05620_/C vssd1 vssd1 vccd1 vccd1 _05619_/B sky130_fd_sc_hd__inv_2
X_09386_ _10130_/A _10129_/A _10157_/B _10158_/B vssd1 vssd1 vccd1 vccd1 _09386_/X
+ sky130_fd_sc_hd__and4_1
XFILLER_0_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06598_ _06463_/Y _06612_/B _06472_/Y vssd1 vssd1 vccd1 vccd1 _06601_/B sky130_fd_sc_hd__a21o_1
X_05549_ _08672_/A _07646_/D vssd1 vssd1 vccd1 vccd1 _05600_/A sky130_fd_sc_hd__nand2_1
X_08337_ _08337_/A vssd1 vssd1 vccd1 vccd1 _09393_/A sky130_fd_sc_hd__inv_2
XFILLER_0_34_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08268_ _08269_/B _08269_/A vssd1 vssd1 vccd1 vccd1 _08297_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ _07222_/A _07222_/B vssd1 vssd1 vccd1 vccd1 _07377_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_21_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10230_ _10230_/A vssd1 vssd1 vccd1 vccd1 _10231_/B sky130_fd_sc_hd__inv_2
XFILLER_0_14_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08199_ _08199_/A _08199_/B _08199_/C vssd1 vssd1 vccd1 vccd1 _08200_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06404__A _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10161_ _10161_/A _10162_/A vssd1 vssd1 vccd1 vccd1 _10163_/A sky130_fd_sc_hd__or2b_1
X_10092_ _10092_/A _10092_/B vssd1 vssd1 vccd1 vccd1 _10094_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08649__A1 _09201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10428_ _10438_/A _10431_/C vssd1 vssd1 vccd1 vccd1 _10430_/A sky130_fd_sc_hd__nand2_1
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10359_ _10359_/A vssd1 vssd1 vccd1 vccd1 _10360_/B sky130_fd_sc_hd__inv_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05872__B _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07570_ _07570_/A _07570_/B vssd1 vssd1 vccd1 vccd1 _07839_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09360__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06521_ _10211_/B _10130_/A vssd1 vssd1 vccd1 vccd1 _07004_/B sky130_fd_sc_hd__nand2_1
X_09240_ _09469_/A _09469_/B _09470_/A vssd1 vssd1 vccd1 vccd1 _09244_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06452_ _06455_/B vssd1 vssd1 vccd1 vccd1 _06457_/B sky130_fd_sc_hd__inv_2
X_09171_ _08593_/C _08593_/B _08587_/Y vssd1 vssd1 vccd1 vccd1 _09172_/B sky130_fd_sc_hd__a21oi_1
X_05403_ _05682_/C vssd1 vssd1 vccd1 vccd1 _05684_/B sky130_fd_sc_hd__inv_2
X_06383_ _06383_/A vssd1 vssd1 vccd1 vccd1 _06384_/B sky130_fd_sc_hd__inv_2
XFILLER_0_43_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08122_ _08185_/C _08185_/B _08197_/B vssd1 vssd1 vccd1 vccd1 _08135_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08053_ _08091_/A _08091_/B _08092_/A vssd1 vssd1 vccd1 vccd1 _08153_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08423__B _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07004_ _07004_/A _07004_/B vssd1 vssd1 vccd1 vccd1 _07006_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06224__A _06229_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ _09002_/B _09080_/B _08955_/C vssd1 vssd1 vccd1 vccd1 _09080_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_11_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07906_ _08061_/B _07906_/B vssd1 vssd1 vccd1 vccd1 _08041_/C sky130_fd_sc_hd__nand2_1
X_08886_ _08963_/A _08964_/A vssd1 vssd1 vccd1 vccd1 _08886_/Y sky130_fd_sc_hd__nand2_1
X_07837_ _07560_/Y _07607_/A _07562_/Y vssd1 vssd1 vccd1 vccd1 _07838_/B sky130_fd_sc_hd__a21o_1
X_07768_ _07768_/A _07768_/B vssd1 vssd1 vccd1 vccd1 _07770_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09507_ _09507_/A _09507_/B vssd1 vssd1 vccd1 vccd1 _09509_/A sky130_fd_sc_hd__nand2_1
X_06719_ _08432_/B _06723_/C vssd1 vssd1 vccd1 vccd1 _06721_/A sky130_fd_sc_hd__nand2_1
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ _07699_/A _07699_/B vssd1 vssd1 vccd1 vccd1 _07702_/A sky130_fd_sc_hd__nand2_1
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ _09438_/A vssd1 vssd1 vccd1 vccd1 _09725_/A sky130_fd_sc_hd__inv_2
XFILLER_0_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09369_ _09368_/B _09369_/B _09369_/C vssd1 vssd1 vccd1 vccd1 _09641_/B sky130_fd_sc_hd__nand3b_2
XFILLER_0_74_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09429__B _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10213_ _10213_/A _10213_/B vssd1 vssd1 vccd1 vccd1 _10214_/B sky130_fd_sc_hd__xnor2_1
X_10144_ _10146_/C vssd1 vssd1 vccd1 vccd1 _10145_/B sky130_fd_sc_hd__inv_2
XFILLER_0_27_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10075_ _10075_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10076_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09164__B _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10103__B _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06979__A _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _10211_/A _09517_/C vssd1 vssd1 vccd1 vccd1 _08741_/C sky130_fd_sc_hd__nand2_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05952_ _05952_/A _06760_/A _06804_/A vssd1 vssd1 vccd1 vccd1 _05957_/B sky130_fd_sc_hd__nand3_1
X_08671_ _09133_/B _08813_/C vssd1 vssd1 vccd1 vccd1 _08811_/A sky130_fd_sc_hd__nand2_1
X_05883_ _06113_/A _06115_/B vssd1 vssd1 vccd1 vccd1 _05883_/Y sky130_fd_sc_hd__nor2_1
X_07622_ _07622_/A _07622_/B _07622_/C vssd1 vssd1 vccd1 vccd1 _07697_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_17_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09090__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07553_ _07614_/A _07613_/A vssd1 vssd1 vccd1 vccd1 _07553_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_75_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07484_ input12/X _07646_/D vssd1 vssd1 vccd1 vccd1 _07489_/A sky130_fd_sc_hd__nand2_1
X_06504_ _06504_/A _06504_/B _06504_/C vssd1 vssd1 vccd1 vccd1 _06659_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_75_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09223_ _09223_/A _09449_/A vssd1 vssd1 vccd1 vccd1 _09225_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_455 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06435_ _06439_/B _06436_/A vssd1 vssd1 vccd1 vccd1 _06438_/A sky130_fd_sc_hd__nand2_1
X_09154_ _09153_/B _09154_/B _09381_/B vssd1 vssd1 vccd1 vccd1 _09381_/A sky130_fd_sc_hd__nand3b_1
X_08105_ _08105_/A _08130_/A vssd1 vssd1 vccd1 vccd1 _08184_/B sky130_fd_sc_hd__nand2_1
X_06366_ _06504_/A _06504_/B vssd1 vssd1 vccd1 vccd1 _06372_/A sky130_fd_sc_hd__nand2_1
X_09085_ _09085_/A _09085_/B vssd1 vssd1 vccd1 vccd1 _09085_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_16_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06297_ _06317_/B _06295_/Y _06296_/Y vssd1 vssd1 vccd1 vccd1 _06494_/A sky130_fd_sc_hd__a21oi_2
X_08036_ _08149_/B _08149_/C vssd1 vssd1 vccd1 vccd1 _08049_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09265__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ _09987_/A vssd1 vssd1 vccd1 vccd1 _09988_/B sky130_fd_sc_hd__inv_2
X_08938_ _08939_/B _08938_/B _08938_/C vssd1 vssd1 vccd1 vccd1 _08998_/B sky130_fd_sc_hd__nand3_1
X_08869_ _08869_/A _08869_/B vssd1 vssd1 vccd1 vccd1 _08964_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09712__B _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05968__A _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ _10693_/A _10693_/B vssd1 vssd1 vccd1 vccd1 hold55/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10127_ _10127_/A _10127_/B vssd1 vssd1 vccd1 vccd1 _10136_/B sky130_fd_sc_hd__nand2_1
X_10058_ _10064_/B _10300_/B vssd1 vssd1 vccd1 vccd1 _10062_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_54_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09622__B _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06220_ _06220_/A _06220_/B vssd1 vssd1 vccd1 vccd1 _06300_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06151_ _06357_/A _06358_/B vssd1 vssd1 vccd1 vccd1 _06361_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_80_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06082_ _06082_/A _06891_/A _06082_/C vssd1 vssd1 vccd1 vccd1 _06084_/B sky130_fd_sc_hd__nand3_1
X_09910_ _10156_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _09916_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10711__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09841_ input50/X vssd1 vssd1 vccd1 vccd1 _10248_/C sky130_fd_sc_hd__inv_2
XFILLER_0_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ _09770_/Y _09541_/B _09771_/Y vssd1 vssd1 vccd1 vccd1 _09902_/A sky130_fd_sc_hd__a21oi_2
X_06984_ _07143_/A _07144_/B vssd1 vssd1 vccd1 vccd1 _06984_/Y sky130_fd_sc_hd__nor2_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _08781_/C _08781_/B _08722_/Y vssd1 vssd1 vccd1 vccd1 _08734_/B sky130_fd_sc_hd__a21oi_1
X_05935_ _05935_/A _06708_/B vssd1 vssd1 vccd1 vccd1 _05961_/A sky130_fd_sc_hd__nand2_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08654_ _08653_/B _08654_/B _09216_/B vssd1 vssd1 vccd1 vccd1 _09216_/A sky130_fd_sc_hd__nand3b_1
X_05866_ _09517_/C _10148_/A vssd1 vssd1 vccd1 vccd1 _05867_/A sky130_fd_sc_hd__nand2_1
X_05797_ _05797_/A vssd1 vssd1 vccd1 vccd1 _05798_/C sky130_fd_sc_hd__inv_2
XFILLER_0_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07605_ _07608_/A _07608_/B vssd1 vssd1 vccd1 vccd1 _07606_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07333__A _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08585_ input19/X vssd1 vssd1 vccd1 vccd1 _08587_/B sky130_fd_sc_hd__inv_2
XFILLER_0_48_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07536_ _07536_/A _07536_/B vssd1 vssd1 vccd1 vccd1 _07668_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07052__B _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09206_ _09206_/A _09206_/B vssd1 vssd1 vccd1 vccd1 _09214_/A sky130_fd_sc_hd__nand2_1
X_07467_ _07621_/A _07620_/A vssd1 vssd1 vccd1 vccd1 _07472_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_63_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07398_ _07398_/A _07398_/B _07398_/C vssd1 vssd1 vccd1 vccd1 _07405_/C sky130_fd_sc_hd__nand3_1
X_06418_ _06418_/A _06418_/B _06418_/C vssd1 vssd1 vccd1 vccd1 _06676_/C sky130_fd_sc_hd__nand3_1
X_06349_ _10040_/B input64/X vssd1 vssd1 vccd1 vccd1 _06545_/A sky130_fd_sc_hd__nand2_2
X_09137_ _09137_/A vssd1 vssd1 vccd1 vccd1 _09142_/B sky130_fd_sc_hd__inv_2
XFILLER_0_71_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09068_ _09068_/A _09068_/B vssd1 vssd1 vccd1 vccd1 _09072_/B sky130_fd_sc_hd__nand2_1
X_08019_ _08024_/A _08024_/C vssd1 vssd1 vccd1 vccd1 _08032_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09426__C _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08330__C _08366_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05970__B _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08339__A _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07897__B _07897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10676_ _10676_/A hold26/X vssd1 vssd1 vccd1 vccd1 hold27/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09489__B2 _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09489__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05720_ _06158_/A _06159_/B vssd1 vssd1 vccd1 vccd1 _06162_/C sky130_fd_sc_hd__nand2_1
X_05651_ _05651_/A _05651_/B vssd1 vssd1 vccd1 vccd1 _05653_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08370_ _10520_/C _08370_/B vssd1 vssd1 vccd1 vccd1 _10525_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07321_ _07321_/A _07321_/B _07321_/C vssd1 vssd1 vccd1 vccd1 _07509_/B sky130_fd_sc_hd__nand3_1
X_05582_ _05583_/B _05583_/A vssd1 vssd1 vccd1 vccd1 _05582_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_73_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07252_ _07250_/Y _07429_/B _07251_/Y vssd1 vssd1 vccd1 vccd1 _07583_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07183_ _07183_/A _07183_/B vssd1 vssd1 vccd1 vccd1 _07185_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06203_ _06203_/A _06203_/B vssd1 vssd1 vccd1 vccd1 _06382_/B sky130_fd_sc_hd__nand2_1
X_06134_ _06145_/B _06250_/A vssd1 vssd1 vccd1 vccd1 _06255_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06065_ _06067_/A _06067_/B vssd1 vssd1 vccd1 vccd1 _06066_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07328__A _08672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09824_ _09824_/A _09824_/B _09835_/A vssd1 vssd1 vccd1 vccd1 _10092_/B sky130_fd_sc_hd__nand3_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09755_ _09755_/A vssd1 vssd1 vccd1 vccd1 _09758_/A sky130_fd_sc_hd__inv_2
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06967_ _06967_/A _06967_/B vssd1 vssd1 vccd1 vccd1 _06969_/A sky130_fd_sc_hd__nand2_1
X_08706_ _09247_/B _08706_/B vssd1 vssd1 vccd1 vccd1 _08709_/A sky130_fd_sc_hd__nand2_1
X_09686_ _09686_/A vssd1 vssd1 vccd1 vccd1 _10022_/B sky130_fd_sc_hd__inv_2
X_06898_ _06898_/A _06898_/B vssd1 vssd1 vccd1 vccd1 _09037_/A sky130_fd_sc_hd__nand2_1
X_05918_ _05933_/A _05933_/B vssd1 vssd1 vccd1 vccd1 _05932_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08637_ _08633_/Y _08635_/Y _08638_/A vssd1 vssd1 vccd1 vccd1 _08643_/B sky130_fd_sc_hd__o21ai_1
X_05849_ _06183_/A _05850_/A vssd1 vssd1 vccd1 vccd1 _06302_/B sky130_fd_sc_hd__or2_1
XANTENNA__10201__B _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08568_ _08568_/A _08868_/A _08868_/B vssd1 vssd1 vccd1 vccd1 _08964_/C sky130_fd_sc_hd__nand3_2
XANTENNA__08455__A2 _09201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07519_ _07519_/A _07519_/B vssd1 vssd1 vccd1 vccd1 _07520_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08499_ _08571_/B _08499_/B vssd1 vssd1 vccd1 vccd1 _08501_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout98 fanout99/X vssd1 vssd1 vccd1 vccd1 fanout98/X sky130_fd_sc_hd__clkbuf_8
X_10530_ _10644_/A _10643_/A _10529_/Y vssd1 vssd1 vccd1 vccd1 _10538_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10461_ _10667_/B vssd1 vssd1 vccd1 vccd1 _10461_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_44_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10392_ _10725_/Q vssd1 vssd1 vccd1 vccd1 _10393_/B sky130_fd_sc_hd__inv_2
XANTENNA__09453__A _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09603__D _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10728_ _10733_/CLK _10728_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold61/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10659_ _10659_/A vssd1 vssd1 vccd1 vccd1 _10716_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__08532__A _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _07870_/A _07870_/B _07870_/C vssd1 vssd1 vccd1 vccd1 _07873_/A sky130_fd_sc_hd__nand3_1
XANTENNA__06987__A _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06821_ _06821_/A _06821_/B vssd1 vssd1 vccd1 vccd1 _06821_/Y sky130_fd_sc_hd__nor2_1
X_09540_ _09539_/Y _09103_/C _09108_/A vssd1 vssd1 vccd1 vccd1 _09541_/B sky130_fd_sc_hd__o21ai_2
X_06752_ _06752_/A vssd1 vssd1 vccd1 vccd1 _06753_/C sky130_fd_sc_hd__inv_2
X_09471_ _09471_/A _09471_/B vssd1 vssd1 vccd1 vccd1 _09473_/A sky130_fd_sc_hd__nand2_1
X_05703_ _06247_/B _05701_/Y _05702_/Y vssd1 vssd1 vccd1 vccd1 _06228_/B sky130_fd_sc_hd__a21oi_4
X_08422_ _08660_/A _08440_/B vssd1 vssd1 vccd1 vccd1 _08757_/B sky130_fd_sc_hd__nand2_1
X_06683_ _06947_/B _06671_/A _06672_/Y vssd1 vssd1 vccd1 vccd1 _06938_/A sky130_fd_sc_hd__a21oi_1
X_05634_ _05634_/A _05634_/B _05634_/C vssd1 vssd1 vccd1 vccd1 _05639_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_58_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05565_ _05709_/A _05709_/B vssd1 vssd1 vccd1 vccd1 _05580_/A sky130_fd_sc_hd__nand2_1
X_08353_ _08347_/B _08353_/B _08353_/C vssd1 vssd1 vccd1 vccd1 _08354_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__09634__A1 _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07304_ _07156_/Y _07314_/B _07170_/Y vssd1 vssd1 vccd1 vccd1 _07305_/A sky130_fd_sc_hd__a21o_1
X_08284_ _08291_/A vssd1 vssd1 vccd1 vccd1 _08285_/B sky130_fd_sc_hd__inv_2
X_05496_ _05496_/A _05496_/B vssd1 vssd1 vccd1 vccd1 _05498_/A sky130_fd_sc_hd__nand2_1
X_07235_ _07235_/A _07235_/B vssd1 vssd1 vccd1 vccd1 _07237_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07166_ _07166_/A vssd1 vssd1 vccd1 vccd1 _07167_/B sky130_fd_sc_hd__inv_2
X_06117_ _06117_/A _06117_/B vssd1 vssd1 vccd1 vccd1 _06179_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07097_ _07097_/A _07097_/B vssd1 vssd1 vccd1 vccd1 _07242_/A sky130_fd_sc_hd__nand2_1
X_06048_ _06047_/Y _09517_/C _09477_/C vssd1 vssd1 vccd1 vccd1 _06869_/B sky130_fd_sc_hd__nand3b_2
X_09807_ _09807_/A vssd1 vssd1 vccd1 vccd1 _09808_/A sky130_fd_sc_hd__inv_2
X_07999_ _07999_/A _07999_/B _07999_/C vssd1 vssd1 vccd1 vccd1 _08010_/B sky130_fd_sc_hd__nand3_1
X_09738_ _09742_/B _10070_/A vssd1 vssd1 vccd1 vccd1 _09741_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10212__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09669_ _09998_/A _09673_/C vssd1 vssd1 vccd1 vccd1 _09672_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10513_ hold23/X vssd1 vssd1 vccd1 vccd1 _10514_/B sky130_fd_sc_hd__inv_2
XANTENNA__06137__A _08453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10444_ _10467_/C _10472_/B vssd1 vssd1 vccd1 vccd1 _10445_/B sky130_fd_sc_hd__nor2_1
X_10375_ _10375_/A _10375_/B vssd1 vssd1 vccd1 vccd1 _10704_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09911__A _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08527__A _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07150__B _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05350_ input11/X vssd1 vssd1 vccd1 vccd1 _10151_/B sky130_fd_sc_hd__buf_4
XANTENNA__06047__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_264 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_223 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07020_ _07185_/C vssd1 vssd1 vccd1 vccd1 _07022_/B sky130_fd_sc_hd__inv_2
XANTENNA__08262__A _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08971_ _09031_/B _09031_/C vssd1 vssd1 vccd1 vccd1 _09030_/A sky130_fd_sc_hd__nand2_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_07922_ _07946_/A _07945_/B vssd1 vssd1 vccd1 vccd1 _07930_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09093__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ _08381_/A _07849_/Y _07852_/Y vssd1 vssd1 vccd1 vccd1 _10446_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__06510__A _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ _06804_/A _06804_/B vssd1 vssd1 vccd1 vccd1 _06804_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__07325__B input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07784_ _07797_/A _07797_/B vssd1 vssd1 vccd1 vccd1 _07795_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09523_ _09525_/B vssd1 vssd1 vccd1 vccd1 _09524_/B sky130_fd_sc_hd__inv_2
X_06735_ _06737_/A vssd1 vssd1 vccd1 vccd1 _06736_/B sky130_fd_sc_hd__inv_2
XFILLER_0_36_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09454_ _09677_/A _10004_/A _09678_/C _10005_/A vssd1 vssd1 vccd1 vccd1 _09454_/X
+ sky130_fd_sc_hd__and4_1
X_06666_ _06666_/A _06666_/B vssd1 vssd1 vccd1 vccd1 _06955_/C sky130_fd_sc_hd__nand2_1
X_08405_ _09922_/B vssd1 vssd1 vccd1 vccd1 _10188_/C sky130_fd_sc_hd__inv_2
X_05617_ _05617_/A _05617_/B vssd1 vssd1 vccd1 vccd1 _05620_/C sky130_fd_sc_hd__nand2_1
X_09385_ _10128_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _09390_/B sky130_fd_sc_hd__nand2_1
X_08336_ _10275_/B vssd1 vssd1 vccd1 vccd1 _09875_/D sky130_fd_sc_hd__inv_2
XFILLER_0_46_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06597_ _06597_/A _06685_/A vssd1 vssd1 vccd1 vccd1 _06948_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05548_ _05716_/C _05716_/B _05547_/Y vssd1 vssd1 vccd1 vccd1 _05564_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_19_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05479_ _05898_/B _05479_/B vssd1 vssd1 vccd1 vccd1 _05497_/A sky130_fd_sc_hd__nand2_1
X_08267_ _08300_/B _08301_/A _08266_/Y vssd1 vssd1 vccd1 vccd1 _08269_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07218_ _09840_/B _10158_/A vssd1 vssd1 vccd1 vccd1 _07222_/B sky130_fd_sc_hd__nand2_1
X_08198_ _08198_/A _08198_/B vssd1 vssd1 vccd1 vccd1 _08200_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08172__A _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07149_ _10212_/B _10108_/B vssd1 vssd1 vccd1 vccd1 _07319_/A sky130_fd_sc_hd__nand2_2
XANTENNA__08900__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10160_ _10160_/A _10160_/B vssd1 vssd1 vccd1 vccd1 _10162_/A sky130_fd_sc_hd__xnor2_1
X_10091_ _10334_/B _10093_/C vssd1 vssd1 vccd1 vccd1 _10092_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_69_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10427_ _10438_/A hold25/X _10438_/B vssd1 vssd1 vccd1 vccd1 _10675_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_33_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10358_ _10705_/B _10356_/X _10704_/B vssd1 vssd1 vccd1 vccd1 _10384_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_20_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10289_ _09884_/B input56/X _10292_/B _09882_/A vssd1 vssd1 vccd1 vccd1 _10290_/A
+ sky130_fd_sc_hd__a31oi_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10736__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06520_ _06649_/A _06650_/A vssd1 vssd1 vccd1 vccd1 _06653_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06451_ _06615_/A _06616_/A vssd1 vssd1 vccd1 vccd1 _06608_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08257__A _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05402_ _08114_/B input9/X vssd1 vssd1 vccd1 vccd1 _05682_/C sky130_fd_sc_hd__nand2_1
X_09170_ _09173_/B _09399_/A vssd1 vssd1 vccd1 vccd1 _09172_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06382_ _06382_/A _06382_/B vssd1 vssd1 vccd1 vccd1 _06384_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08121_ _08118_/C _08121_/B _08121_/C vssd1 vssd1 vccd1 vccd1 _08197_/B sky130_fd_sc_hd__nand3b_2
XFILLER_0_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08052_ _08052_/A _08052_/B vssd1 vssd1 vccd1 vccd1 _08092_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_31_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07003_ _07132_/A _07127_/A vssd1 vssd1 vccd1 vccd1 _07003_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__08720__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08954_ _08954_/A _09002_/B vssd1 vssd1 vccd1 vccd1 _08956_/A sky130_fd_sc_hd__nand2_1
X_07905_ _07905_/A _07905_/B vssd1 vssd1 vccd1 vccd1 _07906_/B sky130_fd_sc_hd__nand2_1
X_08885_ _08961_/A _08969_/A _08969_/B vssd1 vssd1 vccd1 vccd1 _08964_/A sky130_fd_sc_hd__a21boi_2
XFILLER_0_47_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07836_ _07836_/A _07836_/B vssd1 vssd1 vccd1 vccd1 _07838_/A sky130_fd_sc_hd__nand2_1
X_07767_ _07767_/A vssd1 vssd1 vccd1 vccd1 _07770_/A sky130_fd_sc_hd__inv_2
X_09506_ _09505_/B _09506_/B _09506_/C vssd1 vssd1 vccd1 vccd1 _09507_/B sky130_fd_sc_hd__nand3b_1
X_06718_ _06718_/A _06718_/B vssd1 vssd1 vccd1 vccd1 _06723_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07698_ _07701_/A _07701_/B vssd1 vssd1 vccd1 vccd1 _07699_/A sky130_fd_sc_hd__nand2_1
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09437_ _09725_/B _09438_/A vssd1 vssd1 vccd1 vccd1 _09443_/B sky130_fd_sc_hd__nand2_1
X_06649_ _06649_/A _06652_/A vssd1 vssd1 vccd1 vccd1 _06651_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_81_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ _09368_/A _09368_/B vssd1 vssd1 vccd1 vccd1 _09379_/A sky130_fd_sc_hd__nand2_1
X_09299_ _09299_/A _09299_/B vssd1 vssd1 vccd1 vccd1 _09301_/B sky130_fd_sc_hd__nand2_1
X_08319_ _08319_/A _08319_/B _08319_/C vssd1 vssd1 vccd1 vccd1 _08355_/B sky130_fd_sc_hd__nand3_2
XANTENNA__08264__B1 _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10212_ input46/X _10212_/B vssd1 vssd1 vccd1 vccd1 _10213_/B sky130_fd_sc_hd__nand2_1
X_10143_ _09988_/C _09988_/B _09965_/A vssd1 vssd1 vccd1 vccd1 _10146_/C sky130_fd_sc_hd__a21oi_1
X_10074_ _10074_/A _10075_/A _10075_/B vssd1 vssd1 vccd1 vccd1 _10077_/A sky130_fd_sc_hd__nand3_1
XANTENNA__06150__A _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06979__B _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05951_ _06804_/B _05951_/B vssd1 vssd1 vccd1 vccd1 _05957_/A sky130_fd_sc_hd__nand2_1
X_08670_ _08670_/A _08670_/B vssd1 vssd1 vccd1 vccd1 _08813_/C sky130_fd_sc_hd__nand2_2
X_05882_ _06115_/B _06113_/A vssd1 vssd1 vccd1 vccd1 _05882_/Y sky130_fd_sc_hd__nand2_1
X_07621_ _07621_/A _07621_/B vssd1 vssd1 vccd1 vccd1 _07622_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09090__B _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07552_ _07613_/A _07614_/A vssd1 vssd1 vccd1 vccd1 _07612_/C sky130_fd_sc_hd__nand2_1
X_06503_ _06701_/A _07284_/A vssd1 vssd1 vccd1 vccd1 _06699_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07483_ _07493_/A _07493_/B vssd1 vssd1 vccd1 vccd1 _07491_/A sky130_fd_sc_hd__nand2_1
X_09222_ _09222_/A _09223_/A _09449_/A vssd1 vssd1 vccd1 vccd1 _09512_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_63_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06434_ _06437_/B vssd1 vssd1 vccd1 vccd1 _06439_/B sky130_fd_sc_hd__inv_2
XFILLER_0_56_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09153_ _09153_/A _09153_/B vssd1 vssd1 vccd1 vccd1 _09159_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06365_ _06365_/A _06365_/B _06365_/C vssd1 vssd1 vccd1 vccd1 _06504_/B sky130_fd_sc_hd__nand3_1
X_08104_ _08130_/B _08104_/B _08104_/C vssd1 vssd1 vccd1 vccd1 _08130_/A sky130_fd_sc_hd__nand3_1
X_09084_ _09085_/B _09085_/A vssd1 vssd1 vccd1 vccd1 _09084_/Y sky130_fd_sc_hd__nand2_1
X_06296_ _06315_/A _06314_/A vssd1 vssd1 vccd1 vccd1 _06296_/Y sky130_fd_sc_hd__nor2_1
X_08035_ _08033_/A _08033_/B _08052_/A vssd1 vssd1 vccd1 vccd1 _08149_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09265__B _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09986_ _09986_/A _09987_/A vssd1 vssd1 vccd1 vccd1 _09993_/A sky130_fd_sc_hd__nand2_1
X_08937_ _08937_/A _08937_/B vssd1 vssd1 vccd1 vccd1 _08938_/C sky130_fd_sc_hd__nand2_1
X_08868_ _08868_/A _08868_/B vssd1 vssd1 vccd1 vccd1 _08869_/A sky130_fd_sc_hd__nand2_1
X_07819_ _07822_/B vssd1 vssd1 vccd1 vccd1 _07823_/A sky130_fd_sc_hd__inv_2
X_08799_ _08905_/A _08799_/B vssd1 vssd1 vccd1 vccd1 _08800_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09712__C _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10692_ _10694_/A vssd1 vssd1 vccd1 vccd1 _10693_/A sky130_fd_sc_hd__inv_2
XANTENNA__05968__B _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05984__A _07756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ _10140_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10126_/X sky130_fd_sc_hd__and2_1
X_10057_ _10230_/A _10057_/B _10057_/C vssd1 vssd1 vccd1 vccd1 _10300_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09191__A _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10130__A _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06150_ _10210_/B input64/X vssd1 vssd1 vccd1 vccd1 _06358_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_79_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06081_ _06081_/A _06081_/B vssd1 vssd1 vccd1 vccd1 _06084_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09840_ input51/X _09840_/B vssd1 vssd1 vccd1 vccd1 _09846_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _09771_/A _09771_/B vssd1 vssd1 vccd1 vccd1 _09771_/Y sky130_fd_sc_hd__nor2_1
X_06983_ _07145_/C vssd1 vssd1 vccd1 vccd1 _07147_/B sky130_fd_sc_hd__inv_2
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _10248_/B _10202_/C _08722_/C vssd1 vssd1 vccd1 vccd1 _08722_/Y sky130_fd_sc_hd__nor3_1
X_05934_ _05936_/B _05936_/C vssd1 vssd1 vccd1 vccd1 _06708_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_28_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08653_ _08653_/A _08653_/B vssd1 vssd1 vccd1 vccd1 _08657_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05865_ _05868_/A _05868_/B vssd1 vssd1 vccd1 vccd1 _06170_/C sky130_fd_sc_hd__nand2_1
XANTENNA__10040__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05796_ _05796_/A _06040_/A _06020_/A vssd1 vssd1 vccd1 vccd1 _05798_/B sky130_fd_sc_hd__nand3_1
X_08584_ _09156_/B _08597_/C vssd1 vssd1 vccd1 vccd1 _08595_/A sky130_fd_sc_hd__nand2_1
X_07604_ _07604_/A _07604_/B _07604_/C vssd1 vssd1 vccd1 vccd1 _07608_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07333__B _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07535_ _07535_/A _07535_/B _07535_/C vssd1 vssd1 vccd1 vccd1 _07536_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07466_ _07621_/B vssd1 vssd1 vccd1 vccd1 _07620_/A sky130_fd_sc_hd__inv_2
XFILLER_0_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09205_ _09205_/A _09205_/B vssd1 vssd1 vccd1 vccd1 _09206_/B sky130_fd_sc_hd__xor2_1
XFILLER_0_8_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06417_ _06417_/A _06417_/B vssd1 vssd1 vccd1 vccd1 _06676_/B sky130_fd_sc_hd__nand2_1
X_07397_ _07477_/B _07397_/B vssd1 vssd1 vccd1 vccd1 _07408_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06348_ _08725_/A vssd1 vssd1 vccd1 vccd1 _10040_/B sky130_fd_sc_hd__buf_8
X_09136_ _10115_/A input19/X vssd1 vssd1 vccd1 vccd1 _09137_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09067_ _09069_/B vssd1 vssd1 vccd1 vccd1 _09068_/B sky130_fd_sc_hd__inv_2
X_06279_ _06283_/B _06280_/A vssd1 vssd1 vccd1 vccd1 _06282_/A sky130_fd_sc_hd__nand2_1
X_08018_ _08018_/A _08018_/B _08030_/A vssd1 vssd1 vccd1 vccd1 _08024_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_8_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09426__D _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ input17/X vssd1 vssd1 vccd1 vccd1 _09971_/B sky130_fd_sc_hd__inv_2
XFILLER_0_67_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10675_ _10675_/A _10675_/B vssd1 vssd1 vccd1 vccd1 hold26/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10109_ _10109_/A vssd1 vssd1 vccd1 vccd1 _10110_/B sky130_fd_sc_hd__inv_2
XANTENNA__09489__A2 _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05650_ _05650_/A _05650_/B vssd1 vssd1 vccd1 vccd1 _05651_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05581_ _05564_/B _05563_/A _05712_/B vssd1 vssd1 vccd1 vccd1 _05626_/B sky130_fd_sc_hd__o21ai_2
X_07320_ _07322_/A _07320_/B vssd1 vssd1 vccd1 vccd1 _07321_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07251_ _07427_/A _07426_/A vssd1 vssd1 vccd1 vccd1 _07251_/Y sky130_fd_sc_hd__nor2_1
X_07182_ _07357_/C _07182_/B vssd1 vssd1 vccd1 vccd1 _07195_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_26_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06202_ _06202_/A _06202_/B vssd1 vssd1 vccd1 vccd1 _06203_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06133_ _06284_/C _06284_/B _06132_/Y vssd1 vssd1 vccd1 vccd1 _06250_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06064_ input46/X _09778_/D vssd1 vssd1 vccd1 vccd1 _06067_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06513__A _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07328__B _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _09823_/A _09823_/B vssd1 vssd1 vccd1 vccd1 _09827_/B sky130_fd_sc_hd__nand2_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09754_ _09490_/B _10210_/A _10247_/B _09488_/X vssd1 vssd1 vccd1 vccd1 _09755_/A
+ sky130_fd_sc_hd__a31o_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06966_ _07124_/B _07124_/C vssd1 vssd1 vccd1 vccd1 _07123_/A sky130_fd_sc_hd__nand2_1
X_08705_ _09247_/A vssd1 vssd1 vccd1 vccd1 _08706_/B sky130_fd_sc_hd__inv_2
X_09685_ _09687_/B _09687_/A vssd1 vssd1 vccd1 vccd1 _09686_/A sky130_fd_sc_hd__nor2_1
X_06897_ _06899_/C vssd1 vssd1 vccd1 vccd1 _06898_/B sky130_fd_sc_hd__inv_2
X_05917_ _05917_/A _06711_/A _06734_/A vssd1 vssd1 vccd1 vccd1 _05933_/B sky130_fd_sc_hd__nand3_1
X_05848_ _05848_/A _05848_/B vssd1 vssd1 vccd1 vccd1 _05850_/A sky130_fd_sc_hd__xor2_1
X_08636_ _10156_/A _09602_/B vssd1 vssd1 vccd1 vccd1 _08638_/A sky130_fd_sc_hd__nand2_1
X_08567_ _08567_/A _08567_/B _08570_/A vssd1 vssd1 vccd1 vccd1 _08868_/B sky130_fd_sc_hd__nand3_2
X_05779_ _06020_/A vssd1 vssd1 vccd1 vccd1 _05795_/B sky130_fd_sc_hd__inv_2
XFILLER_0_64_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07518_ _07518_/A _07518_/B _07518_/C vssd1 vssd1 vccd1 vccd1 _07667_/B sky130_fd_sc_hd__nand3_2
X_08498_ _08498_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08499_/B sky130_fd_sc_hd__nand2_1
X_07449_ _07449_/A _07449_/B _07449_/C vssd1 vssd1 vccd1 vccd1 _07450_/B sky130_fd_sc_hd__nand3_1
Xfanout99 input65/X vssd1 vssd1 vccd1 vccd1 fanout99/X sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10460_ _10460_/A hold59/X _10460_/C vssd1 vssd1 vccd1 vccd1 _10667_/B sky130_fd_sc_hd__nand3_1
X_09119_ _09119_/A _09119_/B _09544_/A vssd1 vssd1 vccd1 vccd1 _09564_/B sky130_fd_sc_hd__nand3_2
X_10391_ _10394_/A _10394_/B vssd1 vssd1 vccd1 vccd1 _10393_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09453__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10727_ _10733_/CLK hold32/X fanout98/X vssd1 vssd1 vccd1 vccd1 hold31/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10658_ _10658_/A _10660_/A vssd1 vssd1 vccd1 vccd1 _10659_/A sky130_fd_sc_hd__and2_1
XFILLER_0_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10589_ hold8/X _10589_/B vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__nand2_1
XANTENNA__08532__B _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06987__B _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ _06821_/B _06821_/A vssd1 vssd1 vccd1 vccd1 _06820_/Y sky130_fd_sc_hd__nand2_1
X_06751_ _06751_/A _06752_/A vssd1 vssd1 vccd1 vccd1 _06758_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07164__A _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09470_ _09470_/A _09470_/B vssd1 vssd1 vccd1 vccd1 _09471_/B sky130_fd_sc_hd__or2_1
X_06682_ _06948_/C vssd1 vssd1 vccd1 vccd1 _06947_/B sky130_fd_sc_hd__inv_2
X_05702_ _06240_/A _06245_/A vssd1 vssd1 vccd1 vccd1 _05702_/Y sky130_fd_sc_hd__nor2_1
X_08421_ _08421_/A _08421_/B _08421_/C vssd1 vssd1 vccd1 vccd1 _08440_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_25_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05633_ _06106_/B _06106_/C vssd1 vssd1 vccd1 vccd1 _06108_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_25_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05564_ _05564_/A _05564_/B _05564_/C vssd1 vssd1 vccd1 vccd1 _05709_/B sky130_fd_sc_hd__nand3_1
X_08352_ _08352_/A _08352_/B _08352_/C vssd1 vssd1 vccd1 vccd1 _08353_/C sky130_fd_sc_hd__and3_1
X_05495_ _05497_/C vssd1 vssd1 vccd1 vccd1 _05496_/B sky130_fd_sc_hd__inv_2
X_08283_ _08283_/A _08291_/A vssd1 vssd1 vccd1 vccd1 _08330_/B sky130_fd_sc_hd__nand2_1
X_07303_ _07303_/A _07303_/B _07303_/C vssd1 vssd1 vccd1 vccd1 _07308_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07234_ _07405_/B _07234_/B vssd1 vssd1 vccd1 vccd1 _07235_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07165_ _07165_/A _07166_/A vssd1 vssd1 vccd1 vccd1 _07168_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06116_ _06118_/A _06118_/B vssd1 vssd1 vccd1 vccd1 _06117_/A sky130_fd_sc_hd__nand2_1
X_07096_ _07096_/A _07096_/B vssd1 vssd1 vccd1 vccd1 _07097_/B sky130_fd_sc_hd__nand2_1
X_06047_ _09517_/D _09698_/A vssd1 vssd1 vccd1 vccd1 _06047_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_1_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09806_ _09806_/A _09807_/A vssd1 vssd1 vccd1 vccd1 _09813_/B sky130_fd_sc_hd__nand2_1
X_07998_ _07998_/A _07998_/B vssd1 vssd1 vccd1 vccd1 _08010_/C sky130_fd_sc_hd__nand2_1
X_09737_ _09737_/A _09737_/B _10070_/B vssd1 vssd1 vccd1 vccd1 _10070_/A sky130_fd_sc_hd__nand3_2
X_06949_ _07255_/B _07255_/C vssd1 vssd1 vccd1 vccd1 _07254_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10212__B _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09668_ _09668_/A _09668_/B vssd1 vssd1 vccd1 vccd1 _09673_/C sky130_fd_sc_hd__nand2_1
X_09599_ _09600_/B _09600_/A vssd1 vssd1 vccd1 vccd1 _09936_/B sky130_fd_sc_hd__or2_1
X_08619_ _08619_/A _08619_/B vssd1 vssd1 vccd1 vccd1 _08620_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10512_ _10520_/A _10520_/C vssd1 vssd1 vccd1 vccd1 _10514_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06137__B _07785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10443_ _10443_/A _10443_/B _10672_/B vssd1 vssd1 vccd1 vccd1 _10548_/A sky130_fd_sc_hd__nand3_1
X_10374_ _10374_/A _10558_/B vssd1 vssd1 vccd1 vccd1 _10383_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05992__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09911__B _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06047__B _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06063__A _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07159__A _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08262__B _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08970_ _08970_/A _08970_/B vssd1 vssd1 vccd1 vccd1 _09031_/C sky130_fd_sc_hd__nand2_1
X_07921_ _07945_/A _07946_/B vssd1 vssd1 vccd1 vccd1 _07930_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09552__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__B2 _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__B _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ _07852_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _07852_/Y sky130_fd_sc_hd__nor2_1
X_06803_ _06804_/B _06804_/A vssd1 vssd1 vccd1 vccd1 _06803_/Y sky130_fd_sc_hd__nand2_1
Xinput1 a_i[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__buf_4
XANTENNA__05407__A _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ input51/X _10275_/B vssd1 vssd1 vccd1 vccd1 _09525_/B sky130_fd_sc_hd__nand2_1
X_07783_ _07783_/A _07783_/B _07783_/C vssd1 vssd1 vccd1 vccd1 _07797_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08718__A _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06734_ _06734_/A _06734_/B vssd1 vssd1 vccd1 vccd1 _06737_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09453_ _10201_/A _10187_/B vssd1 vssd1 vccd1 vccd1 _09458_/B sky130_fd_sc_hd__nand2_1
X_06665_ _06665_/A _06665_/B _06665_/C vssd1 vssd1 vccd1 vccd1 _06666_/B sky130_fd_sc_hd__nand3_1
X_08404_ _08445_/B _08402_/Y _08444_/A vssd1 vssd1 vccd1 vccd1 _08418_/A sky130_fd_sc_hd__a21oi_1
X_05616_ _05616_/A _05616_/B _05616_/C vssd1 vssd1 vccd1 vccd1 _05617_/B sky130_fd_sc_hd__nand3_1
X_09384_ _09407_/A _09620_/B vssd1 vssd1 vccd1 vccd1 _09405_/A sky130_fd_sc_hd__nand2_1
X_08335_ _08335_/A vssd1 vssd1 vccd1 vccd1 _08353_/B sky130_fd_sc_hd__inv_2
X_06596_ _07081_/B _06685_/B _06596_/C vssd1 vssd1 vccd1 vccd1 _06685_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_61_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05547_ _05547_/A _05547_/B vssd1 vssd1 vccd1 vccd1 _05547_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09549__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08453__A _08453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05478_ _05898_/A vssd1 vssd1 vccd1 vccd1 _05479_/B sky130_fd_sc_hd__inv_2
XFILLER_0_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08266_ _08266_/A _08266_/B vssd1 vssd1 vccd1 vccd1 _08266_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_61_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07217_ _09749_/B _10157_/A vssd1 vssd1 vccd1 vccd1 _07222_/A sky130_fd_sc_hd__nand2_1
X_08197_ _08197_/A _08197_/B vssd1 vssd1 vccd1 vccd1 _08201_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07148_ _07312_/B _07312_/C vssd1 vssd1 vccd1 vccd1 _07311_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08172__B _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08900__B _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07079_ _07079_/A vssd1 vssd1 vccd1 vccd1 _07097_/A sky130_fd_sc_hd__inv_2
X_10090_ _10090_/A _10090_/B vssd1 vssd1 vccd1 vccd1 _10093_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_16_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06148__A _08725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05987__A _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10426_ _10426_/A _10426_/B _10426_/C vssd1 vssd1 vccd1 vccd1 _10438_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_33_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10357_ _10357_/A hold41/X _10357_/C vssd1 vssd1 vccd1 vccd1 _10704_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_20_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10288_ _09882_/A _10274_/Y _10287_/Y vssd1 vssd1 vccd1 vccd1 _10294_/B sky130_fd_sc_hd__o21ai_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09922__A _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08257__B _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06450_ _06625_/C _06625_/B _06449_/Y vssd1 vssd1 vccd1 vccd1 _06616_/A sky130_fd_sc_hd__a21oi_1
X_05401_ _05680_/A _05681_/B vssd1 vssd1 vccd1 vccd1 _05684_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_16_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06381_ _06489_/B _06410_/C vssd1 vssd1 vccd1 vccd1 _06409_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08120_ _08120_/A _08120_/B vssd1 vssd1 vccd1 vccd1 _08121_/C sky130_fd_sc_hd__nand2_1
X_08051_ _08051_/A _08051_/B vssd1 vssd1 vccd1 vccd1 _08091_/B sky130_fd_sc_hd__nand2_1
X_07002_ _07130_/B _07130_/C _07001_/Y vssd1 vssd1 vccd1 vccd1 _07127_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08720__B _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08953_ _08998_/A _08998_/B _08999_/A vssd1 vssd1 vccd1 vccd1 _09002_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06521__A _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07904_ _07905_/B _07905_/A vssd1 vssd1 vccd1 vccd1 _08061_/B sky130_fd_sc_hd__or2_2
X_08884_ _08884_/A _08884_/B _08884_/C vssd1 vssd1 vccd1 vccd1 _08969_/B sky130_fd_sc_hd__nand3_2
X_07835_ _07835_/A _07835_/B _07835_/C vssd1 vssd1 vccd1 vccd1 _07836_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_78_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07766_ _07951_/C vssd1 vssd1 vccd1 vccd1 _07950_/B sky130_fd_sc_hd__inv_2
XFILLER_0_2_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09505_ _09505_/A _09505_/B vssd1 vssd1 vccd1 vccd1 _09507_/A sky130_fd_sc_hd__nand2_1
X_06717_ _06718_/A _06718_/B vssd1 vssd1 vccd1 vccd1 _08432_/B sky130_fd_sc_hd__or2_1
XFILLER_0_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ _09436_/A _09436_/B vssd1 vssd1 vccd1 vccd1 _09438_/A sky130_fd_sc_hd__nand2_1
X_07697_ _07697_/A _07697_/B _07697_/C vssd1 vssd1 vccd1 vccd1 _07701_/B sky130_fd_sc_hd__nand3_1
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06648_ _06642_/C _06642_/B _06518_/Y vssd1 vssd1 vccd1 vccd1 _06652_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_81_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06579_ _06579_/A _06579_/B _06579_/C vssd1 vssd1 vccd1 vccd1 _07078_/B sky130_fd_sc_hd__nand3_1
X_09367_ _09140_/A _09140_/B _09145_/C vssd1 vssd1 vccd1 vccd1 _09368_/B sky130_fd_sc_hd__o21a_1
X_09298_ _08813_/B _08813_/C _09133_/B vssd1 vssd1 vccd1 vccd1 _09299_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_19_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08318_ _08346_/B vssd1 vssd1 vccd1 vccd1 _08319_/C sky130_fd_sc_hd__inv_2
XANTENNA__08264__A1 _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08264__B2 _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08249_ _08249_/A _08275_/B _08249_/C vssd1 vssd1 vccd1 vccd1 _08292_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_15_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10211_ _10211_/A _10211_/B vssd1 vssd1 vccd1 vccd1 _10213_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10142_ _10146_/A _10146_/B vssd1 vssd1 vccd1 vccd1 _10145_/A sky130_fd_sc_hd__nand2_1
X_10073_ _10073_/A _10073_/B _10073_/C vssd1 vssd1 vccd1 vccd1 _10075_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06150__B input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10128__A _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10409_ _10409_/A vssd1 vssd1 vccd1 vccd1 _10410_/B sky130_fd_sc_hd__inv_2
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05950_ _06804_/A vssd1 vssd1 vccd1 vccd1 _05951_/B sky130_fd_sc_hd__inv_2
X_05881_ _05870_/Y _06188_/B _05880_/Y vssd1 vssd1 vccd1 vccd1 _06113_/A sky130_fd_sc_hd__a21oi_1
X_07620_ _07620_/A _07620_/B vssd1 vssd1 vccd1 vccd1 _07622_/A sky130_fd_sc_hd__nand2_1
X_07551_ _07540_/Y _07663_/B _07550_/Y vssd1 vssd1 vccd1 vccd1 _07614_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06502_ _06502_/A _06502_/B _06502_/C vssd1 vssd1 vccd1 vccd1 _07284_/A sky130_fd_sc_hd__nand3_4
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07482_ _07384_/Y _07482_/B _07482_/C vssd1 vssd1 vccd1 vccd1 _07493_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_33_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09221_ _09220_/B _09221_/B _09449_/B vssd1 vssd1 vccd1 vccd1 _09449_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_8_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06433_ _06605_/B _06605_/C vssd1 vssd1 vccd1 vccd1 _06610_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09099__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09152_ _09152_/A _09397_/C vssd1 vssd1 vccd1 vccd1 _09153_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06364_ _06364_/A _06364_/B vssd1 vssd1 vccd1 vccd1 _06504_/A sky130_fd_sc_hd__nand2_1
X_08103_ _08130_/B _08104_/C _08104_/B vssd1 vssd1 vccd1 vccd1 _08105_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06516__A _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09083_ _09081_/Y _08958_/B _09082_/Y vssd1 vssd1 vccd1 vccd1 _09308_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_16_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06295_ _06314_/A _06315_/A vssd1 vssd1 vccd1 vccd1 _06295_/Y sky130_fd_sc_hd__nand2_1
X_08034_ _08052_/A _08052_/B vssd1 vssd1 vccd1 vccd1 _08149_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_12_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09985_ _09985_/A _10166_/A vssd1 vssd1 vccd1 vccd1 _09987_/A sky130_fd_sc_hd__nand2_1
X_08936_ _08949_/B _08949_/A vssd1 vssd1 vccd1 vccd1 _08938_/B sky130_fd_sc_hd__nor2_1
X_08867_ _08967_/C vssd1 vssd1 vccd1 vccd1 _08966_/B sky130_fd_sc_hd__inv_2
X_07818_ _07823_/B vssd1 vssd1 vccd1 vccd1 _07822_/A sky130_fd_sc_hd__inv_2
X_08798_ _08798_/A _08798_/B vssd1 vssd1 vccd1 vccd1 _08799_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09712__D _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07749_ _08725_/A _08114_/B vssd1 vssd1 vccd1 vccd1 _07946_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09419_ _09598_/B _09419_/B vssd1 vssd1 vccd1 vccd1 _09421_/A sky130_fd_sc_hd__and2_1
X_10691_ _10691_/A hold29/X vssd1 vssd1 vccd1 vccd1 hold30/A sky130_fd_sc_hd__xnor2_1
XANTENNA__07810__A _07811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10125_ _10140_/B _10140_/A vssd1 vssd1 vccd1 vccd1 _10125_/Y sky130_fd_sc_hd__nor2_1
X_10056_ _10056_/A vssd1 vssd1 vccd1 vccd1 _10057_/C sky130_fd_sc_hd__inv_2
XANTENNA__09191__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05505__A _07891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06336__A _07756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06080_ _06082_/A vssd1 vssd1 vccd1 vccd1 _06081_/B sky130_fd_sc_hd__inv_2
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ _09771_/B _09771_/A vssd1 vssd1 vccd1 vccd1 _09770_/Y sky130_fd_sc_hd__nand2_1
X_06982_ _10115_/A _09677_/A vssd1 vssd1 vccd1 vccd1 _07145_/C sky130_fd_sc_hd__nand2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _08721_/A vssd1 vssd1 vccd1 vccd1 _08781_/B sky130_fd_sc_hd__inv_2
X_05933_ _05933_/A _05933_/B _05933_/C vssd1 vssd1 vccd1 vccd1 _05936_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_28_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08652_ _09237_/A _08652_/B vssd1 vssd1 vccd1 vccd1 _08653_/B sky130_fd_sc_hd__xor2_1
X_07603_ _07603_/A _07603_/B vssd1 vssd1 vccd1 vccd1 _07608_/A sky130_fd_sc_hd__nand2_1
X_05864_ _07675_/A _10151_/A vssd1 vssd1 vccd1 vccd1 _05868_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10040__B _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05795_ _06020_/B _05795_/B vssd1 vssd1 vccd1 vccd1 _05798_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10720__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08583_ _08583_/A _08583_/B vssd1 vssd1 vccd1 vccd1 _08597_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_48_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07534_ _07534_/A _07534_/B vssd1 vssd1 vccd1 vccd1 _07536_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07465_ _08739_/A _07785_/B vssd1 vssd1 vccd1 vccd1 _07621_/B sky130_fd_sc_hd__nand2_1
X_09204_ _09459_/A _09204_/B vssd1 vssd1 vccd1 vccd1 _09205_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_29_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06416_ _06418_/A _06418_/B vssd1 vssd1 vccd1 vccd1 _06417_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07396_ _07396_/A _07397_/B _07396_/C vssd1 vssd1 vccd1 vccd1 _07477_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06347_ _07675_/A _07646_/D vssd1 vssd1 vccd1 vccd1 _06546_/B sky130_fd_sc_hd__nand2_1
X_09135_ _09135_/A _09135_/B vssd1 vssd1 vccd1 vccd1 _09145_/A sky130_fd_sc_hd__nand2_1
X_09066_ _09064_/Y _09331_/C _09065_/Y vssd1 vssd1 vccd1 vccd1 _09336_/A sky130_fd_sc_hd__a21oi_2
X_06278_ _06281_/B vssd1 vssd1 vccd1 vccd1 _06283_/B sky130_fd_sc_hd__inv_2
X_08017_ _08030_/B _08017_/B vssd1 vssd1 vccd1 vccd1 _08024_/A sky130_fd_sc_hd__nand2_1
X_09968_ _10128_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _09976_/B sky130_fd_sc_hd__nand2_1
X_08919_ input49/X _10284_/B input50/X _08897_/B vssd1 vssd1 vccd1 vccd1 _08920_/B
+ sky130_fd_sc_hd__a22o_1
X_09899_ _10319_/B _09899_/B vssd1 vssd1 vccd1 vccd1 _09907_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08636__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10674_ _10674_/A vssd1 vssd1 vccd1 vccd1 _10720_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10108_ _10112_/A _10108_/B input20/X input21/X vssd1 vssd1 vccd1 vccd1 _10110_/A
+ sky130_fd_sc_hd__and4_1
X_10039_ _10048_/A _10048_/C vssd1 vssd1 vccd1 vccd1 _10046_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05580_ _05580_/A _05580_/B vssd1 vssd1 vccd1 vccd1 _05712_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07250_ _07426_/A _07427_/A vssd1 vssd1 vccd1 vccd1 _07250_/Y sky130_fd_sc_hd__nand2_1
X_07181_ _07182_/B _07181_/B _07181_/C vssd1 vssd1 vccd1 vccd1 _07357_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_26_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06201_ _06201_/A _06202_/B _06202_/A vssd1 vssd1 vccd1 vccd1 _06382_/A sky130_fd_sc_hd__nand3_1
X_06132_ _06280_/A _06281_/B vssd1 vssd1 vccd1 vccd1 _06132_/Y sky130_fd_sc_hd__nor2_1
X_06063_ _10211_/A input1/X vssd1 vssd1 vccd1 vccd1 _06067_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06513__B _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09824__B _09824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09822_ _09824_/A vssd1 vssd1 vccd1 vccd1 _09823_/B sky130_fd_sc_hd__inv_2
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09753_ _09839_/A _09753_/B vssd1 vssd1 vccd1 vccd1 _09758_/B sky130_fd_sc_hd__nand2_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07625__A _08672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08704_ _08394_/A _08703_/Y _08395_/A vssd1 vssd1 vccd1 vccd1 _09247_/A sky130_fd_sc_hd__a21oi_2
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06965_ _06965_/A _06965_/B _06965_/C vssd1 vssd1 vccd1 vccd1 _07124_/C sky130_fd_sc_hd__nand3_2
X_09684_ _10003_/A _09684_/B vssd1 vssd1 vccd1 vccd1 _09687_/A sky130_fd_sc_hd__nand2_1
X_06896_ _06896_/A _06896_/B vssd1 vssd1 vccd1 vccd1 _06899_/C sky130_fd_sc_hd__nand2_1
X_05916_ _06711_/B _05916_/B vssd1 vssd1 vccd1 vccd1 _05933_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09840__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05847_ _05847_/A _05821_/Y vssd1 vssd1 vccd1 vccd1 _05848_/B sky130_fd_sc_hd__nor2b_1
X_08635_ _08639_/C vssd1 vssd1 vccd1 vccd1 _08635_/Y sky130_fd_sc_hd__inv_2
X_08566_ _08566_/A _08566_/B vssd1 vssd1 vccd1 vccd1 _08868_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08456__A _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05778_ _05577_/C _05577_/B _05570_/A vssd1 vssd1 vccd1 vccd1 _06020_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07360__A _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07517_ _07519_/A _07517_/B vssd1 vssd1 vccd1 vccd1 _07518_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08497_ _08498_/A _08498_/B vssd1 vssd1 vccd1 vccd1 _08571_/B sky130_fd_sc_hd__or2_1
X_07448_ _07448_/A _07448_/B vssd1 vssd1 vccd1 vccd1 _07450_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07379_ _10275_/B _10157_/A vssd1 vssd1 vccd1 vccd1 _07384_/A sky130_fd_sc_hd__nand2_1
X_09118_ _09118_/A vssd1 vssd1 vccd1 vccd1 _09119_/A sky130_fd_sc_hd__inv_2
X_10390_ _10389_/B _10390_/B _10390_/C vssd1 vssd1 vccd1 vccd1 _10394_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_32_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09049_ _09069_/B _09068_/A vssd1 vssd1 vccd1 vccd1 _09049_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_67_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10726_ _10733_/CLK _10726_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold54/A sky130_fd_sc_hd__dfrtp_1
X_10657_ _10657_/A _10657_/B vssd1 vssd1 vccd1 vccd1 _10660_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10588_ hold7/X _10588_/B hold15/A vssd1 vssd1 vccd1 vccd1 _10589_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06750_ _10128_/A _09602_/B vssd1 vssd1 vccd1 vccd1 _06752_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07164__B _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06681_ _06938_/B _06938_/C vssd1 vssd1 vccd1 vccd1 _06939_/A sky130_fd_sc_hd__nand2_1
X_05701_ _06245_/A _06240_/A vssd1 vssd1 vccd1 vccd1 _05701_/Y sky130_fd_sc_hd__nand2_1
X_08420_ _08420_/A _08420_/B vssd1 vssd1 vccd1 vccd1 _08421_/C sky130_fd_sc_hd__nand2_1
X_05632_ _05632_/A _05632_/B _05632_/C vssd1 vssd1 vccd1 vccd1 _06106_/C sky130_fd_sc_hd__nand3_1
X_05563_ _05563_/A _05563_/B vssd1 vssd1 vccd1 vccd1 _05709_/A sky130_fd_sc_hd__nand2_1
X_08351_ _08351_/A _10292_/B _10103_/A vssd1 vssd1 vccd1 vccd1 _08352_/C sky130_fd_sc_hd__and3_1
XFILLER_0_58_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05494_ _05494_/A _05494_/B vssd1 vssd1 vccd1 vccd1 _05497_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_6_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07302_ _07432_/B _07432_/C vssd1 vssd1 vccd1 vccd1 _07437_/B sky130_fd_sc_hd__nand2_1
X_08282_ _08282_/A _08287_/A _08287_/B vssd1 vssd1 vccd1 vccd1 _08291_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07233_ _07233_/A _07233_/B vssd1 vssd1 vccd1 vccd1 _07234_/B sky130_fd_sc_hd__or2_1
XFILLER_0_33_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07164_ _10210_/B _10101_/A vssd1 vssd1 vccd1 vccd1 _07166_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06524__A _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06115_ _06115_/A _06115_/B vssd1 vssd1 vccd1 vccd1 _06118_/B sky130_fd_sc_hd__nand2_1
X_07095_ _07095_/A vssd1 vssd1 vccd1 vccd1 _07415_/A sky130_fd_sc_hd__inv_2
XANTENNA__09835__A _09835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06046_ _06075_/A _06075_/B vssd1 vssd1 vccd1 vccd1 _06074_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09805_ _10083_/A _09805_/B vssd1 vssd1 vccd1 vccd1 _09807_/A sky130_fd_sc_hd__nand2_1
X_07997_ _07999_/A _07999_/B vssd1 vssd1 vccd1 vccd1 _07998_/A sky130_fd_sc_hd__nand2_1
X_09736_ _09736_/A vssd1 vssd1 vccd1 vccd1 _09737_/A sky130_fd_sc_hd__inv_2
X_06948_ _06948_/A _06948_/B _06948_/C vssd1 vssd1 vccd1 vccd1 _07255_/C sky130_fd_sc_hd__nand3_1
X_09667_ _09667_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _09668_/A sky130_fd_sc_hd__nand2_1
X_06879_ _06881_/A vssd1 vssd1 vccd1 vccd1 _06880_/B sky130_fd_sc_hd__inv_2
X_08618_ _08618_/A _08618_/B vssd1 vssd1 vccd1 vccd1 _08619_/A sky130_fd_sc_hd__nand2_1
X_09598_ _09598_/A _09598_/B vssd1 vssd1 vccd1 vccd1 _09600_/A sky130_fd_sc_hd__and2_1
X_08549_ _08549_/A _08549_/B vssd1 vssd1 vccd1 vccd1 _08550_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_436 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10511_ _10511_/A _10511_/B vssd1 vssd1 vccd1 vccd1 _10520_/A sky130_fd_sc_hd__or2_1
XFILLER_0_52_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10442_ _10442_/A vssd1 vssd1 vccd1 vccd1 _10672_/B sky130_fd_sc_hd__inv_2
X_10373_ _10558_/A _10558_/B _10373_/C vssd1 vssd1 vccd1 vccd1 _10374_/A sky130_fd_sc_hd__nand3_1
XANTENNA__09745__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05992__B _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05513__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10709_ _10709_/A vssd1 vssd1 vccd1 vccd1 _10730_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_86 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07159__B _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08262__C _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06063__B input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07920_ _07946_/A vssd1 vssd1 vccd1 vccd1 _07945_/A sky130_fd_sc_hd__inv_2
XANTENNA__09552__A2 _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07851_ _07851_/A _07851_/B vssd1 vssd1 vccd1 vccd1 _08385_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07175__A _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06802_ _08822_/A _06808_/C vssd1 vssd1 vccd1 vccd1 _08975_/B sky130_fd_sc_hd__nand2_1
X_07782_ _07782_/A _07782_/B vssd1 vssd1 vccd1 vccd1 _07783_/B sky130_fd_sc_hd__nand2_1
Xinput2 a_i[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__05407__B _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ _09525_/A vssd1 vssd1 vccd1 vccd1 _09524_/A sky130_fd_sc_hd__inv_2
X_06733_ _06737_/B _08478_/A vssd1 vssd1 vccd1 vccd1 _06736_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08718__B _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09452_ _09510_/B _09739_/B vssd1 vssd1 vccd1 vccd1 _09508_/A sky130_fd_sc_hd__nand2_1
X_06664_ _06664_/A vssd1 vssd1 vccd1 vccd1 _06665_/A sky130_fd_sc_hd__inv_2
X_08403_ _09912_/A _10188_/A _08403_/C vssd1 vssd1 vccd1 vccd1 _08444_/A sky130_fd_sc_hd__nor3_1
X_05615_ _05615_/A vssd1 vssd1 vccd1 vccd1 _05616_/B sky130_fd_sc_hd__inv_2
XFILLER_0_46_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09383_ _09382_/B _09383_/B _09641_/A vssd1 vssd1 vccd1 vccd1 _09620_/B sky130_fd_sc_hd__nand3b_1
X_06595_ _06595_/A _07081_/B vssd1 vssd1 vccd1 vccd1 _06597_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05546_ _05546_/A vssd1 vssd1 vccd1 vccd1 _05716_/B sky130_fd_sc_hd__inv_2
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ _08334_/A _08334_/B vssd1 vssd1 vccd1 vccd1 _08335_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08453__B _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08265_ _08299_/B _08265_/B vssd1 vssd1 vccd1 vccd1 _08301_/A sky130_fd_sc_hd__and2_1
X_05477_ _05356_/C _05356_/B _05476_/Y vssd1 vssd1 vccd1 vccd1 _05898_/A sky130_fd_sc_hd__a21oi_2
X_07216_ _07226_/B _07226_/C vssd1 vssd1 vccd1 vccd1 _07233_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08196_ _08271_/B _08272_/A _08195_/Y vssd1 vssd1 vccd1 vccd1 _08206_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07147_ _07147_/A _07147_/B _07147_/C vssd1 vssd1 vccd1 vccd1 _07312_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_14_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07078_ _07078_/A _07078_/B vssd1 vssd1 vccd1 vccd1 _07080_/A sky130_fd_sc_hd__nand2_1
X_06029_ _06841_/B _06033_/C vssd1 vssd1 vccd1 vccd1 _06032_/A sky130_fd_sc_hd__nand2_1
X_09719_ _09719_/A _09719_/B vssd1 vssd1 vccd1 vccd1 _09722_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_69_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06148__B _07646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05987__B _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08363__B _08363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10425_ _10425_/A _10425_/B vssd1 vssd1 vccd1 vccd1 _10438_/A sky130_fd_sc_hd__nand2_1
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10356_ _10375_/A _10375_/B vssd1 vssd1 vccd1 vccd1 _10356_/X sky130_fd_sc_hd__and2_1
X_10287_ _10290_/C _10290_/B vssd1 vssd1 vccd1 vccd1 _10287_/Y sky130_fd_sc_hd__nand2_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09922__B _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06339__A _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05400_ _08574_/A _09602_/B vssd1 vssd1 vccd1 vccd1 _05681_/B sky130_fd_sc_hd__nand2_1
X_06380_ _06380_/A _06380_/B vssd1 vssd1 vccd1 vccd1 _06410_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_43_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08050_ _08212_/B _08148_/A vssd1 vssd1 vccd1 vccd1 _08051_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_22_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_322 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07001_ _07138_/A _07137_/A vssd1 vssd1 vccd1 vccd1 _07001_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09385__A _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08952_ _09005_/B _09005_/A vssd1 vssd1 vccd1 vccd1 _08999_/A sky130_fd_sc_hd__nor2_1
X_08883_ _08883_/A _08883_/B vssd1 vssd1 vccd1 vccd1 _08969_/A sky130_fd_sc_hd__nand2_2
X_07903_ _07976_/A _07903_/B vssd1 vssd1 vccd1 vccd1 _07905_/A sky130_fd_sc_hd__and2_1
XANTENNA__06521__B _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07834_ _07834_/A _07834_/B vssd1 vssd1 vccd1 vccd1 _07836_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08729__A _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09551__C _09551_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07633__A _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07765_ _07765_/A _07782_/A vssd1 vssd1 vccd1 vccd1 _07951_/C sky130_fd_sc_hd__nand2_1
X_09504_ _09251_/B _09250_/A _09285_/A vssd1 vssd1 vccd1 vccd1 _09505_/B sky130_fd_sc_hd__o21ai_2
X_07696_ _07696_/A _07696_/B vssd1 vssd1 vccd1 vccd1 _07701_/A sky130_fd_sc_hd__nand2_1
X_06716_ _10103_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _06718_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09435_ _09439_/A _09615_/A vssd1 vssd1 vccd1 vccd1 _09725_/B sky130_fd_sc_hd__nand2_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06647_ _06962_/A _06957_/A vssd1 vssd1 vccd1 vccd1 _06647_/Y sky130_fd_sc_hd__nand2_1
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09366_ _09369_/B _09369_/C vssd1 vssd1 vccd1 vccd1 _09368_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06578_ _06578_/A _06581_/A vssd1 vssd1 vccd1 vccd1 _07078_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09297_ _09297_/A _09512_/A vssd1 vssd1 vccd1 vccd1 _09299_/A sky130_fd_sc_hd__nand2_1
X_05529_ _05894_/B _05894_/A vssd1 vssd1 vccd1 vccd1 _05530_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08264__A2 _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08317_ _08345_/B _08345_/A vssd1 vssd1 vccd1 vccd1 _08346_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08248_ _08249_/A _08275_/B _08249_/C vssd1 vssd1 vccd1 vccd1 _08292_/A sky130_fd_sc_hd__a21o_1
X_10210_ _10210_/A _10210_/B vssd1 vssd1 vccd1 vccd1 _10214_/A sky130_fd_sc_hd__nand2_1
X_08179_ _08251_/C _08251_/B vssd1 vssd1 vccd1 vccd1 _08252_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10141_ _10141_/A _10141_/B _10141_/C vssd1 vssd1 vccd1 vccd1 _10146_/B sky130_fd_sc_hd__nand3_1
X_10072_ _10072_/A _10072_/B vssd1 vssd1 vccd1 vccd1 _10075_/A sky130_fd_sc_hd__nand2_1
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10408_ _10408_/A _10409_/A vssd1 vssd1 vccd1 vccd1 _10419_/A sky130_fd_sc_hd__nand2_1
X_10339_ _10573_/A _10339_/B _10339_/C vssd1 vssd1 vccd1 vccd1 _10343_/C sky130_fd_sc_hd__nand3_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05880_ _06186_/C _06185_/A vssd1 vssd1 vccd1 vccd1 _05880_/Y sky130_fd_sc_hd__nor2_1
X_07550_ _07656_/A _07661_/A vssd1 vssd1 vccd1 vccd1 _07550_/Y sky130_fd_sc_hd__nor2_1
X_06501_ _07274_/A vssd1 vssd1 vccd1 vccd1 _06502_/C sky130_fd_sc_hd__inv_2
XFILLER_0_75_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09220_ _09220_/A _09220_/B vssd1 vssd1 vccd1 vccd1 _09223_/A sky130_fd_sc_hd__nand2_1
X_07481_ _07384_/Y _07480_/Y _07383_/A vssd1 vssd1 vccd1 vccd1 _07493_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_33_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06432_ _06432_/A _06432_/B _06432_/C vssd1 vssd1 vccd1 vccd1 _06605_/C sky130_fd_sc_hd__nand3_1
X_09151_ _09151_/A _10101_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _09397_/C sky130_fd_sc_hd__nand3_1
X_06363_ _06365_/A vssd1 vssd1 vccd1 vccd1 _06364_/B sky130_fd_sc_hd__inv_2
X_09082_ _09082_/A _09082_/B vssd1 vssd1 vccd1 vccd1 _09082_/Y sky130_fd_sc_hd__nor2_1
X_08102_ _08102_/A vssd1 vssd1 vccd1 vccd1 _08104_/B sky130_fd_sc_hd__inv_2
XANTENNA__06516__B _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08033_ _08033_/A _08033_/B vssd1 vssd1 vccd1 vccd1 _08052_/B sky130_fd_sc_hd__nor2_1
X_06294_ _06417_/B _06292_/Y _06293_/Y vssd1 vssd1 vccd1 vccd1 _06315_/A sky130_fd_sc_hd__a21oi_2
Xinput60 b_i[5] vssd1 vssd1 vccd1 vccd1 input60/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09984_ _10166_/B _09984_/B _09984_/C vssd1 vssd1 vccd1 vccd1 _10166_/A sky130_fd_sc_hd__nand3_1
X_08935_ _08935_/A _08935_/B vssd1 vssd1 vccd1 vccd1 _08949_/A sky130_fd_sc_hd__and2_1
X_08866_ _08866_/A _08866_/B vssd1 vssd1 vccd1 vccd1 _08967_/C sky130_fd_sc_hd__nand2_1
X_08797_ _08797_/A vssd1 vssd1 vccd1 vccd1 _08798_/B sky130_fd_sc_hd__inv_2
X_07817_ _07815_/Y _07967_/B _07816_/Y vssd1 vssd1 vccd1 vccd1 _08067_/B sky130_fd_sc_hd__a21oi_1
X_07748_ _07916_/A _07917_/A vssd1 vssd1 vccd1 vccd1 _07919_/B sky130_fd_sc_hd__nand2_1
X_07679_ _07769_/B vssd1 vssd1 vccd1 vccd1 _07768_/B sky130_fd_sc_hd__inv_2
XFILLER_0_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09418_ _10158_/A _10151_/B _10157_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _09419_/B
+ sky130_fd_sc_hd__a22o_1
X_10690_ _10690_/A _10690_/B vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__nand2_1
X_09349_ _10365_/C vssd1 vssd1 vccd1 vccd1 _09350_/B sky130_fd_sc_hd__inv_2
XFILLER_0_47_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06442__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10124_ _10124_/A _10124_/B vssd1 vssd1 vccd1 vccd1 _10140_/A sky130_fd_sc_hd__nand2_1
X_10055_ _10055_/A _10056_/A vssd1 vssd1 vccd1 vccd1 _10064_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05505__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06336__B _07891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _07143_/A _07144_/B vssd1 vssd1 vccd1 vccd1 _07147_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _08739_/A _10201_/B vssd1 vssd1 vccd1 vccd1 _08721_/A sky130_fd_sc_hd__nand2_1
X_05932_ _05932_/A _05932_/B vssd1 vssd1 vccd1 vccd1 _05936_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_28_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _08651_/A _08651_/B vssd1 vssd1 vccd1 vccd1 _08652_/B sky130_fd_sc_hd__nor2_1
X_05863_ _08739_/A input37/X vssd1 vssd1 vccd1 vccd1 _05868_/A sky130_fd_sc_hd__nand2_1
X_07602_ _07604_/A vssd1 vssd1 vccd1 vccd1 _07603_/B sky130_fd_sc_hd__inv_2
X_05794_ _05794_/A _05794_/B _05797_/A vssd1 vssd1 vccd1 vccd1 _05801_/A sky130_fd_sc_hd__nand3_1
X_08582_ _08501_/B _08501_/A _08571_/B vssd1 vssd1 vccd1 vccd1 _08583_/B sky130_fd_sc_hd__o21a_1
X_07533_ _07535_/A _07535_/C vssd1 vssd1 vccd1 vccd1 _07534_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07464_ _07620_/B vssd1 vssd1 vccd1 vccd1 _07621_/A sky130_fd_sc_hd__inv_2
XFILLER_0_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09203_ _09203_/A vssd1 vssd1 vccd1 vccd1 _09204_/B sky130_fd_sc_hd__inv_2
XANTENNA__06527__A _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06415_ _06415_/A _06415_/B vssd1 vssd1 vccd1 vccd1 _06418_/B sky130_fd_sc_hd__nand2_1
X_09134_ _09134_/A _09134_/B vssd1 vssd1 vccd1 vccd1 _09222_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07395_ _07450_/C vssd1 vssd1 vccd1 vccd1 _07396_/C sky130_fd_sc_hd__inv_2
XFILLER_0_71_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06346_ _06476_/A _06477_/A vssd1 vssd1 vccd1 vccd1 _06346_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09065_ _09328_/C _09327_/A vssd1 vssd1 vccd1 vccd1 _09065_/Y sky130_fd_sc_hd__nor2_1
X_06277_ _06430_/A _06431_/A vssd1 vssd1 vccd1 vccd1 _06422_/B sky130_fd_sc_hd__nand2_1
X_08016_ _08030_/A vssd1 vssd1 vccd1 vccd1 _08017_/B sky130_fd_sc_hd__inv_2
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09967_ _09988_/A _09988_/C vssd1 vssd1 vccd1 vccd1 _09986_/A sky130_fd_sc_hd__nand2_1
X_08918_ _08916_/Y _08925_/C vssd1 vssd1 vccd1 vccd1 _08924_/A sky130_fd_sc_hd__nand2b_1
X_09898_ _10319_/A vssd1 vssd1 vccd1 vccd1 _09899_/B sky130_fd_sc_hd__inv_2
XANTENNA__05606__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08849_ _10210_/A _10284_/B vssd1 vssd1 vccd1 vccd1 _08856_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08636__B _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05341__A _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10673_ _10673_/A _10675_/A vssd1 vssd1 vccd1 vccd1 _10674_/A sky130_fd_sc_hd__and2_1
X_10107_ _10107_/A vssd1 vssd1 vccd1 vccd1 _10123_/B sky130_fd_sc_hd__inv_2
X_10038_ _10259_/B _10259_/A vssd1 vssd1 vccd1 vccd1 _10048_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_77_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06347__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06200_ _06200_/A _06200_/B vssd1 vssd1 vccd1 vccd1 _06202_/A sky130_fd_sc_hd__nand2_1
X_07180_ _07349_/B _07350_/B vssd1 vssd1 vccd1 vccd1 _07181_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09949__A2 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06131_ _06282_/C vssd1 vssd1 vccd1 vccd1 _06284_/B sky130_fd_sc_hd__inv_2
X_06062_ input47/X vssd1 vssd1 vccd1 vccd1 _10211_/A sky130_fd_sc_hd__buf_4
XFILLER_0_53_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07178__A _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09821_ _09821_/A _09821_/B vssd1 vssd1 vccd1 vccd1 _09824_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09824__C _09835_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07906__A _08061_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09752_ _09752_/A _09752_/B vssd1 vssd1 vccd1 vccd1 _09753_/B sky130_fd_sc_hd__nand2_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07625__B _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08703_ _08703_/A vssd1 vssd1 vccd1 vccd1 _08703_/Y sky130_fd_sc_hd__inv_2
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06964_ _06964_/A _06964_/B vssd1 vssd1 vccd1 vccd1 _07124_/B sky130_fd_sc_hd__nand2_1
X_09683_ _09683_/A _09683_/B vssd1 vssd1 vccd1 vccd1 _09684_/B sky130_fd_sc_hd__nand2_1
X_06895_ _06895_/A _06895_/B _06895_/C vssd1 vssd1 vccd1 vccd1 _06896_/B sky130_fd_sc_hd__nand3_1
X_05915_ _06711_/A vssd1 vssd1 vccd1 vccd1 _05916_/B sky130_fd_sc_hd__inv_2
XANTENNA__09840__B _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08634_ _09912_/A _08633_/B _08633_/C vssd1 vssd1 vccd1 vccd1 _08639_/C sky130_fd_sc_hd__o21ai_2
XFILLER_0_55_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05846_ _05846_/A vssd1 vssd1 vccd1 vccd1 _06183_/A sky130_fd_sc_hd__inv_2
X_08565_ _08567_/A vssd1 vssd1 vccd1 vccd1 _08566_/B sky130_fd_sc_hd__inv_2
X_05777_ _05765_/Y _05858_/B _05776_/Y vssd1 vssd1 vccd1 vccd1 _05800_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_49_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08456__B _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07360__B _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07516_ _07516_/A vssd1 vssd1 vccd1 vccd1 _07519_/A sky130_fd_sc_hd__inv_2
XFILLER_0_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08496_ _08574_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _08498_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07447_ _07713_/B _07713_/C vssd1 vssd1 vccd1 vccd1 _07715_/B sky130_fd_sc_hd__nand2_1
X_07378_ _07449_/A _07449_/B vssd1 vssd1 vccd1 vccd1 _07448_/A sky130_fd_sc_hd__nand2_1
X_09117_ _09117_/A _09118_/A vssd1 vssd1 vccd1 vccd1 _09123_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06329_ _08453_/A _08101_/B vssd1 vssd1 vccd1 vccd1 _06456_/C sky130_fd_sc_hd__nand2_1
X_09048_ _09068_/A _09069_/B vssd1 vssd1 vccd1 vccd1 _09048_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__07088__A _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06720__A _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08128__A1 _09551_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09876__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09876__B2 _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08647__A _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08366__B _08366_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10725_ _10733_/CLK hold30/X fanout98/X vssd1 vssd1 vccd1 vccd1 _10725_/Q sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10656_ _10657_/B _10657_/A vssd1 vssd1 vccd1 vccd1 _10658_/A sky130_fd_sc_hd__or2_1
XFILLER_0_35_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10587_ _10587_/A hold7/X vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06630__A _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09941__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06680_ _06939_/B _06938_/B _06938_/C vssd1 vssd1 vccd1 vccd1 _06687_/B sky130_fd_sc_hd__nand3_1
X_05700_ _06243_/B _06243_/C _05699_/Y vssd1 vssd1 vccd1 vccd1 _06240_/A sky130_fd_sc_hd__a21oi_1
X_05631_ _05892_/A _05631_/B _05631_/C vssd1 vssd1 vccd1 vccd1 _05632_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_25_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08350_ _09875_/D _09393_/A _08342_/C vssd1 vssd1 vccd1 vccd1 _08352_/B sky130_fd_sc_hd__o21ai_1
X_05562_ _05564_/B vssd1 vssd1 vccd1 vccd1 _05563_/B sky130_fd_sc_hd__inv_2
XFILLER_0_46_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07301_ _07301_/A _07301_/B _07301_/C vssd1 vssd1 vccd1 vccd1 _07432_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_73_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05493_ _05493_/A _05493_/B _05493_/C vssd1 vssd1 vccd1 vccd1 _05494_/B sky130_fd_sc_hd__nand3_1
X_08281_ _08281_/A _08289_/B vssd1 vssd1 vccd1 vccd1 _08287_/A sky130_fd_sc_hd__nand2_1
X_07232_ _07232_/A _07232_/B vssd1 vssd1 vccd1 vccd1 _07405_/B sky130_fd_sc_hd__nand2_1
X_07163_ _07167_/A _07167_/C vssd1 vssd1 vccd1 vccd1 _07165_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06114_ _05870_/Y _06188_/B _05880_/Y vssd1 vssd1 vccd1 vccd1 _06115_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06524__B _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07094_ _07414_/B _07414_/A vssd1 vssd1 vccd1 vccd1 _07095_/A sky130_fd_sc_hd__nor2_1
X_06045_ _06890_/A _06045_/B _06045_/C vssd1 vssd1 vccd1 vccd1 _06075_/B sky130_fd_sc_hd__nand3_1
X_09804_ _09804_/A _09804_/B _09804_/C vssd1 vssd1 vccd1 vccd1 _09805_/B sky130_fd_sc_hd__nand3_1
X_07996_ _07996_/A _07996_/B vssd1 vssd1 vccd1 vccd1 _07999_/A sky130_fd_sc_hd__nand2_1
X_09735_ _09735_/A _09736_/A vssd1 vssd1 vccd1 vccd1 _09742_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_66_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06947_ _06947_/A _06947_/B vssd1 vssd1 vccd1 vccd1 _07255_/B sky130_fd_sc_hd__nand2_1
X_09666_ _09666_/A _09998_/B _09667_/A vssd1 vssd1 vccd1 vccd1 _09998_/A sky130_fd_sc_hd__nand3_2
X_06878_ _08951_/A _06878_/B vssd1 vssd1 vccd1 vccd1 _06881_/A sky130_fd_sc_hd__nand2_1
X_08617_ _08619_/B _08618_/A _08618_/B vssd1 vssd1 vccd1 vccd1 _08620_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__08530__A1 _09971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05829_ input1/X vssd1 vssd1 vccd1 vccd1 _08897_/B sky130_fd_sc_hd__buf_6
X_09597_ _09918_/A _09597_/B vssd1 vssd1 vccd1 vccd1 _09600_/B sky130_fd_sc_hd__nand2_1
X_08548_ _08567_/B _08570_/A vssd1 vssd1 vccd1 vccd1 _08566_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08479_ _08491_/B vssd1 vssd1 vccd1 vccd1 _08480_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10510_ _10510_/A _10510_/B vssd1 vssd1 vccd1 vccd1 _10540_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10441_ _10441_/A _10675_/B vssd1 vssd1 vccd1 vccd1 _10442_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10372_ _10697_/B vssd1 vssd1 vccd1 vccd1 _10373_/C sky130_fd_sc_hd__inv_2
XANTENNA__09745__B input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10708_ _10708_/A _10708_/B vssd1 vssd1 vccd1 vccd1 _10709_/A sky130_fd_sc_hd__and2_1
XFILLER_0_43_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10639_ _10642_/A _10639_/B vssd1 vssd1 vccd1 vccd1 _10640_/A sky130_fd_sc_hd__and2_1
XFILLER_0_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08262__D _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07456__A _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07850_ _07850_/A _07850_/B vssd1 vssd1 vccd1 vccd1 _07851_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07175__B _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06801_ _06801_/A _06801_/B _06801_/C vssd1 vssd1 vccd1 vccd1 _06808_/C sky130_fd_sc_hd__nand3_1
X_07781_ _07781_/A _07781_/B vssd1 vssd1 vccd1 vccd1 _07797_/A sky130_fd_sc_hd__nand2_1
X_09520_ _09759_/B _09520_/B vssd1 vssd1 vccd1 vccd1 _09525_/A sky130_fd_sc_hd__nand2_1
X_06732_ _06731_/B _08478_/B _06732_/C vssd1 vssd1 vccd1 vccd1 _08478_/A sky130_fd_sc_hd__nand3b_2
Xinput3 a_i[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__05704__A _06229_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09451_ _09450_/B _09451_/B _09670_/A vssd1 vssd1 vccd1 vccd1 _09739_/B sky130_fd_sc_hd__nand3b_2
X_06663_ _06663_/A _06664_/A vssd1 vssd1 vccd1 vccd1 _06666_/A sky130_fd_sc_hd__nand2_1
X_08402_ _08447_/B vssd1 vssd1 vccd1 vccd1 _08402_/Y sky130_fd_sc_hd__inv_2
X_05614_ _05614_/A _05615_/A vssd1 vssd1 vccd1 vccd1 _05617_/A sky130_fd_sc_hd__nand2_1
X_09382_ _09382_/A _09382_/B vssd1 vssd1 vccd1 vccd1 _09407_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06594_ _07078_/A _07078_/B _07079_/A vssd1 vssd1 vccd1 vccd1 _07081_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05545_ _08724_/A input35/X vssd1 vssd1 vccd1 vccd1 _05546_/A sky130_fd_sc_hd__nand2_1
X_08333_ _08315_/A _08316_/B _08315_/C vssd1 vssd1 vccd1 vccd1 _08334_/A sky130_fd_sc_hd__a21o_1
X_08264_ _09840_/B _10103_/A _10292_/B _10103_/B vssd1 vssd1 vccd1 vccd1 _08265_/B
+ sky130_fd_sc_hd__a22o_1
XANTENNA__06535__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05476_ _05476_/A _05476_/B vssd1 vssd1 vccd1 vccd1 _05476_/Y sky130_fd_sc_hd__nor2_1
X_08195_ _08195_/A _08195_/B vssd1 vssd1 vccd1 vccd1 _08195_/Y sky130_fd_sc_hd__nor2_1
X_07215_ _07215_/A _07215_/B _07215_/C vssd1 vssd1 vccd1 vccd1 _07226_/C sky130_fd_sc_hd__nand3_1
X_07146_ _07146_/A _07146_/B vssd1 vssd1 vccd1 vccd1 _07147_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07077_ _07084_/A vssd1 vssd1 vccd1 vccd1 _07083_/A sky130_fd_sc_hd__inv_2
X_06028_ _06028_/A _06028_/B vssd1 vssd1 vccd1 vccd1 _06033_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06270__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09718_ _09718_/A _09718_/B _09718_/C vssd1 vssd1 vccd1 vccd1 _09719_/B sky130_fd_sc_hd__nand3_1
X_07979_ _07979_/A _07979_/B vssd1 vssd1 vccd1 vccd1 _07980_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09700__B1 _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09649_ _09982_/B _09649_/B vssd1 vssd1 vccd1 vccd1 _09651_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06445__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10424_ _10426_/B vssd1 vssd1 vccd1 vccd1 _10425_/B sky130_fd_sc_hd__inv_2
XFILLER_0_33_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09519__B1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10355_ hold41/X vssd1 vssd1 vccd1 vccd1 _10375_/B sky130_fd_sc_hd__inv_2
X_10286_ _10285_/B _10286_/B _10286_/C vssd1 vssd1 vccd1 vccd1 _10290_/B sky130_fd_sc_hd__nand3b_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06339__B _07897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07000_ _07139_/C vssd1 vssd1 vccd1 vccd1 _07130_/C sky130_fd_sc_hd__inv_2
XFILLER_0_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09385__B _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08951_ _08951_/A _08951_/B vssd1 vssd1 vccd1 vccd1 _09005_/A sky130_fd_sc_hd__and2_1
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08882_ _08884_/B vssd1 vssd1 vccd1 vccd1 _08883_/B sky130_fd_sc_hd__inv_2
X_07902_ _07902_/A _07902_/B vssd1 vssd1 vccd1 vccd1 _07903_/B sky130_fd_sc_hd__or2_1
XANTENNA__10714__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07833_ _08084_/A _08384_/A _08083_/B vssd1 vssd1 vccd1 vccd1 _08382_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08729__B _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__D _09782_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07633__B _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _07782_/B _07764_/B _07764_/C vssd1 vssd1 vccd1 vccd1 _07782_/A sky130_fd_sc_hd__nand3_1
X_09503_ _09506_/B _09506_/C vssd1 vssd1 vccd1 vccd1 _09505_/A sky130_fd_sc_hd__nand2_1
X_07695_ _07697_/A vssd1 vssd1 vccd1 vccd1 _07696_/B sky130_fd_sc_hd__inv_2
X_06715_ input16/X vssd1 vssd1 vccd1 vccd1 _10128_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__05434__A _07897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09434_ _09433_/B _09615_/B _09434_/C vssd1 vssd1 vccd1 vccd1 _09615_/A sky130_fd_sc_hd__nand3b_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06646_ _06960_/B _06960_/C _06645_/Y vssd1 vssd1 vccd1 vccd1 _06957_/A sky130_fd_sc_hd__a21oi_1
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ _09365_/A _09365_/B vssd1 vssd1 vccd1 vccd1 _09369_/C sky130_fd_sc_hd__nand2_1
X_06577_ _06579_/B vssd1 vssd1 vccd1 vccd1 _06581_/A sky130_fd_sc_hd__inv_2
X_09296_ _09296_/A _09297_/A _09512_/A vssd1 vssd1 vccd1 vccd1 _09572_/B sky130_fd_sc_hd__nand3_2
X_05528_ _05533_/B vssd1 vssd1 vccd1 vccd1 _05530_/B sky130_fd_sc_hd__inv_2
X_08316_ _08334_/B _08316_/B vssd1 vssd1 vccd1 vccd1 _08345_/A sky130_fd_sc_hd__nand2_1
X_08247_ _08285_/A _08363_/B vssd1 vssd1 vccd1 vccd1 _08283_/A sky130_fd_sc_hd__nand2_1
X_05459_ _05459_/A _05459_/B vssd1 vssd1 vccd1 vccd1 _05639_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08178_ _08175_/A _08175_/B _08176_/Y vssd1 vssd1 vccd1 vccd1 _08251_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07129_ _07137_/B _07138_/C _07138_/B vssd1 vssd1 vccd1 vccd1 _07131_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10140_ _10140_/A _10140_/B vssd1 vssd1 vccd1 vccd1 _10141_/C sky130_fd_sc_hd__nand2_1
X_10071_ _10073_/A vssd1 vssd1 vccd1 vccd1 _10072_/B sky130_fd_sc_hd__inv_2
XFILLER_0_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_69_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08390__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10407_ _10415_/A _10410_/C vssd1 vssd1 vccd1 vccd1 _10408_/A sky130_fd_sc_hd__nand2_1
X_10338_ _10338_/A vssd1 vssd1 vccd1 vccd1 _10339_/B sky130_fd_sc_hd__inv_2
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10269_ _09861_/C _09861_/B _09858_/A vssd1 vssd1 vccd1 vccd1 _10272_/C sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07480_ _07482_/C vssd1 vssd1 vccd1 vccd1 _07480_/Y sky130_fd_sc_hd__inv_2
X_06500_ _06500_/A _07274_/A vssd1 vssd1 vccd1 vccd1 _06701_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06431_ _06431_/A _06431_/B _06431_/C vssd1 vssd1 vccd1 vccd1 _06432_/B sky130_fd_sc_hd__nand3_1
X_09150_ _10101_/A _10158_/B _09151_/A vssd1 vssd1 vccd1 vccd1 _09152_/A sky130_fd_sc_hd__a21o_1
X_06362_ _06365_/B _06365_/C vssd1 vssd1 vccd1 vccd1 _06364_/A sky130_fd_sc_hd__nand2_1
X_09081_ _09082_/B _09082_/A vssd1 vssd1 vccd1 vccd1 _09081_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08101_ _09778_/D _08101_/B vssd1 vssd1 vccd1 vccd1 _08102_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06293_ _06413_/A _06415_/A vssd1 vssd1 vccd1 vccd1 _06293_/Y sky130_fd_sc_hd__nor2_1
X_08032_ _08032_/A _08032_/B vssd1 vssd1 vccd1 vccd1 _08033_/B sky130_fd_sc_hd__and2_1
Xinput50 b_i[25] vssd1 vssd1 vccd1 vccd1 input50/X sky130_fd_sc_hd__buf_4
Xinput61 b_i[6] vssd1 vssd1 vccd1 vccd1 input61/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09983_ _10166_/B _09984_/C _09984_/B vssd1 vssd1 vccd1 vccd1 _09985_/A sky130_fd_sc_hd__a21o_1
X_08934_ input49/X _10292_/B vssd1 vssd1 vccd1 vccd1 _08949_/B sky130_fd_sc_hd__nand2_1
X_08865_ _08864_/B _08865_/B _08865_/C vssd1 vssd1 vccd1 vccd1 _08866_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__08459__B _09201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08796_ _09268_/A _10276_/B _08795_/C vssd1 vssd1 vccd1 vccd1 _08797_/A sky130_fd_sc_hd__o21ai_1
X_07816_ _07964_/A _07965_/B vssd1 vssd1 vccd1 vccd1 _07816_/Y sky130_fd_sc_hd__nor2_1
X_07747_ _09710_/B _08573_/A vssd1 vssd1 vccd1 vccd1 _07917_/A sky130_fd_sc_hd__nand2_1
X_07678_ _08724_/A _08114_/B vssd1 vssd1 vccd1 vccd1 _07769_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09417_ _09417_/A vssd1 vssd1 vccd1 vccd1 _09598_/B sky130_fd_sc_hd__inv_2
X_06629_ _06973_/A _06974_/B vssd1 vssd1 vccd1 vccd1 _06977_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_81_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09348_ _10385_/A _09348_/B vssd1 vssd1 vccd1 vccd1 _10348_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _09285_/A _09285_/B vssd1 vssd1 vccd1 vccd1 _09557_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_229 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10123_ _10123_/A _10123_/B vssd1 vssd1 vccd1 vccd1 _10124_/B sky130_fd_sc_hd__nand2_1
X_10054_ _09617_/C _09617_/B _09612_/Y vssd1 vssd1 vccd1 vccd1 _10056_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09944__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06980_ _10212_/B _10112_/A vssd1 vssd1 vccd1 vccd1 _07144_/B sky130_fd_sc_hd__nand2_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05931_ _05933_/C vssd1 vssd1 vccd1 vccd1 _05932_/B sky130_fd_sc_hd__inv_2
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08650_ _08650_/A vssd1 vssd1 vccd1 vccd1 _08651_/B sky130_fd_sc_hd__inv_2
X_05862_ _06186_/A _06186_/B vssd1 vssd1 vccd1 vccd1 _06185_/A sky130_fd_sc_hd__nand2_1
X_07601_ _10452_/A _10447_/B _10453_/B vssd1 vssd1 vccd1 vccd1 _08386_/C sky130_fd_sc_hd__nand3_1
X_05793_ _05853_/C _05793_/B vssd1 vssd1 vccd1 vccd1 _05797_/A sky130_fd_sc_hd__nand2_1
X_08581_ _09135_/A _08581_/B vssd1 vssd1 vccd1 vccd1 _08583_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07532_ _07532_/A _07532_/B vssd1 vssd1 vccd1 vccd1 _07535_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07463_ _09517_/C _07891_/B vssd1 vssd1 vccd1 vccd1 _07620_/B sky130_fd_sc_hd__nand2_1
X_09202_ _09201_/A _10188_/A _09201_/C vssd1 vssd1 vccd1 vccd1 _09203_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__06527__B _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06414_ _06427_/B _06289_/Y _06290_/Y vssd1 vssd1 vccd1 vccd1 _06415_/B sky130_fd_sc_hd__a21o_1
X_09133_ _09133_/A _09133_/B vssd1 vssd1 vccd1 vccd1 _09296_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07394_ _07561_/A _07394_/B vssd1 vssd1 vccd1 vccd1 _07450_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06345_ _06333_/Y _06468_/B _06344_/Y vssd1 vssd1 vccd1 vccd1 _06477_/A sky130_fd_sc_hd__a21oi_1
X_09064_ _09327_/A _09328_/C vssd1 vssd1 vccd1 vccd1 _09064_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_44_387 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06276_ _06440_/C _06440_/B _06275_/Y vssd1 vssd1 vccd1 vccd1 _06431_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_4_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08015_ _07991_/C _07991_/B _07985_/A vssd1 vssd1 vccd1 vccd1 _08030_/A sky130_fd_sc_hd__a21oi_2
X_09966_ _09966_/A _09966_/B vssd1 vssd1 vccd1 vccd1 _09988_/C sky130_fd_sc_hd__nand2_1
X_08917_ _08917_/A _08917_/B vssd1 vssd1 vccd1 vccd1 _08925_/C sky130_fd_sc_hd__nand2_1
X_09897_ _09895_/Y _09732_/B _09896_/Y vssd1 vssd1 vccd1 vccd1 _10319_/A sky130_fd_sc_hd__a21oi_2
X_08848_ _08859_/A _08859_/C vssd1 vssd1 vccd1 vccd1 _08858_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05606__B input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08779_ _08781_/C vssd1 vssd1 vccd1 vccd1 _08779_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_79_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10741_ _10741_/CLK hold6/X input65/X vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05341__B _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10672_ _10672_/A _10672_/B vssd1 vssd1 vccd1 vccd1 _10675_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10106_ _10106_/A _10106_/B vssd1 vssd1 vccd1 vccd1 _10107_/A sky130_fd_sc_hd__xor2_1
X_10037_ _10037_/A vssd1 vssd1 vccd1 vccd1 _10259_/B sky130_fd_sc_hd__inv_2
XFILLER_0_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06628__A _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06347__B _07646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06130_ _08101_/B input4/X vssd1 vssd1 vccd1 vccd1 _06282_/C sky130_fd_sc_hd__nand2_1
X_06061_ _06071_/A _06071_/B vssd1 vssd1 vccd1 vccd1 _06070_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07178__B _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09820_ _09824_/B _09835_/A vssd1 vssd1 vccd1 vccd1 _09823_/A sky130_fd_sc_hd__nand2_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09751_ _09752_/A _09751_/B vssd1 vssd1 vccd1 vccd1 _09839_/A sky130_fd_sc_hd__nand2b_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06963_ _06965_/A _06965_/B vssd1 vssd1 vccd1 vccd1 _06964_/A sky130_fd_sc_hd__nand2_1
X_08702_ _08707_/A _09229_/A vssd1 vssd1 vccd1 vccd1 _09247_/B sky130_fd_sc_hd__nand2_1
X_05914_ _05474_/C _05474_/B _05913_/Y vssd1 vssd1 vccd1 vccd1 _06711_/A sky130_fd_sc_hd__a21oi_2
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09682_ _09683_/B _09683_/A vssd1 vssd1 vccd1 vccd1 _10003_/A sky130_fd_sc_hd__or2_1
X_06894_ _06894_/A _06894_/B vssd1 vssd1 vccd1 vccd1 _06896_/A sky130_fd_sc_hd__nand2_1
X_08633_ _09912_/A _08633_/B _08633_/C vssd1 vssd1 vccd1 vccd1 _08633_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_55_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05845_ _09778_/D input1/X _09477_/C _09698_/A vssd1 vssd1 vccd1 vccd1 _05846_/A
+ sky130_fd_sc_hd__and4_1
X_08564_ _08884_/C _08878_/B vssd1 vssd1 vccd1 vccd1 _08567_/A sky130_fd_sc_hd__nand2_1
X_05776_ _05854_/A _05855_/A vssd1 vssd1 vccd1 vccd1 _05776_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_49_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07515_ _07519_/B _07516_/A vssd1 vssd1 vccd1 vccd1 _07518_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_479 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08495_ _08573_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _08498_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07446_ _07446_/A _07446_/B _07446_/C vssd1 vssd1 vccd1 vccd1 _07713_/C sky130_fd_sc_hd__nand3_1
X_07377_ _07222_/Y _07377_/B _07377_/C vssd1 vssd1 vccd1 vccd1 _07449_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09116_ _08925_/C _08925_/B _08916_/Y vssd1 vssd1 vccd1 vccd1 _09118_/A sky130_fd_sc_hd__a21oi_1
XANTENNA__06273__A _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06328_ _06454_/A _06455_/B vssd1 vssd1 vccd1 vccd1 _06458_/C sky130_fd_sc_hd__nand2_1
X_09047_ _09039_/Y _09058_/B _09046_/Y vssd1 vssd1 vccd1 vccd1 _09069_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_44_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07088__B _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06259_ _06259_/A _06259_/B _06259_/C vssd1 vssd1 vccd1 vccd1 _06260_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06720__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ _09624_/B _10115_/A input21/X _09622_/X vssd1 vssd1 vccd1 vccd1 _09950_/A
+ sky130_fd_sc_hd__a31o_1
XANTENNA__08128__A2 _09971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09876__A2 _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08647__B _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10724_ _10724_/CLK _10724_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10655_ _10654_/A _10653_/A _10502_/B vssd1 vssd1 vccd1 vccd1 _10657_/A sky130_fd_sc_hd__o21ai_1
X_10586_ _10588_/B hold15/A vssd1 vssd1 vccd1 vccd1 _10587_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05630_ _05892_/B _05630_/B vssd1 vssd1 vccd1 vccd1 _05632_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10739__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05561_ _05564_/A _05564_/C vssd1 vssd1 vccd1 vccd1 _05563_/A sky130_fd_sc_hd__nand2_1
X_07300_ _07300_/A _07300_/B vssd1 vssd1 vccd1 vccd1 _07432_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_73_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05492_ _05492_/A vssd1 vssd1 vccd1 vccd1 _05493_/B sky130_fd_sc_hd__inv_2
X_08280_ _08280_/A _08280_/B vssd1 vssd1 vccd1 vccd1 _08281_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08573__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07231_ _07398_/B vssd1 vssd1 vccd1 vccd1 _07232_/B sky130_fd_sc_hd__inv_2
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07162_ _07187_/A _07187_/B vssd1 vssd1 vccd1 vccd1 _07167_/C sky130_fd_sc_hd__nand2_1
X_06113_ _06113_/A _06113_/B _06113_/C vssd1 vssd1 vccd1 vccd1 _06118_/A sky130_fd_sc_hd__nand3_1
X_07093_ _07230_/B _07228_/A vssd1 vssd1 vccd1 vccd1 _07414_/A sky130_fd_sc_hd__and2_1
XFILLER_0_14_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06044_ _06044_/A _06890_/B vssd1 vssd1 vccd1 vccd1 _06075_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09803_ _09803_/A _09803_/B vssd1 vssd1 vccd1 vccd1 _10083_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07995_ _07995_/A vssd1 vssd1 vccd1 vccd1 _07996_/B sky130_fd_sc_hd__inv_2
X_09734_ _09734_/A _09734_/B vssd1 vssd1 vccd1 vccd1 _09736_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06946_ _06948_/A _06948_/B vssd1 vssd1 vccd1 vccd1 _06947_/A sky130_fd_sc_hd__nand2_1
X_06877_ _06877_/A _06877_/B vssd1 vssd1 vccd1 vccd1 _06878_/B sky130_fd_sc_hd__nand2_1
X_09665_ _09665_/A _09665_/B vssd1 vssd1 vccd1 vccd1 _09667_/A sky130_fd_sc_hd__nand2_1
X_05828_ _05832_/B _06091_/B vssd1 vssd1 vccd1 vccd1 _05831_/A sky130_fd_sc_hd__nand2_1
X_08616_ _08616_/A _08616_/B _09210_/A vssd1 vssd1 vccd1 vccd1 _08618_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_82_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09596_ _09596_/A _09596_/B vssd1 vssd1 vccd1 vccd1 _09597_/B sky130_fd_sc_hd__nand2_1
X_05759_ input41/X vssd1 vssd1 vccd1 vccd1 _10187_/B sky130_fd_sc_hd__clkbuf_8
X_08547_ _08547_/A _08570_/B _08547_/C vssd1 vssd1 vccd1 vccd1 _08570_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08478_ _08478_/A _08478_/B vssd1 vssd1 vccd1 vccd1 _08491_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08483__A _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07429_ _07429_/A _07429_/B vssd1 vssd1 vccd1 vccd1 _07572_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10440_ _10440_/A _10440_/B vssd1 vssd1 vccd1 vccd1 _10441_/A sky130_fd_sc_hd__nand2_1
X_10371_ _10560_/A hold54/X _10560_/B vssd1 vssd1 vccd1 vccd1 _10697_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_32_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09745__C _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10707_ _10707_/A _10707_/B vssd1 vssd1 vccd1 vccd1 _10708_/A sky130_fd_sc_hd__or2_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10638_ _10638_/A _10638_/B vssd1 vssd1 vccd1 vccd1 _10639_/B sky130_fd_sc_hd__nand2_1
X_10569_ _10569_/A _10569_/B _10569_/C vssd1 vssd1 vccd1 vccd1 _10573_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_11_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_305 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07456__B _08453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06800_ _06800_/A _06800_/B _08442_/A vssd1 vssd1 vccd1 vccd1 _06801_/B sky130_fd_sc_hd__nand3_1
X_07780_ _07764_/B _07764_/C _07782_/B vssd1 vssd1 vccd1 vccd1 _07781_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_39_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06731_ _06731_/A _06731_/B vssd1 vssd1 vccd1 vccd1 _06737_/B sky130_fd_sc_hd__nand2_1
Xinput4 a_i[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_4
X_09450_ _09450_/A _09450_/B vssd1 vssd1 vccd1 vccd1 _09510_/B sky130_fd_sc_hd__nand2_1
X_08401_ _10156_/A _10004_/A vssd1 vssd1 vccd1 vccd1 _08447_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_2_1__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _10718_/CLK sky130_fd_sc_hd__clkbuf_16
X_06662_ _06665_/B _06665_/C vssd1 vssd1 vccd1 vccd1 _06663_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05704__B _06228_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05613_ _08725_/A input38/X vssd1 vssd1 vccd1 vccd1 _05615_/A sky130_fd_sc_hd__nand2_1
X_09381_ _09381_/A _09381_/B vssd1 vssd1 vccd1 vccd1 _09382_/B sky130_fd_sc_hd__and2_1
X_06593_ _07096_/B _07096_/A vssd1 vssd1 vccd1 vccd1 _07079_/A sky130_fd_sc_hd__nor2_1
X_05544_ input31/X vssd1 vssd1 vccd1 vccd1 _08724_/A sky130_fd_sc_hd__buf_6
X_08332_ _08332_/A _08346_/B vssd1 vssd1 vccd1 vccd1 _08349_/B sky130_fd_sc_hd__nand2_1
X_08263_ _08331_/A vssd1 vssd1 vccd1 vccd1 _08299_/B sky130_fd_sc_hd__inv_2
XANTENNA__10338__A _10338_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05475_ _05480_/B _05480_/C vssd1 vssd1 vccd1 vccd1 _05898_/B sky130_fd_sc_hd__nand2_1
X_07214_ _07214_/A _07214_/B vssd1 vssd1 vccd1 vccd1 _07215_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06535__B _07646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08194_ _08194_/A vssd1 vssd1 vccd1 vccd1 _08272_/A sky130_fd_sc_hd__inv_2
X_07145_ _07145_/A _07145_/B _07145_/C vssd1 vssd1 vccd1 vccd1 _07312_/B sky130_fd_sc_hd__nand3_1
X_07076_ _07074_/Y _07067_/B _07075_/Y vssd1 vssd1 vccd1 vccd1 _07084_/A sky130_fd_sc_hd__a21oi_1
X_06027_ _06027_/A _06027_/B vssd1 vssd1 vccd1 vccd1 _06841_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06270__B _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07978_ _07978_/A _07978_/B vssd1 vssd1 vccd1 vccd1 _08037_/B sky130_fd_sc_hd__nand2_1
X_09717_ _09717_/A vssd1 vssd1 vccd1 vccd1 _09718_/B sky130_fd_sc_hd__inv_2
X_06929_ _06929_/A _09325_/A _06930_/B vssd1 vssd1 vccd1 vccd1 _09353_/A sky130_fd_sc_hd__nand3_2
XANTENNA__07382__A _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__A1 _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__B2 _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ _10130_/A _10128_/B _10129_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _09649_/B
+ sky130_fd_sc_hd__a22o_1
X_09579_ _09579_/A _09821_/B _09579_/C vssd1 vssd1 vccd1 vccd1 _09821_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06726__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06445__B _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10423_ _10423_/A _10423_/B vssd1 vssd1 vccd1 vccd1 _10557_/A sky130_fd_sc_hd__nor2_1
X_10354_ _10357_/A _10357_/C vssd1 vssd1 vccd1 vccd1 _10375_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09519__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09519__B2 _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10285_ _10285_/A _10285_/B vssd1 vssd1 vccd1 vccd1 _10290_/C sky130_fd_sc_hd__nand2_1
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05805__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09455__B1 _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10158__A _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08851__A _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08950_ _08938_/B _08950_/B vssd1 vssd1 vccd1 vccd1 _09005_/B sky130_fd_sc_hd__nand2b_1
X_08881_ _08881_/A _08881_/B vssd1 vssd1 vccd1 vccd1 _08884_/B sky130_fd_sc_hd__nand2_1
X_07901_ _07935_/A _07936_/C vssd1 vssd1 vccd1 vccd1 _07976_/A sky130_fd_sc_hd__nand2_1
X_07832_ _08087_/B vssd1 vssd1 vccd1 vccd1 _08083_/B sky130_fd_sc_hd__inv_2
X_09502_ _09502_/A _09502_/B _09793_/A vssd1 vssd1 vccd1 vccd1 _09506_/C sky130_fd_sc_hd__nand3_1
X_07763_ _07763_/A vssd1 vssd1 vccd1 vccd1 _07764_/B sky130_fd_sc_hd__inv_2
X_06714_ _08171_/B _10151_/B vssd1 vssd1 vccd1 vccd1 _06718_/A sky130_fd_sc_hd__nand2_1
X_07694_ _07735_/A _07734_/B vssd1 vssd1 vccd1 vccd1 _07733_/C sky130_fd_sc_hd__nand2_1
XANTENNA__05434__B _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09433_ _09433_/A _09433_/B vssd1 vssd1 vccd1 vccd1 _09439_/A sky130_fd_sc_hd__nand2_1
X_06645_ _06968_/A _06967_/A vssd1 vssd1 vccd1 vccd1 _06645_/Y sky130_fd_sc_hd__nor2_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09364_ _09365_/B _09365_/A vssd1 vssd1 vccd1 vccd1 _09369_/B sky130_fd_sc_hd__or2_1
XFILLER_0_59_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08315_ _08315_/A _08316_/B _08315_/C vssd1 vssd1 vccd1 vccd1 _08334_/B sky130_fd_sc_hd__nand3_1
X_06576_ _06579_/A _06579_/C vssd1 vssd1 vccd1 vccd1 _06578_/A sky130_fd_sc_hd__nand2_1
X_09295_ _09294_/B _09512_/B _09295_/C vssd1 vssd1 vccd1 vccd1 _09512_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_34_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05527_ _05527_/A _05527_/B vssd1 vssd1 vccd1 vccd1 _05533_/B sky130_fd_sc_hd__nand2_1
X_08246_ _08246_/A _08287_/B vssd1 vssd1 vccd1 vccd1 _08285_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05458_ _05457_/B _05458_/B _05458_/C vssd1 vssd1 vccd1 vccd1 _05459_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_15_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ _08177_/A _08176_/Y vssd1 vssd1 vccd1 vccd1 _08251_/C sky130_fd_sc_hd__or2b_1
XFILLER_0_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07128_ _07147_/C _07147_/B _06984_/Y vssd1 vssd1 vccd1 vccd1 _07137_/B sky130_fd_sc_hd__a21o_1
X_05389_ _05634_/B _05634_/C vssd1 vssd1 vccd1 vccd1 _05636_/B sky130_fd_sc_hd__nand2_1
X_07059_ _07203_/A _07203_/B vssd1 vssd1 vccd1 vccd1 _07064_/A sky130_fd_sc_hd__nand2_1
X_10070_ _10070_/A _10070_/B vssd1 vssd1 vccd1 vccd1 _10073_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08001__A _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05360__A _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10406_ _10406_/A _10406_/B vssd1 vssd1 vccd1 vccd1 _10415_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06191__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10337_ _10337_/A _10338_/A vssd1 vssd1 vccd1 vccd1 _10343_/A sky130_fd_sc_hd__nand2_1
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10268_ _10272_/A _10272_/B vssd1 vssd1 vccd1 vccd1 _10271_/A sky130_fd_sc_hd__nand2_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10199_ _10199_/A _10199_/B vssd1 vssd1 vccd1 vccd1 _10220_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_17_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06430_ _06430_/A _06430_/B vssd1 vssd1 vccd1 vccd1 _06432_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06361_ _06361_/A _06361_/B _06361_/C vssd1 vssd1 vccd1 vccd1 _06365_/C sky130_fd_sc_hd__nand3_1
X_09080_ _09080_/A _09080_/B vssd1 vssd1 vccd1 vccd1 _09581_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09677__A _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08100_ _08100_/A _08100_/B vssd1 vssd1 vccd1 vccd1 _08104_/C sky130_fd_sc_hd__nand2_1
X_06292_ _06415_/A _06413_/A vssd1 vssd1 vccd1 vccd1 _06292_/Y sky130_fd_sc_hd__nand2_1
Xinput40 b_i[16] vssd1 vssd1 vccd1 vccd1 input40/X sky130_fd_sc_hd__buf_2
X_08031_ _08031_/A vssd1 vssd1 vccd1 vccd1 _08033_/A sky130_fd_sc_hd__inv_2
XFILLER_0_3_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput51 b_i[26] vssd1 vssd1 vccd1 vccd1 input51/X sky130_fd_sc_hd__buf_2
Xinput62 b_i[7] vssd1 vssd1 vccd1 vccd1 input62/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09982_ _09982_/A _09982_/B vssd1 vssd1 vccd1 vccd1 _09984_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08933_ _08933_/A vssd1 vssd1 vccd1 vccd1 _08939_/B sky130_fd_sc_hd__inv_2
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08864_ _08864_/A _08864_/B vssd1 vssd1 vccd1 vccd1 _08866_/A sky130_fd_sc_hd__nand2_1
X_08795_ _09268_/A _10276_/B _08795_/C vssd1 vssd1 vccd1 vccd1 _08798_/A sky130_fd_sc_hd__nor3_1
X_07815_ _07965_/B _07964_/A vssd1 vssd1 vccd1 vccd1 _07815_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__05445__A _07785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07746_ _10247_/B _08574_/A vssd1 vssd1 vccd1 vccd1 _07916_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10277__B2 _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10277__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09416_ _10158_/A _10157_/A _10150_/B _10151_/B vssd1 vssd1 vccd1 vccd1 _09417_/A
+ sky130_fd_sc_hd__and4_1
X_07677_ _07741_/A _07742_/A vssd1 vssd1 vccd1 vccd1 _07744_/B sky130_fd_sc_hd__nand2_1
X_06628_ _08574_/A _10201_/A vssd1 vssd1 vccd1 vccd1 _06974_/B sky130_fd_sc_hd__nand2_1
X_09347_ _09357_/B _10359_/A vssd1 vssd1 vccd1 vccd1 _09348_/B sky130_fd_sc_hd__nor2_1
X_06559_ _07034_/C vssd1 vssd1 vccd1 vccd1 _06560_/B sky130_fd_sc_hd__inv_2
XFILLER_0_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09278_ _09278_/A _09278_/B _09278_/C vssd1 vssd1 vccd1 vccd1 _09285_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08229_ _08373_/A _08229_/B vssd1 vssd1 vccd1 vccd1 _08376_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10122_ _10123_/B _10123_/A vssd1 vssd1 vccd1 vccd1 _10124_/A sky130_fd_sc_hd__or2_1
X_10053_ _10230_/A _10057_/B vssd1 vssd1 vccd1 vccd1 _10055_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_263 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05930_ _05930_/A _06755_/A vssd1 vssd1 vccd1 vccd1 _05933_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_28_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05861_ _05861_/A _05861_/B vssd1 vssd1 vccd1 vccd1 _06186_/A sky130_fd_sc_hd__nand2_1
X_07600_ _07600_/A _07851_/B vssd1 vssd1 vccd1 vccd1 _10447_/B sky130_fd_sc_hd__nand2_1
X_08580_ _08580_/A _09135_/A _08581_/B vssd1 vssd1 vccd1 vccd1 _09156_/B sky130_fd_sc_hd__nand3_1
X_05792_ _06020_/B _06020_/A vssd1 vssd1 vccd1 vccd1 _05794_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_44_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07531_ _07531_/A vssd1 vssd1 vccd1 vccd1 _07532_/B sky130_fd_sc_hd__inv_2
XFILLER_0_44_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07462_ _07544_/A _07545_/C vssd1 vssd1 vccd1 vccd1 _07543_/B sky130_fd_sc_hd__nand2_1
X_09201_ _09201_/A _10188_/A _09201_/C vssd1 vssd1 vccd1 vccd1 _09459_/A sky130_fd_sc_hd__nor3_1
X_07393_ _09551_/C _09201_/A _07391_/C vssd1 vssd1 vccd1 vccd1 _07394_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06413_ _06413_/A _06413_/B _06413_/C vssd1 vssd1 vccd1 vccd1 _06418_/A sky130_fd_sc_hd__nand3_1
X_09132_ _09302_/B vssd1 vssd1 vccd1 vccd1 _09300_/A sky130_fd_sc_hd__inv_2
XFILLER_0_60_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06344_ _06466_/A _06465_/A vssd1 vssd1 vccd1 vccd1 _06344_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__09200__A _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09063_ _09061_/Y _06918_/B _09062_/Y vssd1 vssd1 vccd1 vccd1 _09328_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_44_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06275_ _06436_/A _06437_/B vssd1 vssd1 vccd1 vccd1 _06275_/Y sky130_fd_sc_hd__nor2_1
X_08014_ _08018_/A _08018_/B vssd1 vssd1 vccd1 vccd1 _08030_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09965_ _09965_/A vssd1 vssd1 vccd1 vccd1 _09988_/A sky130_fd_sc_hd__inv_2
X_08916_ _08917_/B _08917_/A vssd1 vssd1 vccd1 vccd1 _08916_/Y sky130_fd_sc_hd__nor2_1
X_09896_ _09896_/A _09896_/B vssd1 vssd1 vccd1 vccd1 _09896_/Y sky130_fd_sc_hd__nor2_1
X_08847_ _08930_/B _08847_/B vssd1 vssd1 vccd1 vccd1 _08859_/C sky130_fd_sc_hd__nand2_1
X_08778_ _08815_/B _08815_/C vssd1 vssd1 vccd1 vccd1 _08805_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07390__A _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05903__A _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07729_ _07735_/A vssd1 vssd1 vccd1 vccd1 _07734_/A sky130_fd_sc_hd__inv_2
X_10740_ _10741_/CLK hold11/X fanout98/X vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__dfrtp_2
XFILLER_0_67_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10671_ _10672_/B _10672_/A vssd1 vssd1 vccd1 vccd1 _10673_/A sky130_fd_sc_hd__or2_1
XFILLER_0_35_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10105_ _10105_/A _10104_/X vssd1 vssd1 vccd1 vccd1 _10106_/B sky130_fd_sc_hd__or2b_1
X_10036_ _10036_/A _10037_/A vssd1 vssd1 vccd1 vccd1 _10048_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05813__A input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06628__B _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_174 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06060_ _06060_/A _06060_/B _06869_/A vssd1 vssd1 vccd1 vccd1 _06071_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09750_ _09752_/B vssd1 vssd1 vccd1 vccd1 _09751_/B sky130_fd_sc_hd__inv_2
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06962_ _06962_/A _06962_/B vssd1 vssd1 vccd1 vccd1 _06965_/B sky130_fd_sc_hd__nand2_1
X_08701_ _08701_/A _08701_/B vssd1 vssd1 vccd1 vccd1 _09229_/A sky130_fd_sc_hd__nand2_1
X_09681_ _10003_/B _09681_/B vssd1 vssd1 vccd1 vccd1 _09683_/A sky130_fd_sc_hd__nand2_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05913_ _05913_/A _05913_/B vssd1 vssd1 vccd1 vccd1 _05913_/Y sky130_fd_sc_hd__nor2_1
X_06893_ _06895_/C vssd1 vssd1 vccd1 vccd1 _06894_/B sky130_fd_sc_hd__inv_2
X_08632_ _10157_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _08633_/C sky130_fd_sc_hd__nand2_1
X_05844_ _05887_/A _05887_/B vssd1 vssd1 vccd1 vccd1 _05886_/A sky130_fd_sc_hd__nand2_1
X_08563_ _08878_/A _08563_/B _08878_/B vssd1 vssd1 vccd1 vccd1 _08884_/C sky130_fd_sc_hd__nand3_1
X_05775_ _06186_/B _05860_/A vssd1 vssd1 vccd1 vccd1 _05858_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_9_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07514_ _07517_/B vssd1 vssd1 vccd1 vccd1 _07519_/B sky130_fd_sc_hd__inv_2
X_08494_ _10115_/A input17/X vssd1 vssd1 vccd1 vccd1 _08501_/B sky130_fd_sc_hd__nand2_1
X_07445_ _07445_/A _07445_/B _07445_/C vssd1 vssd1 vccd1 vccd1 _07446_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_57_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07376_ _07222_/Y _07375_/Y _07221_/A vssd1 vssd1 vccd1 vccd1 _07449_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_17_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09115_ _09119_/B _09544_/A vssd1 vssd1 vccd1 vccd1 _09117_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06327_ _08337_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _06455_/B sky130_fd_sc_hd__nand2_1
X_09046_ _09056_/A _09055_/A vssd1 vssd1 vccd1 vccd1 _09046_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_4_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06273__B _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06258_ _06258_/A _06258_/B vssd1 vssd1 vccd1 vccd1 _06260_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06189_ _06188_/B _06189_/B _06189_/C vssd1 vssd1 vccd1 vccd1 _06217_/C sky130_fd_sc_hd__nand3b_1
X_09948_ _09948_/A _10109_/A vssd1 vssd1 vccd1 vccd1 _09952_/B sky130_fd_sc_hd__nand2_1
X_09879_ _09782_/A _09551_/C _09877_/Y vssd1 vssd1 vccd1 vccd1 _09880_/B sky130_fd_sc_hd__o21ai_1
X_10723_ _10724_/CLK hold38/X fanout99/X vssd1 vssd1 vccd1 vccd1 hold62/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10654_ _10654_/A hold47/X vssd1 vssd1 vccd1 vccd1 hold48/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_130 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10585_ hold15/X _10588_/B vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__xor2_1
XFILLER_0_50_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05808__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10019_ _10184_/A _10019_/B _10019_/C vssd1 vssd1 vccd1 vccd1 _10183_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_58_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05560_ _05560_/A _05560_/B _05560_/C vssd1 vssd1 vccd1 vccd1 _05564_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_18_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05491_ _05491_/A _05492_/A vssd1 vssd1 vccd1 vccd1 _05494_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07230_ _07230_/A _07230_/B vssd1 vssd1 vccd1 vccd1 _07398_/B sky130_fd_sc_hd__nand2_1
X_07161_ _07161_/A _07161_/B vssd1 vssd1 vccd1 vccd1 _07167_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_54_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06112_ _06493_/B _06493_/C vssd1 vssd1 vccd1 vccd1 _06495_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07092_ _07229_/B _07228_/A _07228_/B vssd1 vssd1 vccd1 vccd1 _07230_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06043_ _06045_/B _06045_/C vssd1 vssd1 vccd1 vccd1 _06890_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05718__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09802_ _09804_/B vssd1 vssd1 vccd1 vccd1 _09803_/B sky130_fd_sc_hd__inv_2
XFILLER_0_5_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07994_ _07994_/A vssd1 vssd1 vccd1 vccd1 _07996_/A sky130_fd_sc_hd__inv_2
X_09733_ _09732_/B _09733_/B _09733_/C vssd1 vssd1 vccd1 vccd1 _09734_/B sky130_fd_sc_hd__nand3b_1
X_06945_ _06945_/A _06945_/B vssd1 vssd1 vccd1 vccd1 _06948_/B sky130_fd_sc_hd__nand2_1
X_06876_ _06876_/A _08951_/B vssd1 vssd1 vccd1 vccd1 _06877_/A sky130_fd_sc_hd__nand2_1
X_09664_ _09664_/A vssd1 vssd1 vccd1 vccd1 _09665_/B sky130_fd_sc_hd__inv_2
X_05827_ _05826_/B _05827_/B _06057_/A vssd1 vssd1 vccd1 vccd1 _06091_/B sky130_fd_sc_hd__nand3b_1
X_09595_ _09596_/B _09596_/A vssd1 vssd1 vccd1 vccd1 _09918_/A sky130_fd_sc_hd__or2_1
X_08615_ _09210_/B _08615_/B vssd1 vssd1 vccd1 vccd1 _08618_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08546_ _08546_/A vssd1 vssd1 vccd1 vccd1 _08547_/A sky130_fd_sc_hd__inv_2
X_05758_ input26/X vssd1 vssd1 vccd1 vccd1 _09517_/D sky130_fd_sc_hd__buf_12
XFILLER_0_49_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08477_ _08491_/A _08491_/C vssd1 vssd1 vccd1 vccd1 _08480_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05689_ _06264_/A _06265_/B vssd1 vssd1 vccd1 vccd1 _06268_/C sky130_fd_sc_hd__nand2_1
X_07428_ _07430_/A _07430_/B vssd1 vssd1 vccd1 vccd1 _07429_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10518__B _10638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07359_ _09840_/B _10128_/A vssd1 vssd1 vccd1 vccd1 _07453_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10370_ _10370_/A _10370_/B vssd1 vssd1 vccd1 vccd1 _10560_/A sky130_fd_sc_hd__or2_1
XFILLER_0_32_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09029_ _09069_/A _09069_/C vssd1 vssd1 vccd1 vccd1 _09068_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09745__D _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08004__A _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10706_ _10706_/A _10706_/B vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06194__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10637_ hold5/X _10637_/B vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10568_ _10596_/B _10604_/B vssd1 vssd1 vccd1 vccd1 _10707_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10499_ _10653_/B vssd1 vssd1 vccd1 vccd1 _10499_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_11_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08849__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 a_i[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_4
X_06730_ _10115_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _06731_/B sky130_fd_sc_hd__nand2_1
X_06661_ _06661_/A _06661_/B vssd1 vssd1 vccd1 vccd1 _06665_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_78_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08400_ _09912_/A _10188_/A _08403_/C vssd1 vssd1 vccd1 vccd1 _08445_/B sky130_fd_sc_hd__o21ai_1
X_05612_ _05616_/A _05616_/C vssd1 vssd1 vccd1 vccd1 _05614_/A sky130_fd_sc_hd__nand2_1
X_09380_ _09383_/B _09641_/A vssd1 vssd1 vccd1 vccd1 _09382_/A sky130_fd_sc_hd__nand2_1
X_06592_ _07062_/B _07060_/A vssd1 vssd1 vccd1 vccd1 _07096_/A sky130_fd_sc_hd__and2_1
XFILLER_0_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05543_ _05547_/A _05547_/B vssd1 vssd1 vccd1 vccd1 _05716_/C sky130_fd_sc_hd__nand2_1
X_08331_ _08331_/A _08331_/B vssd1 vssd1 vccd1 vccd1 _08332_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05474_ _05474_/A _05474_/B _05474_/C vssd1 vssd1 vccd1 vccd1 _05480_/C sky130_fd_sc_hd__nand3_1
X_08262_ _09840_/B _10292_/B _10103_/A _10103_/B vssd1 vssd1 vccd1 vccd1 _08331_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_61_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07213_ _07213_/A _07213_/B _07213_/C vssd1 vssd1 vccd1 vccd1 _07226_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_14_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08193_ _08193_/A _08193_/B vssd1 vssd1 vccd1 vccd1 _08194_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06832__A _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07144_ _07146_/A _07144_/B vssd1 vssd1 vccd1 vccd1 _07145_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07075_ _07075_/A _07075_/B vssd1 vssd1 vccd1 vccd1 _07075_/Y sky130_fd_sc_hd__nor2_1
X_06026_ _06028_/B vssd1 vssd1 vccd1 vccd1 _06027_/B sky130_fd_sc_hd__inv_2
XFILLER_0_77_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07977_ _08045_/A _08046_/C vssd1 vssd1 vccd1 vccd1 _07978_/A sky130_fd_sc_hd__nand2_1
X_09716_ _09716_/A _09717_/A vssd1 vssd1 vccd1 vccd1 _09719_/A sky130_fd_sc_hd__nand2_1
X_06928_ _06928_/A _06928_/B _06928_/C vssd1 vssd1 vccd1 vccd1 _06930_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07382__B _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09700__A2 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06859_ _10210_/A _08897_/B vssd1 vssd1 vccd1 vccd1 _06860_/B sky130_fd_sc_hd__nand2_1
X_09647_ _09647_/A vssd1 vssd1 vccd1 vccd1 _09982_/B sky130_fd_sc_hd__inv_2
X_09578_ _09578_/A _09578_/B vssd1 vssd1 vccd1 vccd1 _09584_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08494__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08529_ _09971_/A _08529_/B _08529_/C vssd1 vssd1 vccd1 vccd1 _08604_/B sky130_fd_sc_hd__or3_1
XFILLER_0_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06726__B _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_228 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10422_ _10555_/A _10685_/B vssd1 vssd1 vccd1 vccd1 _10423_/B sky130_fd_sc_hd__nor2_1
X_10353_ _10376_/A _10353_/B _10353_/C vssd1 vssd1 vccd1 vccd1 _10357_/C sky130_fd_sc_hd__nand3_1
XANTENNA__09519__A2 _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05358__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10284_ input56/X _10284_/B vssd1 vssd1 vccd1 vccd1 _10285_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05805__B _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09455__A1 _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09455__B2 _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10158__B _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08851__B _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08880_ _08884_/A _08884_/C vssd1 vssd1 vccd1 vccd1 _08883_/A sky130_fd_sc_hd__nand2_1
X_07900_ _08018_/B _07900_/B vssd1 vssd1 vccd1 vccd1 _07936_/C sky130_fd_sc_hd__nand2_1
X_07831_ _07831_/A _08075_/A _08075_/B vssd1 vssd1 vccd1 vccd1 _08087_/B sky130_fd_sc_hd__nand3_4
X_09501_ _09793_/B _09501_/B vssd1 vssd1 vccd1 vccd1 _09506_/B sky130_fd_sc_hd__nand2_1
X_07762_ _07762_/A _07763_/A vssd1 vssd1 vccd1 vccd1 _07765_/A sky130_fd_sc_hd__nand2_1
X_06713_ _06768_/A vssd1 vssd1 vccd1 vccd1 _06767_/B sky130_fd_sc_hd__inv_2
X_07693_ _07800_/C _07799_/B _07692_/Y vssd1 vssd1 vccd1 vccd1 _07734_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06827__A _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09432_ _09432_/A _09432_/B vssd1 vssd1 vccd1 vccd1 _09433_/B sky130_fd_sc_hd__nand2_1
X_06644_ _06969_/C vssd1 vssd1 vccd1 vccd1 _06960_/C sky130_fd_sc_hd__inv_2
XFILLER_0_59_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06575_ _06575_/A vssd1 vssd1 vccd1 vccd1 _06579_/A sky130_fd_sc_hd__inv_2
XANTENNA__10723__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09363_ _09361_/X _09363_/B vssd1 vssd1 vccd1 vccd1 _09365_/A sky130_fd_sc_hd__nand2b_1
X_08314_ _08314_/A vssd1 vssd1 vccd1 vccd1 _08315_/C sky130_fd_sc_hd__inv_2
X_05526_ _05525_/B _05526_/B _05526_/C vssd1 vssd1 vccd1 vccd1 _05527_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_74_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09294_ _09294_/A _09294_/B vssd1 vssd1 vccd1 vccd1 _09297_/A sky130_fd_sc_hd__nand2_1
X_08245_ _08245_/A _08245_/B vssd1 vssd1 vccd1 vccd1 _08246_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05457_ _05457_/A _05457_/B vssd1 vssd1 vccd1 vccd1 _05459_/A sky130_fd_sc_hd__nand2_1
X_08176_ _08897_/B _10101_/A vssd1 vssd1 vccd1 vccd1 _08176_/Y sky130_fd_sc_hd__nand2_1
X_05388_ _05388_/A _05388_/B _05388_/C vssd1 vssd1 vccd1 vccd1 _05634_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07127_ _07127_/A _07127_/B _07127_/C vssd1 vssd1 vccd1 vccd1 _07135_/A sky130_fd_sc_hd__nand3_1
X_07058_ _07058_/A _07065_/C _07065_/B vssd1 vssd1 vccd1 vccd1 _07203_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06009_ _06008_/B _06009_/B _06009_/C vssd1 vssd1 vccd1 vccd1 _06010_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__08001__B _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05641__A _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05360__B _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10405_ _10414_/A _10414_/C vssd1 vssd1 vccd1 vccd1 _10406_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06191__B input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10336_ _10336_/A _10336_/B vssd1 vssd1 vccd1 vccd1 _10338_/A sky130_fd_sc_hd__nand2_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10267_ _10266_/B _10267_/B _10267_/C vssd1 vssd1 vccd1 vccd1 _10272_/B sky130_fd_sc_hd__nand3b_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08399__A _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10198_ _10198_/A _10198_/B vssd1 vssd1 vccd1 vccd1 _10199_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05551__A _08453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06360_ _06360_/A _06360_/B vssd1 vssd1 vccd1 vccd1 _06361_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09677__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06291_ _06427_/B _06289_/Y _06290_/Y vssd1 vssd1 vccd1 vccd1 _06413_/A sky130_fd_sc_hd__a21oi_1
X_08030_ _08030_/A _08030_/B vssd1 vssd1 vccd1 vccd1 _08031_/A sky130_fd_sc_hd__or2_1
Xinput30 a_i[7] vssd1 vssd1 vccd1 vccd1 input30/X sky130_fd_sc_hd__clkbuf_1
Xinput52 b_i[27] vssd1 vssd1 vccd1 vccd1 input52/X sky130_fd_sc_hd__clkbuf_4
Xinput41 b_i[17] vssd1 vssd1 vccd1 vccd1 input41/X sky130_fd_sc_hd__buf_1
Xinput63 b_i[8] vssd1 vssd1 vccd1 vccd1 input63/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09981_ _09981_/A _09981_/B vssd1 vssd1 vccd1 vccd1 _09984_/C sky130_fd_sc_hd__nand2_1
X_08932_ _08937_/B _08937_/A vssd1 vssd1 vccd1 vccd1 _08933_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08863_ _08840_/C _08839_/A _08980_/A vssd1 vssd1 vccd1 vccd1 _08864_/B sky130_fd_sc_hd__o21ai_1
X_08794_ _10211_/A _09749_/B vssd1 vssd1 vccd1 vccd1 _08795_/C sky130_fd_sc_hd__nand2_1
X_07814_ _07872_/C _07872_/B _07813_/Y vssd1 vssd1 vccd1 vccd1 _07964_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__05445__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07745_ _07769_/A _07768_/B vssd1 vssd1 vccd1 vccd1 _07753_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10277__A2 _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09415_ _09415_/A vssd1 vssd1 vccd1 vccd1 _09421_/B sky130_fd_sc_hd__inv_2
X_07676_ _10040_/B input55/X vssd1 vssd1 vccd1 vccd1 _07742_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06627_ _08573_/A _09677_/A vssd1 vssd1 vccd1 vccd1 _06973_/A sky130_fd_sc_hd__nand2_1
X_09346_ _10389_/B _10385_/B vssd1 vssd1 vccd1 vccd1 _10359_/A sky130_fd_sc_hd__nand2_1
X_06558_ _06558_/A _06558_/B vssd1 vssd1 vccd1 vccd1 _07034_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_35_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09277_ _09277_/A _09277_/B vssd1 vssd1 vccd1 vccd1 _09285_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_62_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06489_ _06489_/A _06489_/B vssd1 vssd1 vccd1 vccd1 _06692_/B sky130_fd_sc_hd__nand2_1
X_05509_ _05509_/A _05509_/B vssd1 vssd1 vccd1 vccd1 _05954_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08228_ _08228_/A _08362_/B vssd1 vssd1 vccd1 vccd1 _08229_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_15_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08159_ _08162_/A _08162_/B vssd1 vssd1 vccd1 vccd1 _08254_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10121_ _10121_/A _10121_/B vssd1 vssd1 vccd1 vccd1 _10123_/A sky130_fd_sc_hd__nand2_1
X_10052_ _10052_/A _10052_/B _10052_/C vssd1 vssd1 vccd1 vccd1 _10057_/B sky130_fd_sc_hd__nand3_1
XANTENNA__05371__A _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09778__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10319_ _10319_/A _10319_/B vssd1 vssd1 vccd1 vccd1 _10321_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05860_ _05860_/A _05860_/B vssd1 vssd1 vccd1 vccd1 _05861_/A sky130_fd_sc_hd__nand2_1
X_05791_ _05796_/A _06040_/A vssd1 vssd1 vccd1 vccd1 _06020_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07761__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07530_ _07530_/A vssd1 vssd1 vccd1 vccd1 _07532_/A sky130_fd_sc_hd__inv_2
XFILLER_0_48_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07461_ _07535_/C _07535_/B _07460_/Y vssd1 vssd1 vccd1 vccd1 _07545_/C sky130_fd_sc_hd__a21oi_2
X_09200_ _10150_/A _10187_/A vssd1 vssd1 vccd1 vccd1 _09201_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_56_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07392_ _07392_/A vssd1 vssd1 vccd1 vccd1 _07561_/A sky130_fd_sc_hd__inv_2
X_06412_ _06679_/C vssd1 vssd1 vccd1 vccd1 _06678_/B sky130_fd_sc_hd__inv_2
X_09131_ _09131_/A _09576_/A vssd1 vssd1 vccd1 vccd1 _09302_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_56_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06343_ _06652_/B _06343_/B vssd1 vssd1 vccd1 vccd1 _06468_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09062_ _09062_/A _09062_/B vssd1 vssd1 vccd1 vccd1 _09062_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_44_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09200__B _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06274_ _06438_/C vssd1 vssd1 vccd1 vccd1 _06440_/B sky130_fd_sc_hd__inv_2
XFILLER_0_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08013_ _07900_/B _07899_/B _07899_/C vssd1 vssd1 vccd1 vccd1 _08018_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09964_ _09966_/B _09966_/A vssd1 vssd1 vccd1 vccd1 _09965_/A sky130_fd_sc_hd__nor2_1
X_08915_ _08802_/B _08802_/C _08802_/A vssd1 vssd1 vccd1 vccd1 _08917_/A sky130_fd_sc_hd__a21boi_1
X_09895_ _09896_/B _09896_/A vssd1 vssd1 vccd1 vccd1 _09895_/Y sky130_fd_sc_hd__nand2_1
X_08846_ _08846_/A _08846_/B vssd1 vssd1 vccd1 vccd1 _08930_/B sky130_fd_sc_hd__nand2_1
X_08777_ _08777_/A _08806_/A _08777_/C vssd1 vssd1 vccd1 vccd1 _08815_/C sky130_fd_sc_hd__nand3_1
X_05989_ _05989_/A vssd1 vssd1 vccd1 vccd1 _05995_/A sky130_fd_sc_hd__inv_2
XANTENNA__07390__B _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07728_ _07963_/B _07963_/C vssd1 vssd1 vccd1 vccd1 _07965_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05903__B _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07659_ _07660_/B _07659_/B _07659_/C vssd1 vssd1 vccd1 vccd1 _07669_/A sky130_fd_sc_hd__nand3_1
X_10670_ _10548_/B _10663_/A _10463_/B vssd1 vssd1 vccd1 vccd1 _10672_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_75_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09329_ _09331_/A _09331_/B vssd1 vssd1 vccd1 vccd1 _09330_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06750__A _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10104_ _10103_/A input25/X _10103_/B input20/X vssd1 vssd1 vccd1 vccd1 _10104_/X
+ sky130_fd_sc_hd__a22o_1
X_10035_ _10035_/A _10035_/B vssd1 vssd1 vccd1 vccd1 _10037_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08677__A _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05813__B _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07756__A _07756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06961_ _07127_/B _06961_/B vssd1 vssd1 vccd1 vccd1 _06962_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09971__A _09971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08700_ _08701_/B _08701_/A vssd1 vssd1 vccd1 vccd1 _08707_/A sky130_fd_sc_hd__or2_1
X_09680_ _10004_/A _10005_/A _10187_/A _09678_/C vssd1 vssd1 vccd1 vccd1 _09681_/B
+ sky130_fd_sc_hd__a22o_1
X_05912_ _05917_/A _06734_/A vssd1 vssd1 vccd1 vccd1 _06711_/B sky130_fd_sc_hd__nand2_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06892_ _06892_/A _06892_/B vssd1 vssd1 vccd1 vccd1 _06895_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_55_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08631_ _08629_/Y _08542_/B _08630_/Y vssd1 vssd1 vccd1 vccd1 _09281_/B sky130_fd_sc_hd__a21oi_2
XFILLER_0_55_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05843_ _05843_/A _05843_/B _05843_/C vssd1 vssd1 vccd1 vccd1 _05887_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08562_ _08562_/A _08562_/B _08562_/C vssd1 vssd1 vccd1 vccd1 _08878_/B sky130_fd_sc_hd__nand3_1
X_05774_ _05861_/B _05860_/A _05860_/B vssd1 vssd1 vccd1 vccd1 _06186_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_49_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08493_ _08562_/C _08549_/B vssd1 vssd1 vccd1 vccd1 _08522_/A sky130_fd_sc_hd__nand2_1
X_07513_ _07656_/B _07656_/C vssd1 vssd1 vccd1 vccd1 _07661_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07444_ _07444_/A _07444_/B vssd1 vssd1 vccd1 vccd1 _07446_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07375_ _07377_/C vssd1 vssd1 vccd1 vccd1 _07375_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09114_ _09544_/B _09114_/B _09114_/C vssd1 vssd1 vccd1 vccd1 _09544_/A sky130_fd_sc_hd__nand3_2
X_06326_ _08171_/B _09677_/A vssd1 vssd1 vccd1 vccd1 _06454_/A sky130_fd_sc_hd__nand2_1
X_09045_ _09071_/B _09044_/Y vssd1 vssd1 vccd1 vccd1 _09058_/B sky130_fd_sc_hd__nor2b_1
XFILLER_0_44_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06257_ _06428_/C vssd1 vssd1 vccd1 vccd1 _06427_/B sky130_fd_sc_hd__inv_2
XFILLER_0_4_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06188_ _06188_/A _06188_/B vssd1 vssd1 vccd1 vccd1 _06217_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_40_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09947_ _09947_/A _09947_/B vssd1 vssd1 vccd1 vccd1 _10109_/A sky130_fd_sc_hd__nand2_1
X_09878_ _09877_/Y input54/X _10284_/B vssd1 vssd1 vccd1 vccd1 _10280_/A sky130_fd_sc_hd__nand3b_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08829_ _08830_/B _08830_/A vssd1 vssd1 vccd1 vccd1 _08829_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10722_ _10724_/CLK _10722_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold36/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__09121__A input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10653_ _10653_/A _10653_/B vssd1 vssd1 vccd1 vccd1 hold47/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ _10584_/A _10584_/B vssd1 vssd1 vccd1 vccd1 _10588_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05808__B _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10018_ _10018_/A _10018_/B vssd1 vssd1 vccd1 vccd1 _10020_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05490_ _08101_/B _09922_/B vssd1 vssd1 vccd1 vccd1 _05492_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07160_ _07187_/B vssd1 vssd1 vccd1 vccd1 _07161_/B sky130_fd_sc_hd__inv_2
XFILLER_0_26_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06111_ _06111_/A _06111_/B _06111_/C vssd1 vssd1 vccd1 vccd1 _06493_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_14_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07091_ _07091_/A _07091_/B vssd1 vssd1 vccd1 vccd1 _07228_/B sky130_fd_sc_hd__nand2_1
X_06042_ _06041_/B _06042_/B _06042_/C vssd1 vssd1 vccd1 vccd1 _06045_/C sky130_fd_sc_hd__nand3b_1
XFILLER_0_14_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06390__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05718__B _07646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09801_ _09801_/A _09801_/B vssd1 vssd1 vccd1 vccd1 _09804_/B sky130_fd_sc_hd__nor2_1
X_09732_ _09732_/A _09732_/B vssd1 vssd1 vccd1 vccd1 _09734_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_76 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07993_ _08199_/C vssd1 vssd1 vccd1 vccd1 _08198_/B sky130_fd_sc_hd__inv_2
XFILLER_0_5_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06944_ _06952_/C _06952_/B _06668_/Y vssd1 vssd1 vccd1 vccd1 _06945_/B sky130_fd_sc_hd__a21o_1
X_06875_ _06877_/B _08951_/B _06876_/A vssd1 vssd1 vccd1 vccd1 _08951_/A sky130_fd_sc_hd__nand3b_1
X_09663_ _09663_/A _09990_/A vssd1 vssd1 vccd1 vccd1 _09665_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05734__A input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05826_ _05826_/A _05826_/B vssd1 vssd1 vccd1 vccd1 _05832_/B sky130_fd_sc_hd__nand2_1
X_09594_ _09918_/B _09594_/B vssd1 vssd1 vccd1 vccd1 _09596_/A sky130_fd_sc_hd__nand2_1
X_08614_ _09210_/A vssd1 vssd1 vccd1 vccd1 _08615_/B sky130_fd_sc_hd__inv_2
X_08545_ _08545_/A _08546_/A vssd1 vssd1 vccd1 vccd1 _08567_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05757_ _05793_/B _05762_/C vssd1 vssd1 vccd1 vccd1 _05761_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05688_ _08574_/A _10187_/A vssd1 vssd1 vccd1 vccd1 _06265_/B sky130_fd_sc_hd__nand2_1
X_08476_ _08476_/A _08476_/B vssd1 vssd1 vccd1 vccd1 _08491_/C sky130_fd_sc_hd__nand2_1
X_07427_ _07427_/A _07427_/B _07427_/C vssd1 vssd1 vccd1 vccd1 _07430_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07358_ _07369_/B _07369_/C vssd1 vssd1 vccd1 vccd1 _07368_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06309_ _06311_/B _06311_/C vssd1 vssd1 vccd1 vccd1 _06310_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07289_ _07289_/A _07289_/B vssd1 vssd1 vccd1 vccd1 _07294_/B sky130_fd_sc_hd__nand2_1
X_09028_ _09028_/A _09028_/B _09028_/C vssd1 vssd1 vccd1 vccd1 _09069_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08004__B _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08020__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05644__A _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08674__B _10188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10705_ _10705_/A _10705_/B vssd1 vssd1 vccd1 vccd1 _10706_/B sky130_fd_sc_hd__nand2_1
X_10636_ _10636_/A hold10/A _10636_/C vssd1 vssd1 vccd1 vccd1 _10637_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06194__B input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10567_ _10694_/A _10593_/C vssd1 vssd1 vccd1 vccd1 _10604_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_51_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05819__A _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10498_ _10504_/A hold46/X _10504_/B vssd1 vssd1 vccd1 vccd1 _10653_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08849__B _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput6 a_i[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_2
XFILLER_0_36_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06660_ _06660_/A _06660_/B vssd1 vssd1 vccd1 vccd1 _06661_/B sky130_fd_sc_hd__nand2_1
X_05611_ _05611_/A _05611_/B vssd1 vssd1 vccd1 vccd1 _05616_/C sky130_fd_sc_hd__nand2_1
X_06591_ _07061_/B _07060_/A _07060_/B vssd1 vssd1 vccd1 vccd1 _07062_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_74_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05542_ _07756_/A _07646_/D vssd1 vssd1 vccd1 vccd1 _05547_/B sky130_fd_sc_hd__nand2_1
X_08330_ _08330_/A _08330_/B _08366_/B vssd1 vssd1 vccd1 vccd1 _08361_/B sky130_fd_sc_hd__nand3_1
X_08261_ _08266_/B _08266_/A vssd1 vssd1 vccd1 vccd1 _08300_/B sky130_fd_sc_hd__nand2_1
X_05473_ _05913_/A _05913_/B vssd1 vssd1 vccd1 vccd1 _05474_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_6_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07212_ _07214_/A _07212_/B vssd1 vssd1 vccd1 vccd1 _07213_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08192_ _08192_/A _08192_/B vssd1 vssd1 vccd1 vccd1 _08193_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06832__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07143_ _07143_/A vssd1 vssd1 vccd1 vccd1 _07146_/A sky130_fd_sc_hd__inv_2
XANTENNA__05729__A _08725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07074_ _07075_/B _07075_/A vssd1 vssd1 vccd1 vccd1 _07074_/Y sky130_fd_sc_hd__nand2_1
X_06025_ _08725_/A _09678_/C vssd1 vssd1 vccd1 vccd1 _06028_/B sky130_fd_sc_hd__nand2_1
X_07976_ _07976_/A _07976_/B vssd1 vssd1 vccd1 vccd1 _08046_/C sky130_fd_sc_hd__nand2_1
X_09715_ _09715_/A _09715_/B vssd1 vssd1 vccd1 vccd1 _09717_/A sky130_fd_sc_hd__xor2_1
X_06927_ _06927_/A _06927_/B vssd1 vssd1 vccd1 vccd1 _09325_/A sky130_fd_sc_hd__nand2_1
X_09646_ _10130_/A _10129_/A _10158_/B _10128_/B vssd1 vssd1 vccd1 vccd1 _09647_/A
+ sky130_fd_sc_hd__and4_1
X_06858_ _06860_/A _10210_/A _08897_/B vssd1 vssd1 vccd1 vccd1 _08935_/A sky130_fd_sc_hd__nand3b_1
X_09577_ _09579_/C vssd1 vssd1 vccd1 vccd1 _09578_/B sky130_fd_sc_hd__inv_2
X_05809_ _05811_/B vssd1 vssd1 vccd1 vccd1 _05810_/B sky130_fd_sc_hd__inv_2
X_06789_ _10156_/A _09677_/A vssd1 vssd1 vccd1 vccd1 _06790_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08528_ _10129_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _08529_/C sky130_fd_sc_hd__nand2_1
X_08459_ _10202_/A _09201_/A _08459_/C vssd1 vssd1 vccd1 vccd1 _08459_/Y sky130_fd_sc_hd__nor3_1
XFILLER_0_9_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10421_ _10681_/A _10418_/Y _10420_/Y vssd1 vssd1 vccd1 vccd1 _10685_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10352_ _10352_/A _10352_/B vssd1 vssd1 vccd1 vccd1 _10357_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05358__B _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10283_ _10286_/B _10286_/C vssd1 vssd1 vccd1 vccd1 _10285_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08685__A _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09455__A2 _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10619_ _10627_/A _10619_/B vssd1 vssd1 vccd1 vccd1 _10632_/A sky130_fd_sc_hd__nor2_1
XANTENNA__05549__A _08672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07830_ _07830_/A _07830_/B vssd1 vssd1 vccd1 vccd1 _08075_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07761_ _09517_/C _08101_/B vssd1 vssd1 vccd1 vccd1 _07763_/A sky130_fd_sc_hd__nand2_1
X_09500_ _09793_/A vssd1 vssd1 vccd1 vccd1 _09501_/B sky130_fd_sc_hd__inv_2
X_06712_ _05932_/B _06710_/Y _06711_/Y vssd1 vssd1 vccd1 vccd1 _06768_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07692_ _07800_/B vssd1 vssd1 vccd1 vccd1 _07692_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_2_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09431_ _09431_/A _09430_/A vssd1 vssd1 vccd1 vccd1 _09432_/B sky130_fd_sc_hd__or2b_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06643_ _06643_/A _06643_/B vssd1 vssd1 vccd1 vccd1 _06969_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06827__B _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06574_ _06685_/B _06596_/C vssd1 vssd1 vccd1 vccd1 _06595_/A sky130_fd_sc_hd__nand2_1
X_09362_ _10112_/A input18/X _10108_/B input19/X vssd1 vssd1 vccd1 vccd1 _09363_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08313_ _09749_/B _10103_/A vssd1 vssd1 vccd1 vccd1 _08314_/A sky130_fd_sc_hd__nand2_1
X_05525_ _05525_/A _05525_/B vssd1 vssd1 vccd1 vccd1 _05527_/A sky130_fd_sc_hd__nand2_1
X_09293_ _09558_/A _09293_/B vssd1 vssd1 vccd1 vccd1 _09294_/B sky130_fd_sc_hd__nand2_1
X_08244_ _08244_/A _08244_/B vssd1 vssd1 vccd1 vccd1 _10467_/A sky130_fd_sc_hd__nor2_1
X_05456_ _05653_/B _05650_/A vssd1 vssd1 vccd1 vccd1 _05457_/B sky130_fd_sc_hd__nand2_2
X_08175_ _08175_/A _08175_/B vssd1 vssd1 vccd1 vccd1 _08177_/A sky130_fd_sc_hd__nand2_1
X_05387_ _05387_/A _05387_/B vssd1 vssd1 vccd1 vccd1 _05634_/B sky130_fd_sc_hd__nand2_1
X_07126_ _07287_/B _07287_/C vssd1 vssd1 vccd1 vccd1 _07289_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07057_ _07057_/A _07065_/A vssd1 vssd1 vccd1 vccd1 _07203_/A sky130_fd_sc_hd__nand2_1
X_06008_ _06008_/A _06008_/B vssd1 vssd1 vccd1 vccd1 _06010_/A sky130_fd_sc_hd__nand2_1
X_07959_ _08060_/B _08059_/B vssd1 vssd1 vccd1 vccd1 _08058_/C sky130_fd_sc_hd__nand2_1
X_09629_ _09629_/A _09629_/B _09629_/C vssd1 vssd1 vccd1 vccd1 _09963_/B sky130_fd_sc_hd__nand3_1
XANTENNA__05641__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10404_ _10404_/A vssd1 vssd1 vccd1 vccd1 _10414_/C sky130_fd_sc_hd__inv_2
XFILLER_0_0_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10335_ _10334_/B _10335_/B _10335_/C vssd1 vssd1 vccd1 vccd1 _10336_/B sky130_fd_sc_hd__nand3b_1
X_10266_ _10266_/A _10266_/B vssd1 vssd1 vccd1 vccd1 _10272_/A sky130_fd_sc_hd__nand2_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08399__B _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10197_ _10199_/B _10198_/B _10198_/A vssd1 vssd1 vccd1 vccd1 _10220_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_17_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05551__B input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06290_ _06425_/A _06424_/A vssd1 vssd1 vccd1 vccd1 _06290_/Y sky130_fd_sc_hd__nor2_1
Xinput31 a_i[8] vssd1 vssd1 vccd1 vccd1 input31/X sky130_fd_sc_hd__clkbuf_1
Xinput20 a_i[27] vssd1 vssd1 vccd1 vccd1 input20/X sky130_fd_sc_hd__buf_2
Xinput53 b_i[28] vssd1 vssd1 vccd1 vccd1 input53/X sky130_fd_sc_hd__buf_2
Xinput42 b_i[18] vssd1 vssd1 vccd1 vccd1 input42/X sky130_fd_sc_hd__buf_1
Xinput64 b_i[9] vssd1 vssd1 vccd1 vccd1 input64/X sky130_fd_sc_hd__buf_4
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09980_ _09980_/A vssd1 vssd1 vccd1 vccd1 _10166_/B sky130_fd_sc_hd__inv_2
X_08931_ _08929_/Y _08858_/B _08930_/Y vssd1 vssd1 vccd1 vccd1 _08937_/A sky130_fd_sc_hd__a21oi_1
X_08862_ _08862_/A _08862_/B vssd1 vssd1 vccd1 vccd1 _08980_/A sky130_fd_sc_hd__nand2_1
X_07813_ _07867_/A _07868_/B vssd1 vssd1 vccd1 vccd1 _07813_/Y sky130_fd_sc_hd__nor2_1
X_08793_ _10210_/A _10275_/B vssd1 vssd1 vccd1 vccd1 _08905_/A sky130_fd_sc_hd__nand2_1
X_07744_ _07744_/A _07744_/B vssd1 vssd1 vccd1 vccd1 _07769_/A sky130_fd_sc_hd__nand2_1
X_07675_ _07675_/A _08574_/A vssd1 vssd1 vccd1 vccd1 _07741_/A sky130_fd_sc_hd__nand2_1
X_09414_ _10156_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _09415_/A sky130_fd_sc_hd__nand2_1
X_06626_ _06968_/B _06968_/C vssd1 vssd1 vccd1 vccd1 _06967_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09345_ _10386_/C vssd1 vssd1 vccd1 vccd1 _10385_/B sky130_fd_sc_hd__inv_2
X_06557_ _06394_/Y _06557_/B _06557_/C vssd1 vssd1 vccd1 vccd1 _06558_/B sky130_fd_sc_hd__nand3b_1
X_09276_ _09278_/B vssd1 vssd1 vccd1 vccd1 _09277_/B sky130_fd_sc_hd__inv_2
X_06488_ _06690_/B _06689_/A vssd1 vssd1 vccd1 vccd1 _06488_/Y sky130_fd_sc_hd__nand2_1
X_05508_ _05510_/B vssd1 vssd1 vccd1 vccd1 _05509_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08227_ _08233_/B _08227_/B vssd1 vssd1 vccd1 vccd1 _08228_/A sky130_fd_sc_hd__nand2_1
X_05439_ _05439_/A _05439_/B vssd1 vssd1 vccd1 vccd1 _05439_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08158_ _10284_/B _10112_/A vssd1 vssd1 vccd1 vccd1 _08162_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08089_ _08089_/A _08382_/B _08089_/C vssd1 vssd1 vccd1 vccd1 _10490_/A sky130_fd_sc_hd__nand3_1
X_07109_ _07267_/A vssd1 vssd1 vccd1 vccd1 _07110_/B sky130_fd_sc_hd__inv_2
XANTENNA_fanout99_A input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10120_ _10120_/A _10120_/B vssd1 vssd1 vccd1 vccd1 _10121_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10051_ _10051_/A _10051_/B vssd1 vssd1 vccd1 vccd1 _10230_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10318_ _10324_/A _10324_/B vssd1 vssd1 vccd1 vccd1 _10323_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10249_ input49/X _10040_/B input50/X _09710_/B vssd1 vssd1 vccd1 vccd1 _10250_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05790_ _05795_/B _06040_/A _05796_/A vssd1 vssd1 vccd1 vccd1 _05794_/A sky130_fd_sc_hd__nand3_1
XANTENNA__07761__B _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06580__A1 _09551_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ _07530_/A _07531_/A vssd1 vssd1 vccd1 vccd1 _07460_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07391_ _09551_/C _09201_/A _07391_/C vssd1 vssd1 vccd1 vccd1 _07392_/A sky130_fd_sc_hd__nor3_1
X_06411_ _06411_/A _06489_/A vssd1 vssd1 vccd1 vccd1 _06679_/C sky130_fd_sc_hd__nand2_1
X_09130_ _09130_/A _09576_/B _09130_/C vssd1 vssd1 vccd1 vccd1 _09576_/A sky130_fd_sc_hd__nand3_1
X_06342_ _06343_/B _06342_/B _06342_/C vssd1 vssd1 vccd1 vccd1 _06652_/B sky130_fd_sc_hd__nand3_1
X_09061_ _09062_/B _09062_/A vssd1 vssd1 vccd1 vccd1 _09061_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_71_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08012_ _08026_/B _08026_/A vssd1 vssd1 vccd1 vccd1 _08142_/C sky130_fd_sc_hd__nand2_1
X_06273_ _08114_/B _09602_/B vssd1 vssd1 vccd1 vccd1 _06438_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_71_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09963_ _09963_/A _09963_/B vssd1 vssd1 vccd1 vccd1 _09966_/A sky130_fd_sc_hd__and2_1
X_08914_ _08914_/A _09111_/A vssd1 vssd1 vccd1 vccd1 _08917_/B sky130_fd_sc_hd__nand2_1
X_09894_ _10306_/A _09900_/B vssd1 vssd1 vccd1 vccd1 _10319_/B sky130_fd_sc_hd__nand2_1
X_08845_ _08930_/A _08846_/A _08846_/B vssd1 vssd1 vccd1 vccd1 _08859_/A sky130_fd_sc_hd__nand3_1
X_08776_ _08806_/B _08776_/B vssd1 vssd1 vccd1 vccd1 _08815_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_79_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05988_ _05990_/A _05990_/B vssd1 vssd1 vccd1 vccd1 _05989_/A sky130_fd_sc_hd__nor2_1
X_07727_ _07727_/A _07727_/B _07727_/C vssd1 vssd1 vccd1 vccd1 _07963_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_67_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08783__A _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07658_ _07666_/B _07667_/C _07667_/B vssd1 vssd1 vccd1 vccd1 _07660_/B sky130_fd_sc_hd__nand3_1
X_07589_ _07857_/B _07597_/B vssd1 vssd1 vccd1 vccd1 _07591_/B sky130_fd_sc_hd__nand2_1
X_06609_ _06957_/B _06609_/B vssd1 vssd1 vccd1 vccd1 _06610_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09328_ _09328_/A _09328_/B _09328_/C vssd1 vssd1 vccd1 vccd1 _09331_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_47_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09259_ _09259_/A _09259_/B vssd1 vssd1 vccd1 vccd1 _09260_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_50_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06750__B _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10103_ _10103_/A _10103_/B input20/X input25/X vssd1 vssd1 vccd1 vccd1 _10105_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__09879__A2 _09551_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10034_ _10259_/A vssd1 vssd1 vccd1 vccd1 _10036_/A sky130_fd_sc_hd__inv_2
XANTENNA__08677__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07756__B _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05557__A _07756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06960_ _06961_/B _06960_/B _06960_/C vssd1 vssd1 vccd1 vccd1 _07127_/B sky130_fd_sc_hd__nand3_1
X_06891_ _06891_/A vssd1 vssd1 vccd1 vccd1 _06892_/B sky130_fd_sc_hd__inv_2
X_05911_ _06734_/B _05911_/B _05911_/C vssd1 vssd1 vccd1 vccd1 _06734_/A sky130_fd_sc_hd__nand3_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08630_ _08630_/A _08630_/B vssd1 vssd1 vccd1 vccd1 _08630_/Y sky130_fd_sc_hd__nor2_1
X_05842_ _05842_/A _05842_/B vssd1 vssd1 vccd1 vccd1 _05887_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08561_ _08879_/B vssd1 vssd1 vccd1 vccd1 _08563_/B sky130_fd_sc_hd__inv_2
X_05773_ _05773_/A _05773_/B vssd1 vssd1 vccd1 vccd1 _05860_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_71_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08492_ _08549_/A _08492_/B _08549_/B vssd1 vssd1 vccd1 vccd1 _08562_/C sky130_fd_sc_hd__nand3_1
X_07512_ _07512_/A _07512_/B _07512_/C vssd1 vssd1 vccd1 vccd1 _07656_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_71_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07443_ _07604_/B _07604_/C vssd1 vssd1 vccd1 vccd1 _07603_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10638__A _10638_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09113_ _09113_/A _09113_/B vssd1 vssd1 vccd1 vccd1 _09119_/B sky130_fd_sc_hd__nand2_1
X_07374_ _07444_/A _07445_/A vssd1 vssd1 vccd1 vccd1 _07435_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_44_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06325_ _06466_/B _06466_/C vssd1 vssd1 vccd1 vccd1 _06465_/A sky130_fd_sc_hd__nand2_1
X_09044_ _09044_/A _09044_/B vssd1 vssd1 vccd1 vccd1 _09044_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06256_ _06256_/A _06256_/B vssd1 vssd1 vccd1 vccd1 _06428_/C sky130_fd_sc_hd__nand2_1
X_06187_ _06189_/B _06189_/C vssd1 vssd1 vccd1 vccd1 _06188_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09946_ _09947_/B _09947_/A vssd1 vssd1 vccd1 vccd1 _09948_/A sky130_fd_sc_hd__or2_1
X_09877_ _10280_/B _09877_/B vssd1 vssd1 vccd1 vccd1 _09877_/Y sky130_fd_sc_hd__nand2_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08828_ _08865_/B _08865_/C vssd1 vssd1 vccd1 vccd1 _08864_/A sky130_fd_sc_hd__nand2_1
X_08759_ _09085_/A vssd1 vssd1 vccd1 vccd1 _08760_/B sky130_fd_sc_hd__inv_2
X_10721_ _10724_/CLK hold27/X fanout99/X vssd1 vssd1 vccd1 vccd1 hold63/A sky130_fd_sc_hd__dfrtp_2
XFILLER_0_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06745__B _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09121__B _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10652_ _10652_/A _10652_/B vssd1 vssd1 vccd1 vccd1 _10654_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10583_ _10595_/A vssd1 vssd1 vccd1 vccd1 _10584_/B sky130_fd_sc_hd__inv_2
XFILLER_0_23_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10017_ _10020_/B _10017_/B _10017_/C vssd1 vssd1 vccd1 vccd1 _10025_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_58_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06110_ _06110_/A _06110_/B vssd1 vssd1 vccd1 vccd1 _06493_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07090_ _07091_/A _07091_/B vssd1 vssd1 vccd1 vccd1 _07228_/A sky130_fd_sc_hd__or2_1
X_06041_ _06041_/A _06041_/B vssd1 vssd1 vccd1 vccd1 _06045_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_10_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06390__B _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09800_ _09800_/A vssd1 vssd1 vccd1 vccd1 _09801_/B sky130_fd_sc_hd__inv_2
X_07992_ _07992_/A _07992_/B vssd1 vssd1 vccd1 vccd1 _08199_/C sky130_fd_sc_hd__nand2_1
X_09731_ _09474_/C _09472_/A _09502_/A vssd1 vssd1 vccd1 vccd1 _09732_/B sky130_fd_sc_hd__o21ai_2
XFILLER_0_5_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06943_ _06943_/A _06943_/B _06943_/C vssd1 vssd1 vccd1 vccd1 _06948_/A sky130_fd_sc_hd__nand3_1
XANTENNA__10717__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06874_ _06874_/A _06874_/B vssd1 vssd1 vccd1 vccd1 _06876_/A sky130_fd_sc_hd__nand2_1
X_09662_ _09664_/A _09663_/A _09990_/A vssd1 vssd1 vccd1 vccd1 _09998_/B sky130_fd_sc_hd__nand3_2
X_05825_ _05821_/Y _05823_/Y _05847_/A vssd1 vssd1 vccd1 vccd1 _05826_/B sky130_fd_sc_hd__a21oi_1
X_09593_ _10158_/A _10156_/B _10157_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _09594_/B
+ sky130_fd_sc_hd__a22o_1
X_08613_ _08513_/B _08516_/B _08511_/A vssd1 vssd1 vccd1 vccd1 _09210_/A sky130_fd_sc_hd__a21oi_2
X_08544_ _08544_/A _08544_/B vssd1 vssd1 vccd1 vccd1 _08546_/A sky130_fd_sc_hd__nand2_1
X_05756_ _05756_/A _05756_/B vssd1 vssd1 vccd1 vccd1 _05762_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_49_246 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05687_ input6/X vssd1 vssd1 vccd1 vccd1 _10187_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_37_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08475_ _08476_/B _08476_/A vssd1 vssd1 vccd1 vccd1 _08491_/A sky130_fd_sc_hd__or2_1
XFILLER_0_9_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07426_ _07426_/A _07426_/B vssd1 vssd1 vccd1 vccd1 _07430_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07357_ _07401_/A _07357_/B _07357_/C vssd1 vssd1 vccd1 vccd1 _07369_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_72_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06308_ _06705_/A _06308_/B _06308_/C vssd1 vssd1 vccd1 vccd1 _06311_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_17_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09027_ _09027_/A _09027_/B vssd1 vssd1 vccd1 vccd1 _09069_/A sky130_fd_sc_hd__nand2_1
X_07288_ _07200_/Y _07300_/B _07239_/Y vssd1 vssd1 vccd1 vccd1 _07289_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_32_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06239_ _06418_/C vssd1 vssd1 vccd1 vccd1 _06417_/B sky130_fd_sc_hd__inv_2
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09929_ _10170_/B _09930_/C _09930_/B vssd1 vssd1 vccd1 vccd1 _09935_/A sky130_fd_sc_hd__a21o_1
XANTENNA__08020__B _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05644__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10704_ _10704_/A _10704_/B vssd1 vssd1 vccd1 vccd1 _10706_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10635_ hold4/X vssd1 vssd1 vccd1 vccd1 _10636_/C sky130_fd_sc_hd__inv_2
XFILLER_0_51_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10566_ _10566_/A _10566_/B vssd1 vssd1 vccd1 vccd1 _10593_/C sky130_fd_sc_hd__nor2_1
XANTENNA__05819__B _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10497_ _10497_/A _10497_/B vssd1 vssd1 vccd1 vccd1 _10504_/A sky130_fd_sc_hd__or2_1
Xinput7 a_i[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__buf_1
X_05610_ _05610_/A vssd1 vssd1 vccd1 vccd1 _05616_/A sky130_fd_sc_hd__inv_2
X_06590_ _06590_/A _06590_/B vssd1 vssd1 vccd1 vccd1 _07060_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_52_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05541_ input34/X vssd1 vssd1 vccd1 vccd1 _07646_/D sky130_fd_sc_hd__buf_6
XFILLER_0_19_408 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05472_ _05472_/A vssd1 vssd1 vccd1 vccd1 _05474_/B sky130_fd_sc_hd__inv_2
X_08260_ _08303_/A _08258_/Y _08304_/B vssd1 vssd1 vccd1 vccd1 _08266_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07211_ _07211_/A vssd1 vssd1 vccd1 vccd1 _07214_/A sky130_fd_sc_hd__inv_2
X_08191_ _08249_/C vssd1 vssd1 vccd1 vccd1 _08193_/A sky130_fd_sc_hd__inv_2
XFILLER_0_27_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07142_ _07146_/B _07143_/A vssd1 vssd1 vccd1 vccd1 _07145_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05729__B input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07073_ _07115_/A _07113_/A vssd1 vssd1 vccd1 vccd1 _07073_/Y sky130_fd_sc_hd__nand2_1
X_06024_ _06028_/A vssd1 vssd1 vccd1 vccd1 _06027_/A sky130_fd_sc_hd__inv_2
XFILLER_0_10_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07975_ _07975_/A _07975_/B _07975_/C vssd1 vssd1 vccd1 vccd1 _07976_/B sky130_fd_sc_hd__nand3_1
X_09714_ _09714_/A _09713_/X vssd1 vssd1 vccd1 vccd1 _09715_/B sky130_fd_sc_hd__or2b_1
X_06926_ _06928_/A _06928_/B vssd1 vssd1 vccd1 vccd1 _06927_/A sky130_fd_sc_hd__nand2_1
X_06857_ input48/X vssd1 vssd1 vccd1 vccd1 _10210_/A sky130_fd_sc_hd__buf_4
X_09645_ _10128_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _09651_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07960__A _08061_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05808_ _09517_/D _09477_/C vssd1 vssd1 vccd1 vccd1 _05811_/B sky130_fd_sc_hd__nand2_1
X_09576_ _09576_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09579_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06788_ _06788_/A _06788_/B vssd1 vssd1 vccd1 vccd1 _06792_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_77_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05739_ _05739_/A _05739_/B vssd1 vssd1 vccd1 vccd1 _06122_/C sky130_fd_sc_hd__nand2_1
X_08527_ _10151_/B vssd1 vssd1 vccd1 vccd1 _08529_/B sky130_fd_sc_hd__inv_2
XFILLER_0_77_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08458_ _08681_/B _08460_/C _08460_/B vssd1 vssd1 vccd1 vccd1 _08461_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_9_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07409_ _07409_/A _07409_/B vssd1 vssd1 vccd1 vccd1 _07446_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_18_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08389_ _08453_/A _10148_/A vssd1 vssd1 vccd1 vccd1 _08703_/A sky130_fd_sc_hd__nand2_1
X_10420_ _10681_/B vssd1 vssd1 vccd1 vccd1 _10420_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10351_ _10353_/B vssd1 vssd1 vccd1 vccd1 _10352_/B sky130_fd_sc_hd__inv_2
XFILLER_0_33_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10282_ _10282_/A _10282_/B vssd1 vssd1 vccd1 vccd1 _10286_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08685__B _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10618_ _10618_/A _10618_/B hold20/X vssd1 vssd1 vccd1 vccd1 _10627_/A sky130_fd_sc_hd__or3b_1
XFILLER_0_24_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05549__B _07646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10549_ _10664_/A _10549_/B vssd1 vssd1 vccd1 vccd1 _10550_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07760_ _07782_/B _07764_/C vssd1 vssd1 vccd1 vccd1 _07762_/A sky130_fd_sc_hd__nand2_1
X_06711_ _06711_/A _06711_/B vssd1 vssd1 vccd1 vccd1 _06711_/Y sky130_fd_sc_hd__nor2_1
X_09430_ _09430_/A _09431_/A vssd1 vssd1 vccd1 vccd1 _09432_/A sky130_fd_sc_hd__or2b_1
X_07691_ _07691_/A _07691_/B vssd1 vssd1 vccd1 vccd1 _07800_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_63_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06642_ _06642_/A _06642_/B _06642_/C vssd1 vssd1 vccd1 vccd1 _06643_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_63_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06573_ _06573_/A _06573_/B vssd1 vssd1 vccd1 vccd1 _06596_/C sky130_fd_sc_hd__nand2_1
X_09361_ _10112_/A _10108_/B input18/X input19/X vssd1 vssd1 vccd1 vccd1 _09361_/X
+ sky130_fd_sc_hd__and4_1
X_09292_ _09292_/A _09292_/B _09292_/C vssd1 vssd1 vccd1 vccd1 _09293_/B sky130_fd_sc_hd__nand3_1
X_08312_ _08312_/A _08312_/B _08312_/C vssd1 vssd1 vccd1 vccd1 _08316_/B sky130_fd_sc_hd__nand3_1
X_05524_ _05524_/A _05524_/B vssd1 vssd1 vccd1 vccd1 _05525_/B sky130_fd_sc_hd__nand2_1
X_08243_ _10487_/B _08378_/B vssd1 vssd1 vccd1 vccd1 _08244_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_19_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05455_ _05650_/A _05455_/B _05650_/B vssd1 vssd1 vccd1 vccd1 _05653_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08174_ _08174_/A _08174_/B vssd1 vssd1 vccd1 vccd1 _08175_/B sky130_fd_sc_hd__nand2_1
X_05386_ _05388_/C vssd1 vssd1 vccd1 vccd1 _05387_/B sky130_fd_sc_hd__inv_2
XFILLER_0_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07125_ _07125_/A _07125_/B _07125_/C vssd1 vssd1 vccd1 vccd1 _07287_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_30_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07056_ _07058_/A vssd1 vssd1 vccd1 vccd1 _07065_/A sky130_fd_sc_hd__inv_2
XANTENNA__10732__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06007_ _05604_/B _05603_/A _05623_/B vssd1 vssd1 vccd1 vccd1 _06008_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__07393__A1 _09551_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ _08040_/B _08041_/A _08041_/B vssd1 vssd1 vccd1 vccd1 _08059_/B sky130_fd_sc_hd__a21boi_4
X_06909_ _06910_/B _06910_/A vssd1 vssd1 vccd1 vccd1 _09040_/B sky130_fd_sc_hd__or2_1
X_07889_ _07889_/A _07902_/A _07889_/C vssd1 vssd1 vccd1 vccd1 _07975_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_69_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09628_ _09629_/A _09629_/C _09629_/B vssd1 vssd1 vccd1 vccd1 _09638_/B sky130_fd_sc_hd__a21o_1
X_09559_ _09559_/A _09559_/B vssd1 vssd1 vccd1 vccd1 _09815_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_65_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10275__B _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10403_ _10425_/A _10403_/B vssd1 vssd1 vccd1 vccd1 _10414_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10334_ _10334_/A _10334_/B vssd1 vssd1 vccd1 vccd1 _10336_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10265_ _10265_/A _10265_/B vssd1 vssd1 vccd1 vccd1 _10266_/B sky130_fd_sc_hd__nand2_1
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10196_ _10196_/A _10196_/B vssd1 vssd1 vccd1 vccd1 _10198_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput10 a_i[18] vssd1 vssd1 vccd1 vccd1 input10/X sky130_fd_sc_hd__buf_1
Xinput21 a_i[28] vssd1 vssd1 vccd1 vccd1 input21/X sky130_fd_sc_hd__clkbuf_2
Xinput54 b_i[29] vssd1 vssd1 vccd1 vccd1 input54/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 b_i[19] vssd1 vssd1 vccd1 vccd1 input43/X sky130_fd_sc_hd__buf_1
XFILLER_0_3_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput32 a_i[9] vssd1 vssd1 vccd1 vccd1 input32/X sky130_fd_sc_hd__clkbuf_1
Xinput65 nrst vssd1 vssd1 vccd1 vccd1 input65/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08930_ _08930_/A _08930_/B vssd1 vssd1 vccd1 vccd1 _08930_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_58_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08861_ _08978_/A vssd1 vssd1 vccd1 vccd1 _08862_/B sky130_fd_sc_hd__inv_2
X_07812_ _07967_/B _07811_/Y vssd1 vssd1 vccd1 vccd1 _07872_/B sky130_fd_sc_hd__nor2b_1
X_08792_ _08791_/B _08792_/B vssd1 vssd1 vccd1 vccd1 _08802_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07743_ _07743_/A _07743_/B vssd1 vssd1 vccd1 vccd1 _07744_/A sky130_fd_sc_hd__nand2_1
X_07674_ _07674_/A _07674_/B vssd1 vssd1 vccd1 vccd1 _07689_/A sky130_fd_sc_hd__nand2_1
X_09413_ _09192_/A _09192_/B _09197_/C vssd1 vssd1 vccd1 vccd1 _09424_/B sky130_fd_sc_hd__o21a_1
X_06625_ _06625_/A _06625_/B _06625_/C vssd1 vssd1 vccd1 vccd1 _06968_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_66_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09344_ _09344_/A _10390_/C vssd1 vssd1 vccd1 vccd1 _10386_/C sky130_fd_sc_hd__nand2_1
X_06556_ _06394_/Y _06555_/Y _06393_/A vssd1 vssd1 vccd1 vccd1 _06558_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09275_ _09275_/A _09534_/A vssd1 vssd1 vccd1 vccd1 _09278_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09230__A _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06487_ _06678_/B _06485_/Y _06486_/Y vssd1 vssd1 vccd1 vccd1 _06689_/A sky130_fd_sc_hd__a21oi_2
X_05507_ _07785_/B _09602_/B vssd1 vssd1 vccd1 vccd1 _05510_/B sky130_fd_sc_hd__nand2_1
X_08226_ _08226_/A _08233_/B _08227_/B vssd1 vssd1 vccd1 vccd1 _08373_/A sky130_fd_sc_hd__nand3_2
X_05438_ _05443_/A _05524_/A vssd1 vssd1 vccd1 vccd1 _05583_/B sky130_fd_sc_hd__nand2_1
X_08157_ _10275_/B _10108_/B vssd1 vssd1 vccd1 vccd1 _08162_/A sky130_fd_sc_hd__nand2_1
X_07108_ _07105_/Y _07579_/C _07107_/Y vssd1 vssd1 vccd1 vccd1 _07267_/A sky130_fd_sc_hd__a21oi_2
X_05369_ _05388_/A _05388_/B vssd1 vssd1 vccd1 vccd1 _05387_/A sky130_fd_sc_hd__nand2_1
X_08088_ _08238_/B vssd1 vssd1 vccd1 vccd1 _08089_/C sky130_fd_sc_hd__inv_2
XFILLER_0_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07039_ _07068_/B _07068_/C vssd1 vssd1 vccd1 vccd1 _07067_/A sky130_fd_sc_hd__nand2_1
X_10050_ _10052_/A vssd1 vssd1 vccd1 vccd1 _10051_/B sky130_fd_sc_hd__inv_2
XANTENNA__09778__C _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10189__B1 _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10317_ _10317_/A _10317_/B _10317_/C vssd1 vssd1 vccd1 vccd1 _10324_/B sky130_fd_sc_hd__nand3_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10248_ _10248_/A _10248_/B _10248_/C _10248_/D vssd1 vssd1 vccd1 vccd1 _10250_/A
+ sky130_fd_sc_hd__or4_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10179_ _10181_/A vssd1 vssd1 vccd1 vccd1 _10180_/B sky130_fd_sc_hd__inv_2
XFILLER_0_28_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06580__A2 _10188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06410_ _06409_/B _06489_/B _06410_/C vssd1 vssd1 vccd1 vccd1 _06489_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_227 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07390_ _08897_/B _10150_/A vssd1 vssd1 vccd1 vccd1 _07391_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06341_ _06506_/B _06507_/B vssd1 vssd1 vccd1 vccd1 _06342_/C sky130_fd_sc_hd__nand2_1
X_09060_ _09328_/A _09328_/B vssd1 vssd1 vccd1 vccd1 _09327_/A sky130_fd_sc_hd__nand2_1
X_06272_ _06436_/A _06437_/B vssd1 vssd1 vccd1 vccd1 _06440_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_8_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08011_ _08198_/B _08199_/B _08199_/A vssd1 vssd1 vccd1 vccd1 _08026_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_4_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09962_ _09962_/A _10100_/A vssd1 vssd1 vccd1 vccd1 _09966_/B sky130_fd_sc_hd__nand2_1
X_08913_ _08913_/A _09111_/B _08913_/C vssd1 vssd1 vccd1 vccd1 _09111_/A sky130_fd_sc_hd__nand3_1
X_09893_ _09893_/A _09893_/B _09893_/C vssd1 vssd1 vccd1 vccd1 _09900_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08844_ _08790_/B _08789_/C _08783_/Y vssd1 vssd1 vccd1 vccd1 _08846_/A sky130_fd_sc_hd__a21bo_1
X_08775_ _08806_/A vssd1 vssd1 vccd1 vccd1 _08776_/B sky130_fd_sc_hd__inv_2
X_05987_ _10212_/B _10151_/A vssd1 vssd1 vccd1 vccd1 _05990_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05753__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07726_ _07726_/A _07726_/B vssd1 vssd1 vccd1 vccd1 _07963_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10104__B1 _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08783__B _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07657_ _07667_/A vssd1 vssd1 vccd1 vccd1 _07666_/B sky130_fd_sc_hd__inv_2
X_07588_ _07595_/B _07595_/C _07594_/B vssd1 vssd1 vccd1 vccd1 _07597_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06584__A _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06608_ _06609_/B _06608_/B _06608_/C vssd1 vssd1 vccd1 vccd1 _06957_/B sky130_fd_sc_hd__nand3_1
X_09327_ _09327_/A _09327_/B vssd1 vssd1 vccd1 vccd1 _09331_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06539_ _09517_/C input35/X vssd1 vssd1 vccd1 vccd1 _07044_/C sky130_fd_sc_hd__nand2_1
X_09258_ _09259_/B _09259_/A vssd1 vssd1 vccd1 vccd1 _09260_/A sky130_fd_sc_hd__or2_1
X_09189_ _09189_/A vssd1 vssd1 vccd1 vccd1 _09194_/B sky130_fd_sc_hd__inv_2
XFILLER_0_50_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08209_ _08249_/A _08249_/C _08275_/B vssd1 vssd1 vccd1 vccd1 _08277_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10102_ _10102_/A vssd1 vssd1 vccd1 vccd1 _10106_/A sky130_fd_sc_hd__inv_2
X_10033_ _10206_/A _10033_/B vssd1 vssd1 vccd1 vccd1 _10259_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05557__B _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06890_ _06890_/A _06890_/B vssd1 vssd1 vccd1 vccd1 _06892_/A sky130_fd_sc_hd__nor2_1
X_05910_ _05910_/A vssd1 vssd1 vccd1 vccd1 _05911_/B sky130_fd_sc_hd__inv_2
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05841_ _05843_/A vssd1 vssd1 vccd1 vccd1 _05842_/B sky130_fd_sc_hd__inv_2
X_08560_ _08560_/A _08560_/B vssd1 vssd1 vccd1 vccd1 _08879_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05772_ _05773_/A _05773_/B vssd1 vssd1 vccd1 vccd1 _05860_/A sky130_fd_sc_hd__or2_1
X_08491_ _08491_/A _08491_/B _08491_/C vssd1 vssd1 vccd1 vccd1 _08549_/B sky130_fd_sc_hd__nand3_1
X_07511_ _07511_/A _07511_/B vssd1 vssd1 vccd1 vccd1 _07656_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_76_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07442_ _07442_/A _07442_/B _07442_/C vssd1 vssd1 vccd1 vccd1 _07604_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07373_ _07348_/Y _07504_/B _07372_/Y vssd1 vssd1 vccd1 vccd1 _07445_/A sky130_fd_sc_hd__a21oi_2
X_09112_ _09114_/C vssd1 vssd1 vccd1 vccd1 _09113_/B sky130_fd_sc_hd__inv_2
XFILLER_0_17_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06324_ _06324_/A _06324_/B _06324_/C vssd1 vssd1 vccd1 vccd1 _06466_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09043_ _09044_/B _09044_/A vssd1 vssd1 vccd1 vccd1 _09071_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_44_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06255_ _06255_/A _06255_/B _06255_/C vssd1 vssd1 vccd1 vccd1 _06256_/B sky130_fd_sc_hd__nand3_1
X_06186_ _06186_/A _06186_/B _06186_/C vssd1 vssd1 vccd1 vccd1 _06189_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_0_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09945_ _09945_/A _09945_/B vssd1 vssd1 vccd1 vccd1 _09947_/A sky130_fd_sc_hd__xor2_1
X_09876_ input52/X _09749_/B input53/X _10275_/B vssd1 vssd1 vccd1 vccd1 _09877_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08827_ _08894_/A _08827_/B _08827_/C vssd1 vssd1 vccd1 vccd1 _08865_/C sky130_fd_sc_hd__nand3_1
XANTENNA__08794__A _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08758_ _08756_/Y _08465_/B _08757_/Y vssd1 vssd1 vccd1 vccd1 _09085_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08689_ _08691_/B _08689_/B vssd1 vssd1 vccd1 vccd1 _08767_/A sky130_fd_sc_hd__nand2_1
X_07709_ _07823_/B _07822_/B vssd1 vssd1 vccd1 vccd1 _07821_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_67_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10720_ _10724_/CLK _10720_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__06745__C _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10651_ _10651_/A vssd1 vssd1 vccd1 vccd1 _10714_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10582_ _10582_/A _10591_/C vssd1 vssd1 vccd1 vccd1 _10595_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05658__A _08672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_361 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10016_ _10184_/A _10018_/B _10019_/B vssd1 vssd1 vccd1 vccd1 _10017_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_25_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06040_ _06040_/A _06040_/B vssd1 vssd1 vccd1 vccd1 _06041_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05568__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07991_ _07991_/A _07991_/B _07991_/C vssd1 vssd1 vccd1 vccd1 _07992_/B sky130_fd_sc_hd__nand3_1
X_09730_ _09733_/B _09733_/C vssd1 vssd1 vccd1 vccd1 _09732_/A sky130_fd_sc_hd__nand2_1
X_06942_ _07111_/B _07111_/C vssd1 vssd1 vccd1 vccd1 _07267_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06399__A _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06873_ _06873_/A vssd1 vssd1 vccd1 vccd1 _06874_/B sky130_fd_sc_hd__inv_2
X_09661_ _09660_/B _09661_/B _09990_/B vssd1 vssd1 vccd1 vccd1 _09990_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05824_ _05824_/A _05824_/B vssd1 vssd1 vccd1 vccd1 _05847_/A sky130_fd_sc_hd__nor2_1
X_09592_ _09592_/A vssd1 vssd1 vccd1 vccd1 _09918_/B sky130_fd_sc_hd__inv_2
X_08612_ _08616_/A _08616_/B vssd1 vssd1 vccd1 vccd1 _09210_/B sky130_fd_sc_hd__nand2_1
X_08543_ _08542_/B _08543_/B _08543_/C vssd1 vssd1 vccd1 vccd1 _08544_/B sky130_fd_sc_hd__nand3b_1
X_05755_ _05755_/A _05755_/B vssd1 vssd1 vccd1 vccd1 _05793_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05686_ _08573_/A _09602_/B vssd1 vssd1 vccd1 vccd1 _06264_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08474_ _08474_/A _08474_/B vssd1 vssd1 vccd1 vccd1 _08476_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07425_ _07427_/A vssd1 vssd1 vccd1 vccd1 _07426_/B sky130_fd_sc_hd__inv_2
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06862__A _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07356_ _07401_/B _07356_/B vssd1 vssd1 vccd1 vccd1 _07369_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_72_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07287_ _07287_/A _07287_/B _07287_/C vssd1 vssd1 vccd1 vccd1 _07294_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_17_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06307_ _06298_/Y _06497_/B _06304_/Y vssd1 vssd1 vccd1 vccd1 _06705_/A sky130_fd_sc_hd__a21oi_1
X_09026_ _09028_/A _09028_/B vssd1 vssd1 vccd1 vccd1 _09027_/A sky130_fd_sc_hd__nand2_1
X_06238_ _06238_/A _06238_/B vssd1 vssd1 vccd1 vccd1 _06418_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_17_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06169_ _05868_/Y _06168_/Y _05867_/A vssd1 vssd1 vccd1 vccd1 _06171_/A sky130_fd_sc_hd__o21ai_1
X_09928_ _09928_/A vssd1 vssd1 vccd1 vccd1 _09930_/B sky130_fd_sc_hd__inv_2
X_09859_ _09859_/A _09859_/B vssd1 vssd1 vccd1 vccd1 _09861_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08029__A _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10703_ _10703_/A vssd1 vssd1 vccd1 vccd1 _10728_/D sky130_fd_sc_hd__clkbuf_1
X_10634_ _10634_/A vssd1 vssd1 vccd1 vccd1 _10636_/A sky130_fd_sc_hd__inv_2
XFILLER_0_63_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10565_ _10698_/A _10694_/B vssd1 vssd1 vccd1 vccd1 _10566_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10496_ _10496_/A _10496_/B vssd1 vssd1 vccd1 vccd1 _10652_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput8 a_i[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__dlymetal6s2s_1
X_05540_ input32/X vssd1 vssd1 vccd1 vccd1 _07756_/A sky130_fd_sc_hd__buf_6
XANTENNA__10188__B _10188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05471_ _05471_/A _05471_/B vssd1 vssd1 vccd1 vccd1 _05474_/A sky130_fd_sc_hd__nand2_1
X_07210_ _07214_/B _07211_/A vssd1 vssd1 vccd1 vccd1 _07213_/A sky130_fd_sc_hd__nand2_1
X_08190_ _08192_/B _08192_/A vssd1 vssd1 vccd1 vccd1 _08249_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07141_ _07144_/B vssd1 vssd1 vccd1 vccd1 _07146_/B sky130_fd_sc_hd__inv_2
XFILLER_0_54_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07072_ _07122_/C _07122_/B _07071_/Y vssd1 vssd1 vccd1 vccd1 _07113_/A sky130_fd_sc_hd__a21oi_1
X_06023_ _07675_/A _10005_/A vssd1 vssd1 vccd1 vccd1 _06028_/A sky130_fd_sc_hd__nand2_1
X_07974_ _08046_/A _08046_/B vssd1 vssd1 vccd1 vccd1 _08045_/A sky130_fd_sc_hd__nand2_1
X_09713_ input46/X _10210_/B _10211_/A _10040_/B vssd1 vssd1 vccd1 vccd1 _09713_/X
+ sky130_fd_sc_hd__a22o_1
X_06925_ _09324_/A _06925_/B _06925_/C vssd1 vssd1 vccd1 vccd1 _06928_/B sky130_fd_sc_hd__nand3_1
X_06856_ _08935_/B _06856_/B vssd1 vssd1 vccd1 vccd1 _06860_/A sky130_fd_sc_hd__nand2_1
X_09644_ _09375_/B _10101_/A _10128_/B _09373_/Y vssd1 vssd1 vccd1 vccd1 _09655_/B
+ sky130_fd_sc_hd__a31oi_1
XANTENNA__09233__A _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05807_ input42/X vssd1 vssd1 vccd1 vccd1 _09477_/C sky130_fd_sc_hd__buf_4
X_09575_ _09579_/A _09821_/B vssd1 vssd1 vccd1 vccd1 _09578_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06787_ _06787_/A _06787_/B vssd1 vssd1 vccd1 vccd1 _08442_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08526_ _08570_/B _08547_/C vssd1 vssd1 vccd1 vccd1 _08545_/A sky130_fd_sc_hd__nand2_1
X_05738_ _05730_/Y _05738_/B _05738_/C vssd1 vssd1 vccd1 vccd1 _05739_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_77_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08457_ _08457_/A vssd1 vssd1 vccd1 vccd1 _08460_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05669_ _05669_/A _05669_/B vssd1 vssd1 vccd1 vccd1 _06248_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_80_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07408_ _07408_/A _07408_/B vssd1 vssd1 vccd1 vccd1 _07409_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08388_ _10386_/A _10386_/B vssd1 vssd1 vccd1 vccd1 _10385_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07339_ _07343_/A _07343_/C vssd1 vssd1 vccd1 vccd1 _07341_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10350_ _10376_/A _10353_/C vssd1 vssd1 vccd1 vccd1 _10352_/A sky130_fd_sc_hd__nand2_1
X_10281_ _10282_/B _10282_/A vssd1 vssd1 vccd1 vccd1 _10286_/B sky130_fd_sc_hd__or2_1
X_09009_ _09041_/A _09018_/B _09009_/C vssd1 vssd1 vccd1 vccd1 _09018_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_20_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10617_ _10617_/A hold13/X vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__nand2_1
X_10548_ _10548_/A _10548_/B vssd1 vssd1 vccd1 vccd1 _10549_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_11_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10479_ _10479_/A _10479_/B vssd1 vssd1 vccd1 vccd1 _10481_/A sky130_fd_sc_hd__nand2_1
X_06710_ _06711_/B _06711_/A vssd1 vssd1 vccd1 vccd1 _06710_/Y sky130_fd_sc_hd__nand2_1
X_07690_ _07690_/A vssd1 vssd1 vccd1 vccd1 _07691_/B sky130_fd_sc_hd__inv_2
XFILLER_0_78_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06641_ _06641_/A _06641_/B vssd1 vssd1 vccd1 vccd1 _06642_/A sky130_fd_sc_hd__nand2_1
X_09360_ _10115_/A input20/X vssd1 vssd1 vccd1 vccd1 _09365_/B sky130_fd_sc_hd__nand2_1
X_06572_ _06572_/A _06572_/B vssd1 vssd1 vccd1 vccd1 _06573_/A sky130_fd_sc_hd__nand2_1
X_09291_ _09291_/A _09291_/B vssd1 vssd1 vccd1 vccd1 _09558_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08311_ _08311_/A _08341_/A vssd1 vssd1 vccd1 vccd1 _08315_/A sky130_fd_sc_hd__nand2_1
X_05523_ _05526_/B _05526_/C vssd1 vssd1 vccd1 vccd1 _05525_/A sky130_fd_sc_hd__nand2_1
X_08242_ _10497_/A _10490_/A _10490_/B vssd1 vssd1 vccd1 vccd1 _08378_/B sky130_fd_sc_hd__nand3_1
X_05454_ _05454_/A _05454_/B vssd1 vssd1 vccd1 vccd1 _05650_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08173_ _08174_/A _08174_/B vssd1 vssd1 vccd1 vccd1 _08175_/A sky130_fd_sc_hd__or2_1
X_05385_ _05385_/A _05385_/B vssd1 vssd1 vccd1 vccd1 _05388_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07124_ _07124_/A _07124_/B _07124_/C vssd1 vssd1 vccd1 vccd1 _07125_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_42_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07055_ _07215_/C _07215_/B _07054_/Y vssd1 vssd1 vccd1 vccd1 _07058_/A sky130_fd_sc_hd__a21oi_1
X_06006_ _06009_/B _06009_/C vssd1 vssd1 vccd1 vccd1 _06008_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07957_ _07957_/A _07957_/B vssd1 vssd1 vccd1 vccd1 _08041_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07393__A2 _09201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ _06060_/A _06058_/A _06072_/A vssd1 vssd1 vccd1 vccd1 _06910_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_69_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07888_ _07902_/B _07888_/B vssd1 vssd1 vccd1 vccd1 _07975_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06587__A _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06839_ _06839_/A _08772_/A _08830_/A vssd1 vssd1 vccd1 vccd1 _06843_/C sky130_fd_sc_hd__nand3_1
X_09627_ _09363_/B _10115_/A input20/X _09361_/X vssd1 vssd1 vccd1 vccd1 _09629_/B
+ sky130_fd_sc_hd__a31o_1
X_09558_ _09558_/A vssd1 vssd1 vccd1 vccd1 _09559_/B sky130_fd_sc_hd__inv_2
XFILLER_0_77_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08509_ _10103_/B _10157_/B vssd1 vssd1 vccd1 vccd1 _08510_/C sky130_fd_sc_hd__nand2_1
X_09489_ input46/X _10040_/B _10211_/A _09710_/B vssd1 vssd1 vccd1 vccd1 _09490_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08307__A _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10402_ _10426_/A _10426_/C vssd1 vssd1 vccd1 vccd1 _10425_/A sky130_fd_sc_hd__nand2_1
X_10333_ _10335_/B _10335_/C vssd1 vssd1 vccd1 vccd1 _10334_/A sky130_fd_sc_hd__nand2_1
X_10264_ _10267_/B _10267_/C vssd1 vssd1 vccd1 vccd1 _10266_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09138__A _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10195_ _10195_/A _10195_/B vssd1 vssd1 vccd1 vccd1 _10196_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07881__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput22 a_i[29] vssd1 vssd1 vccd1 vccd1 input22/X sky130_fd_sc_hd__clkbuf_2
Xinput11 a_i[19] vssd1 vssd1 vccd1 vccd1 input11/X sky130_fd_sc_hd__clkbuf_1
Xinput55 b_i[2] vssd1 vssd1 vccd1 vccd1 input55/X sky130_fd_sc_hd__buf_2
Xinput44 b_i[1] vssd1 vssd1 vccd1 vccd1 input44/X sky130_fd_sc_hd__buf_1
Xinput33 b_i[0] vssd1 vssd1 vccd1 vccd1 input33/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08860_ _08860_/A _08860_/B vssd1 vssd1 vccd1 vccd1 _08978_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07811_ _07811_/A _07811_/B vssd1 vssd1 vccd1 vccd1 _07811_/Y sky130_fd_sc_hd__nand2_1
X_08791_ _08792_/B _08791_/B vssd1 vssd1 vccd1 vccd1 _08802_/A sky130_fd_sc_hd__nand2b_1
XFILLER_0_74_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07742_ _07742_/A vssd1 vssd1 vccd1 vccd1 _07743_/B sky130_fd_sc_hd__inv_2
X_07673_ _07682_/A _07682_/C vssd1 vssd1 vccd1 vccd1 _07674_/A sky130_fd_sc_hd__nand2_1
X_09412_ _09447_/B _09670_/B vssd1 vssd1 vccd1 vccd1 _09445_/A sky130_fd_sc_hd__nand2_1
X_06624_ _06624_/A _06624_/B vssd1 vssd1 vccd1 vccd1 _06625_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09343_ _09353_/A _09354_/A _09343_/C vssd1 vssd1 vccd1 vccd1 _10390_/C sky130_fd_sc_hd__nand3b_1
X_06555_ _06557_/C vssd1 vssd1 vccd1 vccd1 _06555_/Y sky130_fd_sc_hd__inv_2
X_09274_ _09534_/B _09274_/B _09274_/C vssd1 vssd1 vccd1 vccd1 _09534_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_74_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09230__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06486_ _06676_/A _06675_/A vssd1 vssd1 vccd1 vccd1 _06486_/Y sky130_fd_sc_hd__nor2_1
X_05506_ _05510_/A vssd1 vssd1 vccd1 vccd1 _05509_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08225_ _08225_/A _08225_/B _08225_/C vssd1 vssd1 vccd1 vccd1 _08227_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05437_ _05524_/B _05437_/B _05437_/C vssd1 vssd1 vccd1 vccd1 _05524_/A sky130_fd_sc_hd__nand3_1
X_08156_ _08276_/C _08276_/B vssd1 vssd1 vccd1 vccd1 _08277_/B sky130_fd_sc_hd__nand2_1
X_05368_ _05501_/A _05368_/B _05368_/C vssd1 vssd1 vccd1 vccd1 _05388_/B sky130_fd_sc_hd__nand3_1
X_07107_ _07255_/A _07254_/A vssd1 vssd1 vccd1 vccd1 _07107_/Y sky130_fd_sc_hd__nor2_1
X_08087_ _08087_/A _08087_/B vssd1 vssd1 vccd1 vccd1 _08089_/A sky130_fd_sc_hd__nand2_1
X_07038_ _07075_/B _07038_/B vssd1 vssd1 vccd1 vccd1 _07068_/C sky130_fd_sc_hd__nand2_1
X_08989_ _08989_/A _08989_/B vssd1 vssd1 vccd1 vccd1 _09034_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09778__D _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10189__B2 _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10189__A1 _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10316_ _10316_/A _10316_/B vssd1 vssd1 vccd1 vccd1 _10324_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10247_ input51/X _10247_/B vssd1 vssd1 vccd1 vccd1 _10251_/A sky130_fd_sc_hd__nand2_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10178_ _09994_/A _09995_/A _09995_/B vssd1 vssd1 vccd1 vccd1 _10181_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_69_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06340_ _06508_/C vssd1 vssd1 vccd1 vccd1 _06342_/B sky130_fd_sc_hd__inv_2
XFILLER_0_60_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06271_ _08574_/A _10004_/A vssd1 vssd1 vccd1 vccd1 _06437_/B sky130_fd_sc_hd__nand2_1
X_08010_ _08010_/A _08010_/B _08010_/C vssd1 vssd1 vccd1 vccd1 _08199_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_8_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_75 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09961_ _10100_/B _09961_/B _09961_/C vssd1 vssd1 vccd1 vccd1 _10100_/A sky130_fd_sc_hd__nand3_1
X_08912_ _08912_/A _08920_/A vssd1 vssd1 vccd1 vccd1 _08914_/A sky130_fd_sc_hd__nand2_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09892_ _09892_/A _09892_/B vssd1 vssd1 vccd1 vccd1 _10306_/A sky130_fd_sc_hd__nand2_1
X_08843_ _08847_/B vssd1 vssd1 vccd1 vccd1 _08930_/A sky130_fd_sc_hd__inv_2
XANTENNA__08410__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08774_ _08771_/Y _08835_/B _08773_/Y vssd1 vssd1 vccd1 vccd1 _08806_/A sky130_fd_sc_hd__a21oi_2
X_05986_ _10211_/B _10150_/A vssd1 vssd1 vccd1 vccd1 _05990_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05753__B input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07725_ _07727_/A _07727_/B vssd1 vssd1 vccd1 vccd1 _07726_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10104__A1 _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07656_ _07656_/A _07656_/B _07656_/C vssd1 vssd1 vccd1 vccd1 _07664_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_47_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07587_ _07587_/A _07599_/B _07599_/A vssd1 vssd1 vccd1 vccd1 _10453_/B sky130_fd_sc_hd__nand3_2
XANTENNA__06584__B _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06607_ _06615_/B _06616_/C _06616_/B vssd1 vssd1 vccd1 vccd1 _06609_/B sky130_fd_sc_hd__nand3_1
X_09326_ _09328_/C vssd1 vssd1 vccd1 vccd1 _09327_/B sky130_fd_sc_hd__inv_2
X_06538_ _07043_/B _07042_/A vssd1 vssd1 vccd1 vccd1 _07046_/C sky130_fd_sc_hd__nand2_1
X_09257_ _09257_/A _09257_/B vssd1 vssd1 vccd1 vccd1 _09259_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_62_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08208_ _08208_/A _08208_/B vssd1 vssd1 vccd1 vccd1 _08275_/B sky130_fd_sc_hd__nand2_1
X_06469_ _06468_/B _06469_/B _06469_/C vssd1 vssd1 vccd1 vccd1 _06470_/B sky130_fd_sc_hd__nand3b_1
X_09188_ _10156_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09189_/A sky130_fd_sc_hd__nand2_1
X_08139_ _08139_/A _08139_/B _08139_/C vssd1 vssd1 vccd1 vccd1 _08142_/B sky130_fd_sc_hd__nand3_1
X_10101_ _10101_/A input19/X vssd1 vssd1 vccd1 vccd1 _10102_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05944__A _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10032_ _10032_/A _10032_/B vssd1 vssd1 vccd1 vccd1 _10033_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09416__A _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06775__A _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05840_ _05838_/Y _05743_/B _05839_/Y vssd1 vssd1 vccd1 vccd1 _05843_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_55_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05771_ _09517_/D _10005_/A vssd1 vssd1 vccd1 vccd1 _05773_/B sky130_fd_sc_hd__nand2_1
X_07510_ _07512_/A _07512_/B vssd1 vssd1 vccd1 vccd1 _07511_/A sky130_fd_sc_hd__nand2_1
X_08490_ _08550_/B vssd1 vssd1 vccd1 vccd1 _08492_/B sky130_fd_sc_hd__inv_2
X_07441_ _07834_/B _07441_/B vssd1 vssd1 vccd1 vccd1 _07442_/C sky130_fd_sc_hd__nand2_1
X_07372_ _07500_/A _07502_/B vssd1 vssd1 vccd1 vccd1 _07372_/Y sky130_fd_sc_hd__nor2_1
X_09111_ _09111_/A _09111_/B vssd1 vssd1 vccd1 vccd1 _09114_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06323_ _06323_/A _06323_/B vssd1 vssd1 vccd1 vccd1 _06324_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_44_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09042_ _06887_/A _06888_/C _06896_/A vssd1 vssd1 vccd1 vccd1 _09044_/A sky130_fd_sc_hd__o21a_1
XANTENNA__08405__A _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06254_ _06254_/A _06254_/B vssd1 vssd1 vccd1 vccd1 _06256_/A sky130_fd_sc_hd__nand2_1
X_06185_ _06185_/A _06185_/B vssd1 vssd1 vccd1 vccd1 _06189_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09944_ _10112_/A input20/X vssd1 vssd1 vccd1 vccd1 _09945_/B sky130_fd_sc_hd__nand2_1
X_09875_ _10276_/A _10276_/C _10276_/D _09875_/D vssd1 vssd1 vccd1 vccd1 _10280_/B
+ sky130_fd_sc_hd__or4_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08826_ _08894_/B _08826_/B vssd1 vssd1 vccd1 vccd1 _08865_/B sky130_fd_sc_hd__nand2_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08794__B _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08757_ _08757_/A _08757_/B vssd1 vssd1 vccd1 vccd1 _08757_/Y sky130_fd_sc_hd__nor2_1
X_05969_ _05973_/A vssd1 vssd1 vccd1 vccd1 _05972_/A sky130_fd_sc_hd__inv_2
X_08688_ _08688_/A _08688_/B vssd1 vssd1 vccd1 vccd1 _08689_/B sky130_fd_sc_hd__nand2_1
X_07708_ _07726_/B _07706_/Y _07707_/Y vssd1 vssd1 vccd1 vccd1 _07822_/B sky130_fd_sc_hd__a21oi_2
X_07639_ _07783_/C _07777_/A vssd1 vssd1 vccd1 vccd1 _07699_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10650_ _10650_/A _10653_/A vssd1 vssd1 vccd1 vccd1 _10651_/A sky130_fd_sc_hd__and2_1
X_09309_ _09309_/A _09309_/B _09572_/A vssd1 vssd1 vccd1 vccd1 _09310_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10581_ _10591_/A _10581_/B _10591_/C vssd1 vssd1 vccd1 vccd1 _10582_/A sky130_fd_sc_hd__nand3_1
XANTENNA__05939__A _07785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05658__B _07897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10015_ _10018_/A _10019_/C vssd1 vssd1 vccd1 vccd1 _10017_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05568__B input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07990_ _07990_/A vssd1 vssd1 vccd1 vccd1 _07991_/B sky130_fd_sc_hd__inv_2
X_06941_ _06941_/A _06941_/B _06941_/C vssd1 vssd1 vccd1 vccd1 _07111_/C sky130_fd_sc_hd__nand3_1
X_09660_ _09660_/A _09660_/B vssd1 vssd1 vccd1 vccd1 _09663_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06399__B _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06872_ _08842_/A _06872_/B vssd1 vssd1 vccd1 vccd1 _06874_/A sky130_fd_sc_hd__nand2_1
X_08611_ _08611_/A _08611_/B vssd1 vssd1 vccd1 vccd1 _08616_/B sky130_fd_sc_hd__nand2_1
X_05823_ _05848_/A vssd1 vssd1 vccd1 vccd1 _05823_/Y sky130_fd_sc_hd__inv_2
X_09591_ _10158_/A _10157_/A _10151_/B _10156_/B vssd1 vssd1 vccd1 vccd1 _09592_/A
+ sky130_fd_sc_hd__and4_1
XFILLER_0_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08542_ _08542_/A _08542_/B vssd1 vssd1 vccd1 vccd1 _08544_/A sky130_fd_sc_hd__nand2_1
X_05754_ _05756_/B vssd1 vssd1 vccd1 vccd1 _05755_/B sky130_fd_sc_hd__inv_2
XFILLER_0_49_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08473_ _08473_/A _08473_/B vssd1 vssd1 vccd1 vccd1 _08474_/B sky130_fd_sc_hd__nand2_1
X_07424_ _07422_/Y _07835_/C _07423_/Y vssd1 vssd1 vccd1 vccd1 _07431_/A sky130_fd_sc_hd__a21o_1
X_05685_ _06259_/B _06259_/C vssd1 vssd1 vccd1 vccd1 _06258_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10726__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06862__B _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07355_ _07401_/A vssd1 vssd1 vccd1 vccd1 _07356_/B sky130_fd_sc_hd__inv_2
X_07286_ _07286_/A _07286_/B vssd1 vssd1 vccd1 vccd1 _07863_/A sky130_fd_sc_hd__nand2_1
X_06306_ _06705_/B _06306_/B vssd1 vssd1 vccd1 vccd1 _06311_/B sky130_fd_sc_hd__nand2_1
X_09025_ _09025_/A _09025_/B _09025_/C vssd1 vssd1 vccd1 vccd1 _09028_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_60_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06237_ _06236_/B _06237_/B _06237_/C vssd1 vssd1 vccd1 vccd1 _06238_/B sky130_fd_sc_hd__nand3b_1
X_06168_ _06170_/C vssd1 vssd1 vccd1 vccd1 _06168_/Y sky130_fd_sc_hd__inv_2
X_06099_ _05749_/Y _06110_/B _05890_/Y vssd1 vssd1 vccd1 vccd1 _06921_/A sky130_fd_sc_hd__a21oi_1
X_09927_ _09927_/A _09927_/B vssd1 vssd1 vccd1 vccd1 _09928_/A sky130_fd_sc_hd__xor2_1
X_09858_ _09858_/A vssd1 vssd1 vccd1 vccd1 _09861_/A sky130_fd_sc_hd__inv_2
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09789_ _09789_/A _09789_/B vssd1 vssd1 vccd1 vccd1 _09903_/A sky130_fd_sc_hd__nand2_1
X_08809_ _08808_/B _08809_/B _08809_/C vssd1 vssd1 vccd1 vccd1 _08810_/B sky130_fd_sc_hd__nand3b_1
X_10702_ _10702_/A _10705_/A vssd1 vssd1 vccd1 vccd1 _10703_/A sky130_fd_sc_hd__and2_1
XANTENNA__08029__B _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_3__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10633_ _10633_/A hold4/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10564_ _10693_/B vssd1 vssd1 vccd1 vccd1 _10694_/B sky130_fd_sc_hd__inv_2
XFILLER_0_23_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10495_ hold60/X vssd1 vssd1 vccd1 vccd1 _10496_/B sky130_fd_sc_hd__inv_2
Xinput9 a_i[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__buf_1
XFILLER_0_36_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05470_ _05470_/A _05470_/B _05472_/A vssd1 vssd1 vccd1 vccd1 _05480_/B sky130_fd_sc_hd__nand3_1
X_07140_ _07303_/B _07303_/C vssd1 vssd1 vccd1 vccd1 _07305_/B sky130_fd_sc_hd__nand2_1
X_07071_ _07124_/A _07123_/A vssd1 vssd1 vccd1 vccd1 _07071_/Y sky130_fd_sc_hd__nor2_1
X_06022_ _06890_/A vssd1 vssd1 vccd1 vccd1 _06044_/A sky130_fd_sc_hd__inv_2
XFILLER_0_77_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09712_ input46/X _10211_/A _10210_/B _10040_/B vssd1 vssd1 vccd1 vccd1 _09714_/A
+ sky130_fd_sc_hd__and4_1
X_07973_ _08225_/B _08225_/C vssd1 vssd1 vccd1 vccd1 _08064_/A sky130_fd_sc_hd__nand2_1
X_06924_ _09324_/B _06924_/B vssd1 vssd1 vccd1 vccd1 _06928_/A sky130_fd_sc_hd__nand2_1
X_06855_ _06855_/A _06855_/B vssd1 vssd1 vccd1 vccd1 _06856_/B sky130_fd_sc_hd__nand2_1
X_09643_ _09661_/B _09990_/B vssd1 vssd1 vccd1 vccd1 _09660_/A sky130_fd_sc_hd__nand2_1
X_09574_ _09573_/B _09574_/B _09810_/A vssd1 vssd1 vccd1 vccd1 _09821_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__09233__B _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05806_ _05811_/A vssd1 vssd1 vccd1 vccd1 _05810_/A sky130_fd_sc_hd__inv_2
X_06786_ _06788_/B vssd1 vssd1 vccd1 vccd1 _06787_/B sky130_fd_sc_hd__inv_2
X_08525_ _08525_/A _08525_/B vssd1 vssd1 vccd1 vccd1 _08547_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_26_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05737_ _05737_/A vssd1 vssd1 vccd1 vccd1 _05738_/B sky130_fd_sc_hd__inv_2
X_08456_ _10212_/B _10148_/A vssd1 vssd1 vccd1 vccd1 _08457_/A sky130_fd_sc_hd__nand2_1
X_05668_ _05667_/B _05668_/B _05668_/C vssd1 vssd1 vccd1 vccd1 _05669_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07407_ _07407_/A _07407_/B vssd1 vssd1 vccd1 vccd1 _07408_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08387_ _08387_/A _10466_/A _10401_/A vssd1 vssd1 vccd1 vccd1 _10386_/B sky130_fd_sc_hd__nand3_1
X_05599_ _05604_/A _05966_/A vssd1 vssd1 vccd1 vccd1 _05603_/A sky130_fd_sc_hd__nand2_1
X_07338_ _07353_/A _07353_/B vssd1 vssd1 vccd1 vccd1 _07343_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_33_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07269_ _07269_/A _07269_/B vssd1 vssd1 vccd1 vccd1 _07856_/A sky130_fd_sc_hd__nand2_1
X_10280_ _10280_/A _10280_/B vssd1 vssd1 vccd1 vccd1 _10282_/A sky130_fd_sc_hd__nand2_1
X_09008_ _09008_/A _09041_/A vssd1 vssd1 vccd1 vccd1 _09010_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09688__A2 _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06783__A _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10616_ _10616_/A hold12/X vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10547_ _10664_/B _10667_/A _10667_/B vssd1 vssd1 vccd1 vccd1 _10548_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10478_ _10660_/B _10661_/A _10484_/B vssd1 vssd1 vccd1 vccd1 _10503_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__06023__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10289__A3 _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ _06640_/A _06640_/B _06640_/C vssd1 vssd1 vccd1 vccd1 _06643_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06571_ _06571_/A _06572_/A _06572_/B vssd1 vssd1 vccd1 vccd1 _06685_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09290_ _09292_/C vssd1 vssd1 vccd1 vccd1 _09291_/B sky130_fd_sc_hd__inv_2
XFILLER_0_59_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08310_ _08312_/C vssd1 vssd1 vccd1 vccd1 _08341_/A sky130_fd_sc_hd__inv_2
X_05522_ _05522_/A _05954_/A _06001_/A vssd1 vssd1 vccd1 vccd1 _05526_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_74_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08241_ _08241_/A vssd1 vssd1 vccd1 vccd1 _10497_/A sky130_fd_sc_hd__inv_2
X_05453_ _05651_/B vssd1 vssd1 vccd1 vccd1 _05455_/B sky130_fd_sc_hd__inv_2
XFILLER_0_74_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08172_ _10247_/B _08337_/A vssd1 vssd1 vccd1 vccd1 _08174_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_27_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05384_ _05384_/A _05384_/B _05384_/C vssd1 vssd1 vccd1 vccd1 _05385_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_42_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07123_ _07123_/A _07123_/B vssd1 vssd1 vccd1 vccd1 _07125_/A sky130_fd_sc_hd__nand2_1
X_07054_ _07211_/A _07212_/B vssd1 vssd1 vccd1 vccd1 _07054_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06005_ _06884_/A _06005_/B _06810_/A vssd1 vssd1 vccd1 vccd1 _06009_/C sky130_fd_sc_hd__nand3_1
XANTENNA__09228__B _10188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07956_ _07956_/A _07956_/B vssd1 vssd1 vccd1 vccd1 _07957_/B sky130_fd_sc_hd__nand2_1
X_06907_ _06919_/A _06919_/B vssd1 vssd1 vccd1 vccd1 _06918_/A sky130_fd_sc_hd__nand2_1
X_07887_ _07902_/A vssd1 vssd1 vccd1 vccd1 _07888_/B sky130_fd_sc_hd__inv_2
XANTENNA__06587__B _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10741__RESET_B input65/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06838_ _08830_/B _06838_/B vssd1 vssd1 vccd1 vccd1 _06843_/B sky130_fd_sc_hd__nand2_1
X_09626_ _09626_/A _09626_/B vssd1 vssd1 vccd1 vccd1 _09629_/C sky130_fd_sc_hd__nand2_1
X_09557_ _09557_/A _09557_/B vssd1 vssd1 vccd1 vccd1 _09559_/A sky130_fd_sc_hd__nor2_1
X_06769_ _06769_/A _06769_/B _06769_/C vssd1 vssd1 vccd1 vccd1 _06817_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_77_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09488_ input46/X _10211_/A _10040_/B _09710_/B vssd1 vssd1 vccd1 vccd1 _09488_/X
+ sky130_fd_sc_hd__and4_1
X_08508_ input18/X vssd1 vssd1 vccd1 vccd1 _08510_/B sky130_fd_sc_hd__inv_2
X_08439_ _08757_/B _08439_/B vssd1 vssd1 vccd1 vccd1 _08466_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_80_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08307__B _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10401_ _10401_/A _10466_/A vssd1 vssd1 vccd1 vccd1 _10426_/A sky130_fd_sc_hd__nand2_1
X_10332_ _10331_/B _10332_/B _10332_/C vssd1 vssd1 vccd1 vccd1 _10335_/C sky130_fd_sc_hd__nand3b_1
X_10263_ _10263_/A _10263_/B _10263_/C vssd1 vssd1 vccd1 vccd1 _10267_/C sky130_fd_sc_hd__nand3_1
X_10194_ _10196_/B _10195_/A _10195_/B vssd1 vssd1 vccd1 vccd1 _10198_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_68_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 a_i[1] vssd1 vssd1 vccd1 vccd1 input12/X sky130_fd_sc_hd__clkbuf_4
Xinput45 b_i[20] vssd1 vssd1 vccd1 vccd1 input45/X sky130_fd_sc_hd__buf_1
Xinput34 b_i[10] vssd1 vssd1 vccd1 vccd1 input34/X sky130_fd_sc_hd__buf_1
Xinput23 a_i[2] vssd1 vssd1 vccd1 vccd1 input23/X sky130_fd_sc_hd__clkbuf_1
Xinput56 b_i[30] vssd1 vssd1 vccd1 vccd1 input56/X sky130_fd_sc_hd__buf_1
XFILLER_0_12_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08790_ _08846_/B _08790_/B vssd1 vssd1 vccd1 vccd1 _08791_/B sky130_fd_sc_hd__nand2_1
X_07810_ _07811_/B _07811_/A vssd1 vssd1 vccd1 vccd1 _07967_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_74_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07741_ _07741_/A vssd1 vssd1 vccd1 vccd1 _07743_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07672_ _07672_/A _07672_/B vssd1 vssd1 vccd1 vccd1 _07682_/A sky130_fd_sc_hd__nand2_1
X_09411_ _09410_/B _09411_/B _09620_/A vssd1 vssd1 vccd1 vccd1 _09670_/B sky130_fd_sc_hd__nand3b_2
X_06623_ _06623_/A _06623_/B _06623_/C vssd1 vssd1 vccd1 vccd1 _06968_/B sky130_fd_sc_hd__nand3_1
X_09342_ _09353_/B _09353_/A vssd1 vssd1 vccd1 vccd1 _09344_/A sky130_fd_sc_hd__nand2_1
X_06554_ _07034_/A _07034_/B vssd1 vssd1 vccd1 vccd1 _06560_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05505_ _07891_/B input6/X vssd1 vssd1 vccd1 vccd1 _05510_/A sky130_fd_sc_hd__nand2_1
X_09273_ _09534_/B _09274_/C _09274_/B vssd1 vssd1 vccd1 vccd1 _09275_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_74_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06485_ _06675_/A _06676_/A vssd1 vssd1 vccd1 vccd1 _06485_/Y sky130_fd_sc_hd__nand2_1
X_08224_ _08245_/B _08224_/B vssd1 vssd1 vccd1 vccd1 _08226_/A sky130_fd_sc_hd__nor2_1
X_05436_ _05436_/A vssd1 vssd1 vccd1 vccd1 _05437_/B sky130_fd_sc_hd__inv_2
X_08155_ _08155_/A _08155_/B vssd1 vssd1 vccd1 vccd1 _08276_/C sky130_fd_sc_hd__nand2_1
X_05367_ _05501_/B _05367_/B vssd1 vssd1 vccd1 vccd1 _05388_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05767__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07106_ _07106_/A _07106_/B vssd1 vssd1 vccd1 vccd1 _07579_/C sky130_fd_sc_hd__nand2_2
XFILLER_0_30_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08086_ _10490_/B vssd1 vssd1 vccd1 vccd1 _08086_/Y sky130_fd_sc_hd__inv_2
X_07037_ _07031_/Y _07024_/B _07032_/Y vssd1 vssd1 vccd1 vccd1 _07038_/B sky130_fd_sc_hd__a21o_1
XANTENNA__07982__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08988_ _08988_/A _08988_/B _08988_/C vssd1 vssd1 vccd1 vccd1 _08989_/B sky130_fd_sc_hd__nand3_1
X_07939_ _08046_/B _08045_/B _07938_/Y vssd1 vssd1 vccd1 vccd1 _07944_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_3_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09609_ _09608_/B _09936_/B _09609_/C vssd1 vssd1 vccd1 vccd1 _09936_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_65_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10189__A2 _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10315_ _10317_/C _10317_/B vssd1 vssd1 vccd1 vccd1 _10316_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10246_ _10246_/A vssd1 vssd1 vccd1 vccd1 _10253_/B sky130_fd_sc_hd__inv_2
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10177_ _10181_/B _10181_/C vssd1 vssd1 vccd1 vccd1 _10180_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06270_ _08573_/A _10187_/A vssd1 vssd1 vccd1 vccd1 _06436_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09960_ _10100_/B _09961_/C _09961_/B vssd1 vssd1 vccd1 vccd1 _09962_/A sky130_fd_sc_hd__a21o_1
X_08911_ _08913_/C vssd1 vssd1 vccd1 vccd1 _08920_/A sky130_fd_sc_hd__inv_2
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09891_ _09893_/C vssd1 vssd1 vccd1 vccd1 _09892_/B sky130_fd_sc_hd__inv_2
X_08842_ _08842_/A _08842_/B vssd1 vssd1 vccd1 vccd1 _08847_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08410__B _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08773_ _08833_/A _08832_/A vssd1 vssd1 vccd1 vccd1 _08773_/Y sky130_fd_sc_hd__nor2_1
X_05985_ input37/X vssd1 vssd1 vccd1 vccd1 _10150_/A sky130_fd_sc_hd__clkbuf_8
X_07724_ _07724_/A _07724_/B _07724_/C vssd1 vssd1 vccd1 vccd1 _07727_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09522__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07655_ _07727_/C vssd1 vssd1 vccd1 vccd1 _07726_/B sky130_fd_sc_hd__inv_2
XFILLER_0_79_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06606_ _06625_/C _06625_/B _06449_/Y vssd1 vssd1 vccd1 vccd1 _06615_/B sky130_fd_sc_hd__a21o_1
X_07586_ _07593_/B _07848_/A vssd1 vssd1 vccd1 vccd1 _07599_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09325_ _09325_/A vssd1 vssd1 vccd1 vccd1 _09339_/B sky130_fd_sc_hd__inv_2
X_06537_ _09710_/B _10158_/A vssd1 vssd1 vccd1 vccd1 _07042_/A sky130_fd_sc_hd__nand2_1
X_09256_ _10211_/B _09477_/C vssd1 vssd1 vccd1 vccd1 _09257_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_62_124 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06468_ _06468_/A _06468_/B vssd1 vssd1 vccd1 vccd1 _06470_/A sky130_fd_sc_hd__nand2_1
X_08207_ _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08208_/B sky130_fd_sc_hd__nand2_1
X_05419_ _05676_/C vssd1 vssd1 vccd1 vccd1 _05675_/B sky130_fd_sc_hd__inv_2
X_09187_ _09221_/B _09449_/B vssd1 vssd1 vccd1 vccd1 _09220_/A sky130_fd_sc_hd__nand2_1
X_06399_ _08897_/B _10005_/A vssd1 vssd1 vccd1 vccd1 _06400_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08138_ _08138_/A _08199_/A vssd1 vssd1 vccd1 vccd1 _08139_/A sky130_fd_sc_hd__nand2_1
X_08069_ _08069_/A _08069_/B vssd1 vssd1 vccd1 vccd1 _08072_/A sky130_fd_sc_hd__nor2_1
X_10100_ _10100_/A _10100_/B vssd1 vssd1 vccd1 vccd1 _10140_/B sky130_fd_sc_hd__nand2_1
X_10031_ _10212_/B _10201_/B vssd1 vssd1 vccd1 vccd1 _10032_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09416__B _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05944__B _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07217__A _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06775__B _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09151__B _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10229_ _10229_/A _10229_/B vssd1 vssd1 vccd1 vccd1 _10231_/A sky130_fd_sc_hd__nor2_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06031__A _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05770_ input40/X vssd1 vssd1 vccd1 vccd1 _10005_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07440_ _07835_/C vssd1 vssd1 vccd1 vccd1 _07834_/B sky130_fd_sc_hd__inv_2
X_07371_ _07505_/C vssd1 vssd1 vccd1 vccd1 _07504_/B sky130_fd_sc_hd__inv_2
X_09110_ _09544_/B _09114_/B vssd1 vssd1 vccd1 vccd1 _09113_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06322_ _06322_/A _06322_/B vssd1 vssd1 vccd1 vccd1 _06324_/A sky130_fd_sc_hd__nand2_1
X_09041_ _09041_/A _09041_/B vssd1 vssd1 vccd1 vccd1 _09044_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06253_ _06466_/C _06253_/B vssd1 vssd1 vccd1 vccd1 _06254_/B sky130_fd_sc_hd__and2_1
X_06184_ _06186_/C vssd1 vssd1 vccd1 vccd1 _06185_/B sky130_fd_sc_hd__inv_2
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09517__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09943_ _10108_/B input21/X vssd1 vssd1 vccd1 vccd1 _09945_/A sky130_fd_sc_hd__nand2_1
X_09874_ _09874_/A vssd1 vssd1 vccd1 vccd1 _09883_/B sky130_fd_sc_hd__inv_2
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _08894_/A vssd1 vssd1 vccd1 vccd1 _08826_/B sky130_fd_sc_hd__inv_2
XANTENNA__09479__B1 _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08756_ _08757_/B _08757_/A vssd1 vssd1 vccd1 vccd1 _08756_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__05780__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05968_ _10157_/A _09677_/A vssd1 vssd1 vccd1 vccd1 _05973_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08687_ _08688_/A _08688_/B vssd1 vssd1 vccd1 vccd1 _08691_/B sky130_fd_sc_hd__or2_1
X_05899_ _05897_/Y _05496_/B _05898_/Y vssd1 vssd1 vccd1 vccd1 _06708_/A sky130_fd_sc_hd__a21oi_2
X_07707_ _07724_/A _07723_/A vssd1 vssd1 vccd1 vccd1 _07707_/Y sky130_fd_sc_hd__nor2_1
X_07638_ _07777_/A _07638_/B _07777_/B vssd1 vssd1 vccd1 vccd1 _07783_/C sky130_fd_sc_hd__nand3_1
X_07569_ _07835_/A _07835_/B _07834_/B vssd1 vssd1 vccd1 vccd1 _07570_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09308_ _09308_/A _09308_/B vssd1 vssd1 vccd1 vccd1 _09310_/A sky130_fd_sc_hd__nand2_1
X_10580_ _10580_/A vssd1 vssd1 vccd1 vccd1 _10581_/B sky130_fd_sc_hd__inv_2
X_09239_ _09469_/A _09469_/B _09470_/A vssd1 vssd1 vccd1 vccd1 _09244_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_63_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10014_ _10018_/B vssd1 vssd1 vccd1 vccd1 _10019_/C sky130_fd_sc_hd__inv_2
XANTENNA__05690__A _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10101__A _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06940_ _06940_/A vssd1 vssd1 vccd1 vccd1 _06941_/C sky130_fd_sc_hd__inv_2
X_06871_ _08842_/A _06873_/A _06872_/B vssd1 vssd1 vccd1 vccd1 _08951_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_66_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05822_ input1/X _10201_/B vssd1 vssd1 vccd1 vccd1 _05848_/A sky130_fd_sc_hd__nand2_1
X_08610_ _08611_/B _08611_/A vssd1 vssd1 vccd1 vccd1 _08616_/A sky130_fd_sc_hd__or2_1
X_09590_ _10156_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _09596_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05753_ _08739_/A input39/X vssd1 vssd1 vccd1 vccd1 _05756_/B sky130_fd_sc_hd__nand2_1
X_08541_ _08556_/B _08541_/B vssd1 vssd1 vccd1 vccd1 _08542_/B sky130_fd_sc_hd__nand2_1
X_05684_ _05684_/A _05684_/B _05684_/C vssd1 vssd1 vccd1 vccd1 _06259_/C sky130_fd_sc_hd__nand3_1
X_08472_ _08473_/A _08473_/B vssd1 vssd1 vccd1 vccd1 _08474_/A sky130_fd_sc_hd__or2_1
X_07423_ _07566_/A _07565_/A vssd1 vssd1 vccd1 vccd1 _07423_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07354_ _07343_/C _07343_/B _07353_/Y vssd1 vssd1 vccd1 vccd1 _07401_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07285_ _07282_/Y _07283_/Y _07284_/Y vssd1 vssd1 vccd1 vccd1 _07286_/B sky130_fd_sc_hd__a21oi_1
X_06305_ _06298_/Y _06497_/B _06304_/Y vssd1 vssd1 vccd1 vccd1 _06306_/B sky130_fd_sc_hd__a21o_1
X_09024_ _09024_/A _09024_/B vssd1 vssd1 vccd1 vccd1 _09028_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06236_ _06236_/A _06236_/B vssd1 vssd1 vccd1 vccd1 _06238_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06167_ _06320_/A _06320_/B vssd1 vssd1 vccd1 vccd1 _06173_/A sky130_fd_sc_hd__nand2_1
X_06098_ _06103_/B _06103_/C vssd1 vssd1 vccd1 vccd1 _06921_/B sky130_fd_sc_hd__nand2_1
X_09926_ _09926_/A _09925_/X vssd1 vssd1 vccd1 vccd1 _09927_/B sky130_fd_sc_hd__or2b_1
X_09857_ _09863_/A _09864_/B vssd1 vssd1 vccd1 vccd1 _09858_/A sky130_fd_sc_hd__nor2_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09788_ _09790_/C vssd1 vssd1 vccd1 vccd1 _09789_/B sky130_fd_sc_hd__inv_2
X_08808_ _08808_/A _08808_/B vssd1 vssd1 vccd1 vccd1 _08810_/A sky130_fd_sc_hd__nand2_1
X_08739_ _08739_/A vssd1 vssd1 vccd1 vccd1 _09842_/D sky130_fd_sc_hd__inv_2
XANTENNA__09710__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10701_ _10701_/A _10701_/B vssd1 vssd1 vccd1 vccd1 _10705_/A sky130_fd_sc_hd__nand2_1
X_10632_ _10632_/A hold10/A _10632_/C vssd1 vssd1 vccd1 vccd1 _10633_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_36_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10563_ _10563_/A _10697_/B vssd1 vssd1 vccd1 vccd1 _10693_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_36_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10494_ _10500_/A _10500_/C vssd1 vssd1 vccd1 vccd1 _10496_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07070_ _07125_/C vssd1 vssd1 vccd1 vccd1 _07122_/B sky130_fd_sc_hd__inv_2
X_06021_ _05794_/B _05797_/A _06020_/Y vssd1 vssd1 vccd1 vccd1 _06890_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_14_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__05595__A _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09711_ _09711_/A vssd1 vssd1 vccd1 vccd1 _09715_/A sky130_fd_sc_hd__inv_2
XFILLER_0_10_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07972_ _07972_/A _08069_/B vssd1 vssd1 vccd1 vccd1 _08225_/C sky130_fd_sc_hd__nand2_1
X_06923_ _09324_/A vssd1 vssd1 vccd1 vccd1 _06924_/B sky130_fd_sc_hd__inv_2
X_06854_ _06855_/A _06855_/B vssd1 vssd1 vccd1 vccd1 _08935_/B sky130_fd_sc_hd__or2_1
X_09642_ _09642_/A _09963_/A _09642_/C vssd1 vssd1 vccd1 vccd1 _09990_/B sky130_fd_sc_hd__nand3_1
X_09573_ _09573_/A _09573_/B vssd1 vssd1 vccd1 vccd1 _09579_/A sky130_fd_sc_hd__nand2_1
X_05805_ _08112_/A _09698_/A vssd1 vssd1 vccd1 vccd1 _05811_/A sky130_fd_sc_hd__nand2_1
X_06785_ _10158_/A _10187_/A vssd1 vssd1 vccd1 vccd1 _06788_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05736_ _05730_/Y _05732_/Y _05737_/A vssd1 vssd1 vccd1 vccd1 _05739_/A sky130_fd_sc_hd__o21ai_1
X_08524_ _08549_/A _08492_/B _08549_/B vssd1 vssd1 vccd1 vccd1 _08525_/B sky130_fd_sc_hd__a21boi_1
X_08455_ _10202_/A _09201_/A _08459_/C vssd1 vssd1 vccd1 vccd1 _08460_/C sky130_fd_sc_hd__o21ai_1
X_05667_ _05667_/A _05667_/B vssd1 vssd1 vccd1 vccd1 _05669_/A sky130_fd_sc_hd__nand2_1
X_05598_ _05966_/B _05598_/B _05598_/C vssd1 vssd1 vccd1 vccd1 _05966_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_9_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07406_ _07408_/B _07407_/B _07407_/A vssd1 vssd1 vccd1 vccd1 _07409_/A sky130_fd_sc_hd__nand3b_1
X_08386_ _10467_/C _10472_/B _08386_/C vssd1 vssd1 vccd1 vccd1 _10401_/A sky130_fd_sc_hd__nor3_1
XANTENNA__07050__A _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07337_ _07337_/A _07337_/B vssd1 vssd1 vccd1 vccd1 _07343_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07268_ _07270_/C vssd1 vssd1 vccd1 vccd1 _07269_/B sky130_fd_sc_hd__inv_2
X_09007_ _09040_/B _09040_/A vssd1 vssd1 vccd1 vccd1 _09041_/A sky130_fd_sc_hd__or2_1
XFILLER_0_60_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07199_ _07172_/Y _07307_/B _07198_/Y vssd1 vssd1 vccd1 vccd1 _07298_/A sky130_fd_sc_hd__a21oi_2
X_06219_ _06379_/B _06376_/B vssd1 vssd1 vccd1 vccd1 _06220_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09909_ _10076_/B vssd1 vssd1 vccd1 vccd1 _10074_/A sky130_fd_sc_hd__inv_2
XANTENNA__09688__A3 _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06783__B _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10615_ _10615_/A _10618_/A vssd1 vssd1 vccd1 vccd1 _10617_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08056__A _08059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10546_ _10663_/B vssd1 vssd1 vccd1 vccd1 _10664_/B sky130_fd_sc_hd__inv_2
XFILLER_0_51_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10477_ _10484_/A _10484_/B vssd1 vssd1 vccd1 vccd1 _10661_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06023__B _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_79 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06570_ _06570_/A _06570_/B _06570_/C vssd1 vssd1 vccd1 vccd1 _06572_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_59_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05521_ _06001_/B _05521_/B vssd1 vssd1 vccd1 vccd1 _05526_/B sky130_fd_sc_hd__nand2_1
X_08240_ _08240_/A _10493_/B vssd1 vssd1 vccd1 vccd1 _08241_/A sky130_fd_sc_hd__nand2_1
X_05452_ _10201_/A _07897_/B vssd1 vssd1 vccd1 vccd1 _05651_/B sky130_fd_sc_hd__nand2_1
X_08171_ _09778_/D _08171_/B vssd1 vssd1 vccd1 vccd1 _08174_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07122_ _07122_/A _07122_/B _07122_/C vssd1 vssd1 vccd1 vccd1 _07287_/B sky130_fd_sc_hd__nand3_1
X_05383_ _05383_/A vssd1 vssd1 vccd1 vccd1 _05384_/B sky130_fd_sc_hd__inv_2
X_07053_ _07213_/C vssd1 vssd1 vccd1 vccd1 _07215_/B sky130_fd_sc_hd__inv_2
X_06004_ _06884_/B _06004_/B vssd1 vssd1 vccd1 vccd1 _06009_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07955_ _07978_/B _08046_/A vssd1 vssd1 vccd1 vccd1 _07957_/A sky130_fd_sc_hd__nand2_1
X_06906_ _09062_/A _09037_/A _06906_/C vssd1 vssd1 vccd1 vccd1 _06919_/B sky130_fd_sc_hd__nand3_1
X_07886_ _07913_/B _07913_/C _07913_/A vssd1 vssd1 vccd1 vccd1 _07902_/A sky130_fd_sc_hd__a21boi_2
X_09625_ _09626_/B _09626_/A vssd1 vssd1 vccd1 vccd1 _09629_/A sky130_fd_sc_hd__or2_1
X_06837_ _08830_/A vssd1 vssd1 vccd1 vccd1 _06838_/B sky130_fd_sc_hd__inv_2
X_09556_ _09800_/A _09562_/B vssd1 vssd1 vccd1 vccd1 _09815_/B sky130_fd_sc_hd__nand2_1
X_06768_ _06768_/A _06768_/B _08552_/A vssd1 vssd1 vccd1 vccd1 _06769_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_77_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09487_ _10210_/A _10247_/B vssd1 vssd1 vccd1 vccd1 _09491_/A sky130_fd_sc_hd__nand2_1
X_08507_ _08521_/B _08601_/B vssd1 vssd1 vccd1 vccd1 _08519_/A sky130_fd_sc_hd__nand2_1
X_06699_ _06699_/A _06700_/A vssd1 vssd1 vccd1 vccd1 _06702_/A sky130_fd_sc_hd__nand2_1
X_05719_ _07756_/A input64/X vssd1 vssd1 vccd1 vccd1 _06159_/B sky130_fd_sc_hd__nand2_1
X_08438_ _08757_/A vssd1 vssd1 vccd1 vccd1 _08439_/B sky130_fd_sc_hd__inv_2
XANTENNA__10710__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08369_ _08366_/B _08369_/B vssd1 vssd1 vccd1 vccd1 _08370_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_33_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10400_ _10687_/B _10400_/B _10400_/C vssd1 vssd1 vccd1 vccd1 _10555_/A sky130_fd_sc_hd__nand3_1
X_10331_ _10331_/A _10331_/B vssd1 vssd1 vccd1 vccd1 _10335_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10262_ _10262_/A _10262_/B vssd1 vssd1 vccd1 vccd1 _10267_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10193_ _10193_/A _10193_/B vssd1 vssd1 vccd1 vccd1 _10195_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput13 a_i[20] vssd1 vssd1 vccd1 vccd1 input13/X sky130_fd_sc_hd__buf_1
Xinput46 b_i[21] vssd1 vssd1 vccd1 vccd1 input46/X sky130_fd_sc_hd__buf_4
Xinput35 b_i[11] vssd1 vssd1 vccd1 vccd1 input35/X sky130_fd_sc_hd__clkbuf_4
Xinput24 a_i[30] vssd1 vssd1 vccd1 vccd1 input24/X sky130_fd_sc_hd__buf_1
XANTENNA__08514__A _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_233 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput57 b_i[31] vssd1 vssd1 vccd1 vccd1 input57/X sky130_fd_sc_hd__clkbuf_1
X_10529_ _10529_/A hold51/X vssd1 vssd1 vccd1 vccd1 _10529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_24_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07740_ _07768_/A _07769_/B vssd1 vssd1 vccd1 vccd1 _07753_/A sky130_fd_sc_hd__nand2_1
X_07671_ _07671_/A vssd1 vssd1 vccd1 vccd1 _07672_/B sky130_fd_sc_hd__inv_2
X_09410_ _09410_/A _09410_/B vssd1 vssd1 vccd1 vccd1 _09447_/B sky130_fd_sc_hd__nand2_1
X_06622_ _06624_/A _06622_/B vssd1 vssd1 vccd1 vccd1 _06623_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09341_ _09354_/A _09343_/C vssd1 vssd1 vccd1 vccd1 _09353_/B sky130_fd_sc_hd__nand2_1
X_06553_ _06553_/A _06553_/B _06553_/C vssd1 vssd1 vccd1 vccd1 _07034_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05504_ _05531_/A _05532_/A vssd1 vssd1 vccd1 vccd1 _05530_/A sky130_fd_sc_hd__nand2_1
X_09272_ _09272_/A vssd1 vssd1 vccd1 vccd1 _09274_/B sky130_fd_sc_hd__inv_2
XFILLER_0_47_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06484_ _06600_/C _06600_/B _06483_/Y vssd1 vssd1 vccd1 vccd1 _06676_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08223_ _08363_/B _08362_/A _08362_/B vssd1 vssd1 vccd1 vccd1 _08376_/B sky130_fd_sc_hd__nand3b_2
X_05435_ _05435_/A _05436_/A vssd1 vssd1 vccd1 vccd1 _05443_/A sky130_fd_sc_hd__nand2_1
X_08154_ _08154_/A _08154_/B vssd1 vssd1 vccd1 vccd1 _08155_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05366_ _05501_/A vssd1 vssd1 vccd1 vccd1 _05367_/B sky130_fd_sc_hd__inv_2
XANTENNA__08424__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05767__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08085_ _08085_/A _08085_/B _08238_/B vssd1 vssd1 vccd1 vccd1 _10490_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_15_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07105_ _07254_/A _07255_/A vssd1 vssd1 vccd1 vccd1 _07105_/Y sky130_fd_sc_hd__nand2_1
X_07036_ _07036_/A _07036_/B vssd1 vssd1 vccd1 vccd1 _07075_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07982__B _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09255__A _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05783__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _08987_/A _08987_/B vssd1 vssd1 vccd1 vccd1 _08989_/A sky130_fd_sc_hd__nand2_1
X_07938_ _07938_/A _07938_/B vssd1 vssd1 vccd1 vccd1 _07938_/Y sky130_fd_sc_hd__nor2_1
Xclkbuf_2_2__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _10733_/CLK sky130_fd_sc_hd__clkbuf_16
X_07869_ _07872_/B vssd1 vssd1 vccd1 vccd1 _07870_/C sky130_fd_sc_hd__inv_2
X_09608_ _09608_/A _09608_/B vssd1 vssd1 vccd1 vccd1 _09610_/A sky130_fd_sc_hd__nand2_1
X_09539_ _09539_/A _09539_/B vssd1 vssd1 vccd1 vccd1 _09539_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_38_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10314_ _10314_/A _10314_/B _10314_/C vssd1 vssd1 vccd1 vccd1 _10317_/B sky130_fd_sc_hd__nand3_1
X_10245_ _10043_/X _10045_/A _10044_/A vssd1 vssd1 vccd1 vccd1 _10246_/A sky130_fd_sc_hd__a21oi_1
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06789__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10176_ _10176_/A _10176_/B _10176_/C vssd1 vssd1 vccd1 vccd1 _10181_/C sky130_fd_sc_hd__nand3_1
XANTENNA__09165__A _09971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08509__A _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ _09890_/A _10331_/B vssd1 vssd1 vccd1 vccd1 _09893_/C sky130_fd_sc_hd__nand2_1
X_08910_ input49/X input50/X _09778_/D input1/X vssd1 vssd1 vccd1 vccd1 _08913_/C
+ sky130_fd_sc_hd__and4_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08841_ _08978_/B _08978_/C vssd1 vssd1 vccd1 vccd1 _08862_/A sky130_fd_sc_hd__nand2_1
X_08772_ _08772_/A _08772_/B vssd1 vssd1 vccd1 vccd1 _08835_/B sky130_fd_sc_hd__nand2_1
X_05984_ _07756_/A vssd1 vssd1 vccd1 vccd1 _10211_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07723_ _07723_/A _07723_/B vssd1 vssd1 vccd1 vccd1 _07727_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09522__B _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07654_ _07654_/A _07710_/A vssd1 vssd1 vccd1 vccd1 _07727_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06605_ _06605_/A _06605_/B _06605_/C vssd1 vssd1 vccd1 vccd1 _06613_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_47_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07585_ _07594_/B _07585_/B vssd1 vssd1 vccd1 vccd1 _07593_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09324_ _09324_/A _09324_/B vssd1 vssd1 vccd1 vccd1 _09339_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_47_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06536_ _07675_/A vssd1 vssd1 vccd1 vccd1 _09710_/B sky130_fd_sc_hd__buf_8
X_09255_ _10210_/B _09698_/A vssd1 vssd1 vccd1 vccd1 _09257_/A sky130_fd_sc_hd__nand2_1
X_06467_ _06469_/B _06469_/C vssd1 vssd1 vccd1 vccd1 _06468_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08206_ _08206_/A vssd1 vssd1 vccd1 vccd1 _08208_/A sky130_fd_sc_hd__inv_2
XFILLER_0_28_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05418_ _05418_/A _05418_/B vssd1 vssd1 vccd1 vccd1 _05676_/C sky130_fd_sc_hd__nand2_1
X_09186_ _09186_/A _09186_/B _09409_/A vssd1 vssd1 vccd1 vccd1 _09449_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06398_ _09678_/C vssd1 vssd1 vccd1 vccd1 _10188_/B sky130_fd_sc_hd__inv_2
X_08137_ _08145_/A vssd1 vssd1 vccd1 vccd1 _08144_/A sky130_fd_sc_hd__inv_2
X_05349_ input44/X vssd1 vssd1 vccd1 vccd1 _08114_/B sky130_fd_sc_hd__buf_6
XFILLER_0_70_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08068_ _08076_/B _08072_/C vssd1 vssd1 vccd1 vccd1 _08079_/B sky130_fd_sc_hd__nand2_1
X_07019_ _09710_/B _10128_/A vssd1 vssd1 vccd1 vccd1 _07185_/C sky130_fd_sc_hd__nand2_1
X_10030_ _10032_/A _10212_/B _10201_/B vssd1 vssd1 vccd1 vccd1 _10206_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__09416__C _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07217__B _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09151__C _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05688__A _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10228_ _10234_/A _10234_/B vssd1 vssd1 vccd1 vccd1 _10233_/A sky130_fd_sc_hd__nand2_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06031__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10159_ _10159_/A _10159_/B vssd1 vssd1 vccd1 vccd1 _10160_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07370_ _07370_/A _07370_/B vssd1 vssd1 vccd1 vccd1 _07505_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06982__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06321_ _06477_/B _06477_/C vssd1 vssd1 vccd1 vccd1 _06476_/A sky130_fd_sc_hd__nand2_1
X_09040_ _09040_/A _09040_/B vssd1 vssd1 vccd1 vccd1 _09041_/B sky130_fd_sc_hd__nand2_1
X_06252_ _06255_/A _06255_/B vssd1 vssd1 vccd1 vccd1 _06254_/A sky130_fd_sc_hd__nand2_1
X_06183_ _06183_/A _06183_/B vssd1 vssd1 vccd1 vccd1 _06377_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09942_ _09942_/A vssd1 vssd1 vccd1 vccd1 _09947_/B sky130_fd_sc_hd__inv_2
XANTENNA__09517__B input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09873_ _09873_/A _09873_/B vssd1 vssd1 vccd1 vccd1 _09874_/A sky130_fd_sc_hd__nand2_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _08821_/Y _08874_/B _08823_/Y vssd1 vssd1 vccd1 vccd1 _08894_/A sky130_fd_sc_hd__a21oi_2
X_08755_ _09288_/A _08761_/C vssd1 vssd1 vccd1 vccd1 _09085_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09479__A1 _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09479__B2 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05780__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ _07723_/A _07724_/A vssd1 vssd1 vccd1 vccd1 _07706_/Y sky130_fd_sc_hd__nand2_1
X_05967_ _07646_/D vssd1 vssd1 vccd1 vccd1 _10157_/A sky130_fd_sc_hd__clkbuf_8
X_08686_ _10211_/B _09678_/C vssd1 vssd1 vccd1 vccd1 _08688_/B sky130_fd_sc_hd__nand2_1
X_05898_ _05898_/A _05898_/B vssd1 vssd1 vccd1 vccd1 _05898_/Y sky130_fd_sc_hd__nor2_1
X_07637_ _07637_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _07777_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07568_ _07834_/A _07835_/C vssd1 vssd1 vccd1 vccd1 _07570_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07988__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09307_ _09581_/C _09583_/B _09581_/B vssd1 vssd1 vccd1 vccd1 _09317_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06519_ _06642_/C _06642_/B _06518_/Y vssd1 vssd1 vccd1 vccd1 _06650_/A sky130_fd_sc_hd__a21oi_1
X_07499_ _07615_/C vssd1 vssd1 vccd1 vccd1 _07612_/B sky130_fd_sc_hd__inv_2
XFILLER_0_63_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09238_ _08650_/A _09237_/Y _08651_/A vssd1 vssd1 vccd1 vccd1 _09470_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09169_ _09169_/A _09169_/B vssd1 vssd1 vccd1 vccd1 _09399_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10013_ _09607_/A _10012_/Y _09606_/A vssd1 vssd1 vccd1 vccd1 _10018_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_58_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06870_ _06870_/A _06870_/B vssd1 vssd1 vccd1 vccd1 _06872_/B sky130_fd_sc_hd__nand2_1
X_05821_ _05824_/A _05824_/B vssd1 vssd1 vccd1 vccd1 _05821_/Y sky130_fd_sc_hd__nand2_1
X_05752_ _05756_/A vssd1 vssd1 vccd1 vccd1 _05755_/A sky130_fd_sc_hd__inv_2
X_08540_ _08543_/B _08543_/C vssd1 vssd1 vccd1 vccd1 _08542_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05683_ _05683_/A _05683_/B vssd1 vssd1 vccd1 vccd1 _05684_/A sky130_fd_sc_hd__nand2_1
X_08471_ _10112_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _08473_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_9_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07422_ _07565_/A _07566_/A vssd1 vssd1 vccd1 vccd1 _07422_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07353_ _07353_/A _07353_/B vssd1 vssd1 vccd1 vccd1 _07353_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_72_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07284_ _07284_/A _07284_/B vssd1 vssd1 vccd1 vccd1 _07284_/Y sky130_fd_sc_hd__nor2_1
X_06304_ _06494_/A _06495_/B vssd1 vssd1 vccd1 vccd1 _06304_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_72_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09023_ _09025_/A vssd1 vssd1 vccd1 vccd1 _09024_/B sky130_fd_sc_hd__inv_2
X_06235_ _06237_/B _06237_/C vssd1 vssd1 vccd1 vccd1 _06236_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06166_ _06166_/A _06166_/B _06166_/C vssd1 vssd1 vccd1 vccd1 _06320_/B sky130_fd_sc_hd__nand3_1
X_06097_ _06104_/C vssd1 vssd1 vccd1 vccd1 _06101_/B sky130_fd_sc_hd__inv_2
XFILLER_0_40_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10735__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09925_ _10151_/A _10150_/B _10150_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _09925_/X
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07048__A _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09856_ _09862_/B _10265_/A vssd1 vssd1 vccd1 vccd1 _09864_/B sky130_fd_sc_hd__nand2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _08827_/B _08807_/B vssd1 vssd1 vccd1 vccd1 _08808_/B sky130_fd_sc_hd__nand2_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09787_ _09888_/B _09787_/B vssd1 vssd1 vccd1 vccd1 _09790_/C sky130_fd_sc_hd__nand2_1
X_06999_ _06999_/A _06999_/B vssd1 vssd1 vccd1 vccd1 _07139_/C sky130_fd_sc_hd__nand2_1
X_08738_ input46/X vssd1 vssd1 vccd1 vccd1 _09268_/A sky130_fd_sc_hd__inv_2
X_08669_ _08568_/A _08868_/A _08868_/B vssd1 vssd1 vccd1 vccd1 _08670_/B sky130_fd_sc_hd__a21boi_1
XANTENNA__09710__B _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08675__A2 _10188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10700_ _10701_/B _10701_/A vssd1 vssd1 vccd1 vccd1 _10702_/A sky130_fd_sc_hd__or2_1
XFILLER_0_48_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08607__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10631_ hold10/X _10634_/A vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__xnor2_1
X_10562_ _10562_/A _10562_/B vssd1 vssd1 vccd1 vccd1 _10563_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06127__A _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10493_ _10504_/B _10493_/B _10493_/C vssd1 vssd1 vccd1 vccd1 _10500_/C sky130_fd_sc_hd__nand3_1
XANTENNA__08342__A _09875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08061__B _08061_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10112__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__B1 _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06020_ _06020_/A _06020_/B vssd1 vssd1 vccd1 vccd1 _06020_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__05595__B _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07971_ _07971_/A _07971_/B vssd1 vssd1 vccd1 vccd1 _08069_/B sky130_fd_sc_hd__nand2_1
X_09710_ _10210_/A _09710_/B vssd1 vssd1 vccd1 vccd1 _09711_/A sky130_fd_sc_hd__nand2_1
X_06922_ _06101_/C _06101_/B _06921_/Y vssd1 vssd1 vccd1 vccd1 _09324_/A sky130_fd_sc_hd__a21oi_2
X_06853_ input46/X _08112_/A vssd1 vssd1 vccd1 vccd1 _06855_/B sky130_fd_sc_hd__nand2_1
X_09641_ _09641_/A _09641_/B vssd1 vssd1 vccd1 vccd1 _09642_/C sky130_fd_sc_hd__nand2_1
X_09572_ _09572_/A _09572_/B vssd1 vssd1 vccd1 vccd1 _09573_/B sky130_fd_sc_hd__and2_1
X_05804_ input43/X vssd1 vssd1 vccd1 vccd1 _09698_/A sky130_fd_sc_hd__buf_4
X_06784_ _06788_/A vssd1 vssd1 vccd1 vccd1 _06787_/A sky130_fd_sc_hd__inv_2
XFILLER_0_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05735_ _08739_/A _10148_/A vssd1 vssd1 vccd1 vccd1 _05737_/A sky130_fd_sc_hd__nand2_1
X_08523_ _08523_/A _08601_/A vssd1 vssd1 vccd1 vccd1 _08525_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08454_ _10202_/A _09201_/A _08459_/C vssd1 vssd1 vccd1 vccd1 _08681_/B sky130_fd_sc_hd__or3_1
X_05666_ _06251_/B _06124_/A vssd1 vssd1 vccd1 vccd1 _05667_/B sky130_fd_sc_hd__nand2_2
X_05597_ _05597_/A vssd1 vssd1 vccd1 vccd1 _05598_/B sky130_fd_sc_hd__inv_2
XFILLER_0_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07405_ _07405_/A _07405_/B _07405_/C vssd1 vssd1 vccd1 vccd1 _07407_/A sky130_fd_sc_hd__nand3_1
X_08385_ _08385_/A _08385_/B vssd1 vssd1 vccd1 vccd1 _10472_/B sky130_fd_sc_hd__xor2_2
XFILLER_0_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07050__B _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ _07353_/B vssd1 vssd1 vccd1 vccd1 _07337_/B sky130_fd_sc_hd__inv_2
XFILLER_0_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09006_ _09006_/A _09006_/B vssd1 vssd1 vccd1 vccd1 _09040_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07267_ _07267_/A _07267_/B vssd1 vssd1 vccd1 vccd1 _07270_/C sky130_fd_sc_hd__nor2_1
X_07198_ _07303_/A _07305_/B vssd1 vssd1 vccd1 vccd1 _07198_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06218_ _06377_/B _06376_/A _06376_/B vssd1 vssd1 vccd1 vccd1 _06379_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06149_ _08724_/A vssd1 vssd1 vccd1 vccd1 _10210_/B sky130_fd_sc_hd__clkbuf_8
X_09908_ _10320_/A _09908_/B vssd1 vssd1 vccd1 vccd1 _10076_/B sky130_fd_sc_hd__nand2_1
X_09839_ _09839_/A _09839_/B vssd1 vssd1 vccd1 vccd1 _09855_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_68_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08337__A _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10614_ hold12/X vssd1 vssd1 vccd1 vccd1 _10618_/A sky130_fd_sc_hd__inv_2
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10545_ _10545_/A _10668_/B vssd1 vssd1 vccd1 vccd1 _10663_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10476_ _10476_/A hold57/X _10476_/C vssd1 vssd1 vccd1 vccd1 _10484_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09631__A _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05520_ _06001_/A vssd1 vssd1 vccd1 vccd1 _05521_/B sky130_fd_sc_hd__inv_2
X_05451_ _08453_/A vssd1 vssd1 vccd1 vccd1 _10201_/A sky130_fd_sc_hd__clkbuf_8
X_08170_ _08181_/B _08180_/A _08180_/B vssd1 vssd1 vccd1 vccd1 _08252_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_27_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07121_ _07123_/B _07124_/B _07124_/C vssd1 vssd1 vccd1 vccd1 _07122_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_27_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05382_ _05382_/A _05383_/A vssd1 vssd1 vccd1 vccd1 _05385_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07052_ _09749_/B _10156_/A vssd1 vssd1 vccd1 vccd1 _07213_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_30_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06003_ _06884_/A vssd1 vssd1 vccd1 vccd1 _06004_/B sky130_fd_sc_hd__inv_2
XFILLER_0_2_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07954_ _08046_/A _08046_/B _08045_/B vssd1 vssd1 vccd1 vccd1 _07978_/B sky130_fd_sc_hd__nand3_1
X_06905_ _09062_/B _06905_/B vssd1 vssd1 vccd1 vccd1 _06919_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07326__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07885_ _07885_/A _07885_/B vssd1 vssd1 vccd1 vccd1 _07913_/A sky130_fd_sc_hd__nand2_1
X_06836_ _05995_/C _05995_/B _05989_/A vssd1 vssd1 vccd1 vccd1 _08830_/A sky130_fd_sc_hd__a21oi_2
X_09624_ _09622_/X _09624_/B vssd1 vssd1 vccd1 vccd1 _09626_/A sky130_fd_sc_hd__nand2b_1
X_09555_ _09555_/A _09555_/B _09555_/C vssd1 vssd1 vccd1 vccd1 _09562_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_77_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06767_ _06767_/A _06767_/B vssd1 vssd1 vccd1 vccd1 _06769_/A sky130_fd_sc_hd__nand2_1
X_09486_ _09486_/A _09486_/B vssd1 vssd1 vccd1 vccd1 _09494_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05718_ _08724_/A _07646_/D vssd1 vssd1 vccd1 vccd1 _06158_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08157__A _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06698_ _07273_/B _07274_/A _07274_/B vssd1 vssd1 vccd1 vccd1 _06700_/A sky130_fd_sc_hd__nand3_1
X_08506_ _08506_/A _08571_/A _08506_/C vssd1 vssd1 vccd1 vccd1 _08601_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08437_ _08434_/Y _08558_/B _08436_/Y vssd1 vssd1 vccd1 vccd1 _08757_/A sky130_fd_sc_hd__a21oi_2
X_05649_ _05654_/B _05695_/B _05695_/A vssd1 vssd1 vccd1 vccd1 _05706_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_65_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08368_ _10511_/B _10511_/A vssd1 vssd1 vccd1 vccd1 _10520_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_18_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07319_ _07319_/A vssd1 vssd1 vccd1 vccd1 _07322_/A sky130_fd_sc_hd__inv_2
X_08299_ _08331_/B _08299_/B vssd1 vssd1 vccd1 vccd1 _08319_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10330_ _10332_/B _10332_/C vssd1 vssd1 vccd1 vccd1 _10331_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06405__A _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10261_ _10263_/B vssd1 vssd1 vccd1 vccd1 _10262_/B sky130_fd_sc_hd__inv_2
XFILLER_0_14_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10192_ _10193_/B _10193_/A vssd1 vssd1 vccd1 vccd1 _10195_/A sky130_fd_sc_hd__or2_1
XANTENNA__06140__A _07756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput36 b_i[12] vssd1 vssd1 vccd1 vccd1 input36/X sky130_fd_sc_hd__clkbuf_4
Xinput25 a_i[31] vssd1 vssd1 vccd1 vccd1 input25/X sky130_fd_sc_hd__buf_1
XFILLER_0_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput14 a_i[21] vssd1 vssd1 vccd1 vccd1 input14/X sky130_fd_sc_hd__clkbuf_1
Xinput47 b_i[22] vssd1 vssd1 vccd1 vccd1 input47/X sky130_fd_sc_hd__clkbuf_1
Xinput58 b_i[3] vssd1 vssd1 vccd1 vccd1 input58/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__08514__B _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10528_ hold51/X _10529_/A vssd1 vssd1 vccd1 vccd1 _10643_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10459_ _10668_/B vssd1 vssd1 vccd1 vccd1 _10459_/Y sky130_fd_sc_hd__inv_2
XANTENNA__06050__A _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07670_ _07670_/A vssd1 vssd1 vccd1 vccd1 _07672_/A sky130_fd_sc_hd__inv_2
XFILLER_0_59_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09361__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06621_ _06621_/A vssd1 vssd1 vccd1 vccd1 _06624_/A sky130_fd_sc_hd__inv_2
X_09340_ _09340_/A _09340_/B _09340_/C vssd1 vssd1 vccd1 vccd1 _09343_/C sky130_fd_sc_hd__nand3_1
X_06552_ _06552_/A _06552_/B vssd1 vssd1 vccd1 vccd1 _07034_/A sky130_fd_sc_hd__nand2_1
X_09271_ _09271_/A _09271_/B vssd1 vssd1 vccd1 vccd1 _09272_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05503_ _05894_/A vssd1 vssd1 vccd1 vccd1 _05532_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08222_ _08245_/B _08222_/B _08225_/A vssd1 vssd1 vccd1 vccd1 _08362_/B sky130_fd_sc_hd__nand3b_2
X_06483_ _06602_/A _06601_/A vssd1 vssd1 vccd1 vccd1 _06483_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_7_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05434_ _07897_/B _09677_/A vssd1 vssd1 vccd1 vccd1 _05436_/A sky130_fd_sc_hd__nand2_1
X_08153_ _08153_/A _08153_/B _08153_/C vssd1 vssd1 vccd1 vccd1 _08245_/B sky130_fd_sc_hd__nand3_4
XFILLER_0_15_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05365_ _05396_/C _05396_/B _05364_/Y vssd1 vssd1 vccd1 vccd1 _05501_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08424__B _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08084_ _08084_/A _08384_/A _08087_/B vssd1 vssd1 vccd1 vccd1 _08085_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_15_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07104_ _07073_/Y _07117_/B _07103_/Y vssd1 vssd1 vccd1 vccd1 _07255_/A sky130_fd_sc_hd__a21oi_2
X_07035_ _07075_/A _07036_/A _07036_/B vssd1 vssd1 vccd1 vccd1 _07068_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06225__A _06228_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09255__B _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _08988_/C vssd1 vssd1 vccd1 vccd1 _08987_/B sky130_fd_sc_hd__inv_2
XANTENNA__05783__B input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07937_ _07937_/A _07937_/B vssd1 vssd1 vccd1 vccd1 _08045_/B sky130_fd_sc_hd__nand2_1
X_07868_ _07871_/B _07868_/B vssd1 vssd1 vccd1 vccd1 _07870_/B sky130_fd_sc_hd__nand2_1
X_09607_ _09607_/A _09607_/B vssd1 vssd1 vccd1 vccd1 _09608_/B sky130_fd_sc_hd__xnor2_1
X_06819_ _09036_/B _09036_/C vssd1 vssd1 vccd1 vccd1 _06823_/A sky130_fd_sc_hd__nand2_1
X_07799_ _07799_/A _07799_/B vssd1 vssd1 vccd1 vccd1 _07801_/A sky130_fd_sc_hd__nand2_1
X_09538_ _09542_/B _09542_/C vssd1 vssd1 vccd1 vccd1 _09541_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10210__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09469_ _09469_/A _09469_/B vssd1 vssd1 vccd1 vccd1 _09470_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_65_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10043__B1 _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10313_ _10313_/A _10313_/B vssd1 vssd1 vccd1 vccd1 _10317_/C sky130_fd_sc_hd__nand2_1
XANTENNA__06135__A _08672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10244_ _10314_/A _10314_/C vssd1 vssd1 vccd1 vccd1 _10313_/A sky130_fd_sc_hd__nand2_1
X_10175_ _10175_/A _10175_/B vssd1 vssd1 vccd1 vccd1 _10181_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06789__B _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08509__B _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _08840_/A _08840_/B _08840_/C vssd1 vssd1 vccd1 vccd1 _08978_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_20_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08771_ _08832_/A _08833_/A vssd1 vssd1 vccd1 vccd1 _08771_/Y sky130_fd_sc_hd__nand2_1
X_05983_ _06810_/B _05998_/C vssd1 vssd1 vccd1 vccd1 _05997_/A sky130_fd_sc_hd__nand2_1
X_07722_ _07724_/A vssd1 vssd1 vccd1 vccd1 _07723_/B sky130_fd_sc_hd__inv_2
X_07653_ _07653_/A _07710_/B _07653_/C vssd1 vssd1 vccd1 vccd1 _07710_/A sky130_fd_sc_hd__nand3_1
X_06604_ _06943_/B _06943_/C vssd1 vssd1 vccd1 vccd1 _06945_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09323_ _10370_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _09357_/B sky130_fd_sc_hd__nand2_1
X_07584_ _07584_/A _07594_/B _07585_/B vssd1 vssd1 vccd1 vccd1 _07599_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_47_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06535_ _08739_/A _07646_/D vssd1 vssd1 vccd1 vccd1 _07043_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_34_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09254_ _09254_/A vssd1 vssd1 vccd1 vccd1 _09259_/B sky130_fd_sc_hd__inv_2
XFILLER_0_47_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06466_ _06466_/A _06466_/B _06466_/C vssd1 vssd1 vccd1 vccd1 _06469_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_62_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09185_ _09185_/A _09185_/B vssd1 vssd1 vccd1 vccd1 _09186_/A sky130_fd_sc_hd__nand2_1
X_08205_ _08206_/A _08207_/A _08207_/B vssd1 vssd1 vccd1 vccd1 _08249_/A sky130_fd_sc_hd__nand3_1
X_05417_ _05417_/A _05417_/B _05417_/C vssd1 vssd1 vccd1 vccd1 _05418_/B sky130_fd_sc_hd__nand3_1
X_06397_ _09778_/D vssd1 vssd1 vccd1 vccd1 _09551_/C sky130_fd_sc_hd__clkinv_4
X_08136_ _08204_/B _08203_/B _08135_/Y vssd1 vssd1 vccd1 vccd1 _08145_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05348_ _05353_/A _05476_/B vssd1 vssd1 vccd1 vccd1 _05352_/B sky130_fd_sc_hd__nand2_1
X_08067_ _08067_/A _08067_/B vssd1 vssd1 vccd1 vccd1 _08072_/C sky130_fd_sc_hd__nand2_1
X_07018_ _07184_/A _07183_/A vssd1 vssd1 vccd1 vccd1 _07023_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09416__D _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _08969_/A _08969_/B vssd1 vssd1 vccd1 vccd1 _08970_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__05688__B _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10227_ _10227_/A _10227_/B _10227_/C vssd1 vssd1 vccd1 vccd1 _10234_/B sky130_fd_sc_hd__nand3_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10115__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
X_10158_ _10158_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _10159_/B sky130_fd_sc_hd__nand2_1
X_10089_ _10089_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10090_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06982__B _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06320_ _06320_/A _06320_/B _06320_/C vssd1 vssd1 vccd1 vccd1 _06477_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06251_ _06251_/A _06251_/B _06251_/C vssd1 vssd1 vccd1 vccd1 _06255_/A sky130_fd_sc_hd__nand3_1
XANTENNA__10007__B1 _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06182_ _10284_/B _09477_/C _08897_/B _09698_/A vssd1 vssd1 vccd1 vccd1 _06183_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09941_ _10115_/A input22/X vssd1 vssd1 vccd1 vccd1 _09942_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09517__C _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09872_ input56/X _10292_/B vssd1 vssd1 vccd1 vccd1 _10274_/A sky130_fd_sc_hd__nand2_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _08872_/C _08871_/A vssd1 vssd1 vccd1 vccd1 _08823_/Y sky130_fd_sc_hd__nor2_1
X_08754_ _08754_/A _08754_/B _08754_/C vssd1 vssd1 vccd1 vccd1 _08761_/C sky130_fd_sc_hd__nand3_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05966_ _05966_/A _05966_/B vssd1 vssd1 vccd1 vccd1 _05979_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09479__A2 _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07705_ _07733_/C _07733_/B _07704_/Y vssd1 vssd1 vccd1 vccd1 _07724_/A sky130_fd_sc_hd__a21oi_4
X_08685_ _10210_/B _10005_/A vssd1 vssd1 vccd1 vccd1 _08688_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05897_ _05898_/B _05898_/A vssd1 vssd1 vccd1 vccd1 _05897_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07636_ _07778_/B vssd1 vssd1 vccd1 vccd1 _07638_/B sky130_fd_sc_hd__inv_2
X_07567_ _07835_/A _07835_/B vssd1 vssd1 vccd1 vccd1 _07834_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07988__B _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09306_ _09308_/A _09309_/B vssd1 vssd1 vccd1 vccd1 _09581_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06518_ _06638_/A _06639_/B vssd1 vssd1 vccd1 vccd1 _06518_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_63_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09237_ _09237_/A vssd1 vssd1 vccd1 vccd1 _09237_/Y sky130_fd_sc_hd__inv_2
X_07498_ _07498_/A _07498_/B vssd1 vssd1 vccd1 vccd1 _07615_/C sky130_fd_sc_hd__nand2_1
X_06449_ _06621_/A _06622_/B vssd1 vssd1 vccd1 vccd1 _06449_/Y sky130_fd_sc_hd__nor2_1
X_09168_ _09169_/B _09169_/A vssd1 vssd1 vccd1 vccd1 _09173_/B sky130_fd_sc_hd__or2_1
XFILLER_0_16_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ input49/X vssd1 vssd1 vccd1 vccd1 _10248_/A sky130_fd_sc_hd__inv_2
X_08119_ _08119_/A _08119_/B vssd1 vssd1 vccd1 vccd1 _08121_/B sky130_fd_sc_hd__nand2_1
X_10012_ _10012_/A vssd1 vssd1 vccd1 vccd1 _10012_/Y sky130_fd_sc_hd__inv_2
XANTENNA__08059__B _08059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_58_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05820_ _08112_/A _09477_/C vssd1 vssd1 vccd1 vccd1 _05824_/B sky130_fd_sc_hd__nand2_1
X_05751_ _09517_/C input40/X vssd1 vssd1 vccd1 vccd1 _05756_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06993__A _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05682_ _05682_/A _05682_/B _05682_/C vssd1 vssd1 vccd1 vccd1 _06259_/B sky130_fd_sc_hd__nand3_1
X_08470_ _08573_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _08473_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07421_ _07413_/Y _07439_/B _07420_/Y vssd1 vssd1 vccd1 vccd1 _07566_/A sky130_fd_sc_hd__a21oi_2
X_07352_ _07357_/B _07357_/C vssd1 vssd1 vccd1 vccd1 _07401_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06303_ _06310_/B _06302_/Y vssd1 vssd1 vccd1 vccd1 _06497_/B sky130_fd_sc_hd__nor2b_1
XANTENNA__05402__A _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07283_ _10410_/C vssd1 vssd1 vccd1 vccd1 _07283_/Y sky130_fd_sc_hd__inv_2
X_09022_ _09053_/B _09053_/C vssd1 vssd1 vccd1 vccd1 _09052_/A sky130_fd_sc_hd__nand2_1
X_06234_ _06234_/A _06234_/B _06234_/C vssd1 vssd1 vccd1 vccd1 _06237_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_60_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06165_ _06165_/A _06165_/B vssd1 vssd1 vccd1 vccd1 _06320_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06096_ _06928_/C _06096_/B vssd1 vssd1 vccd1 vccd1 _06104_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_40_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09924_ _10151_/A _10150_/A _10148_/B _10150_/B vssd1 vssd1 vccd1 vccd1 _09926_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__07048__B _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09855_ _09855_/A _09855_/B _10265_/B vssd1 vssd1 vccd1 vccd1 _10265_/A sky130_fd_sc_hd__nand3_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08806_ _08806_/A _08806_/B vssd1 vssd1 vccd1 vccd1 _08807_/B sky130_fd_sc_hd__or2_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09786_ _09786_/A _09786_/B vssd1 vssd1 vccd1 vccd1 _09787_/B sky130_fd_sc_hd__nand2_1
X_06998_ _06998_/A _06998_/B _06998_/C vssd1 vssd1 vccd1 vccd1 _06999_/B sky130_fd_sc_hd__nand3_1
X_08737_ _08737_/A vssd1 vssd1 vccd1 vccd1 _08745_/B sky130_fd_sc_hd__inv_2
X_05949_ _05493_/C _05493_/B _05948_/Y vssd1 vssd1 vccd1 vccd1 _06804_/A sky130_fd_sc_hd__a21oi_2
X_08668_ _08668_/A _09134_/A vssd1 vssd1 vccd1 vccd1 _08670_/A sky130_fd_sc_hd__nand2_1
X_07619_ _07644_/B _07644_/C vssd1 vssd1 vccd1 vccd1 _07642_/A sky130_fd_sc_hd__nand2_1
X_10630_ _10630_/A _10630_/B _10632_/C vssd1 vssd1 vccd1 vccd1 _10634_/A sky130_fd_sc_hd__nand3_1
XANTENNA__08607__B _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08599_ _08521_/A _08521_/B _08601_/B vssd1 vssd1 vccd1 vccd1 _08600_/B sky130_fd_sc_hd__a21boi_1
XFILLER_0_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10561_ hold54/X vssd1 vssd1 vccd1 vccd1 _10562_/B sky130_fd_sc_hd__inv_2
X_10492_ _10492_/A _10492_/B vssd1 vssd1 vccd1 vccd1 _10500_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06127__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09454__A _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07874__A1 _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07874__B2 _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06053__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07149__A _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07970_ _08058_/C _08058_/B _07961_/Y vssd1 vssd1 vccd1 vccd1 _07972_/A sky130_fd_sc_hd__a21o_1
XANTENNA__10006__C _10188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06921_ _06921_/A _06921_/B vssd1 vssd1 vccd1 vccd1 _06921_/Y sky130_fd_sc_hd__nor2_1
X_06852_ _10211_/A _09778_/D vssd1 vssd1 vccd1 vccd1 _06855_/A sky130_fd_sc_hd__nand2_1
X_09640_ _09640_/A _09641_/B _09641_/A vssd1 vssd1 vccd1 vccd1 _09661_/B sky130_fd_sc_hd__nand3_1
X_09571_ _09574_/B _09810_/A vssd1 vssd1 vccd1 vccd1 _09573_/A sky130_fd_sc_hd__nand2_1
X_06783_ _10157_/A _10004_/A vssd1 vssd1 vccd1 vccd1 _06788_/A sky130_fd_sc_hd__nand2_1
X_05803_ _05836_/A _05836_/B vssd1 vssd1 vccd1 vccd1 _05835_/A sky130_fd_sc_hd__nand2_1
X_08522_ _08522_/A _08523_/A _08601_/A vssd1 vssd1 vccd1 vccd1 _08570_/B sky130_fd_sc_hd__nand3_2
X_05734_ input38/X vssd1 vssd1 vccd1 vccd1 _10148_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_77_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08453_ _08453_/A _10150_/A vssd1 vssd1 vccd1 vccd1 _08459_/C sky130_fd_sc_hd__nand2_1
X_07404_ _07400_/Y _07368_/B _07401_/Y vssd1 vssd1 vccd1 vccd1 _07405_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05665_ _06125_/B _06124_/A _06124_/B vssd1 vssd1 vccd1 vccd1 _06251_/B sky130_fd_sc_hd__nand3b_2
X_05596_ _05596_/A _05597_/A vssd1 vssd1 vccd1 vccd1 _05604_/A sky130_fd_sc_hd__nand2_1
X_08384_ _08384_/A _08384_/B vssd1 vssd1 vccd1 vccd1 _08385_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_18_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07335_ _10103_/A _09677_/A vssd1 vssd1 vccd1 vccd1 _07353_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_60_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07266_ _07270_/A _07274_/C vssd1 vssd1 vccd1 vccd1 _07269_/A sky130_fd_sc_hd__nand2_1
X_09005_ _09005_/A _09005_/B vssd1 vssd1 vccd1 vccd1 _09006_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_26_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06217_ _06217_/A _06217_/B _06217_/C vssd1 vssd1 vccd1 vccd1 _06376_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_41_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07197_ _07308_/C vssd1 vssd1 vccd1 vccd1 _07307_/B sky130_fd_sc_hd__inv_2
X_06148_ _08725_/A _07646_/D vssd1 vssd1 vccd1 vccd1 _06357_/A sky130_fd_sc_hd__nand2_2
X_06079_ _06077_/Y _05626_/B _06078_/Y vssd1 vssd1 vccd1 vccd1 _06082_/A sky130_fd_sc_hd__a21oi_2
X_09907_ _09907_/A _09907_/B _09907_/C vssd1 vssd1 vccd1 vccd1 _09908_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_6_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09838_ _09718_/A _09718_/B _09718_/C vssd1 vssd1 vccd1 vccd1 _09863_/A sky130_fd_sc_hd__a21boi_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09769_ _09775_/A _09775_/B vssd1 vssd1 vccd1 vccd1 _09902_/B sky130_fd_sc_hd__nand2_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07522__A _08725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10613_ hold21/X _10615_/A vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__nor2_1
X_10544_ _10544_/A _10544_/B vssd1 vssd1 vccd1 vccd1 _10545_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10475_ _10475_/A _10475_/B vssd1 vssd1 vccd1 vccd1 _10484_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08528__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08247__B _08363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05450_ input3/X vssd1 vssd1 vccd1 vccd1 _08453_/A sky130_fd_sc_hd__buf_6
XFILLER_0_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05381_ _08101_/B input7/X vssd1 vssd1 vccd1 vccd1 _05383_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07120_ _07003_/Y _07134_/B _07028_/Y vssd1 vssd1 vccd1 vccd1 _07123_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_82_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07051_ _07211_/A _07212_/B vssd1 vssd1 vccd1 vccd1 _07215_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06002_ _06000_/Y _05525_/B _06001_/Y vssd1 vssd1 vccd1 vccd1 _06884_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07953_ _07953_/A _07953_/B vssd1 vssd1 vccd1 vccd1 _08046_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06511__A _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06904_ _09062_/A vssd1 vssd1 vccd1 vccd1 _06905_/B sky130_fd_sc_hd__inv_2
X_07884_ _07884_/A vssd1 vssd1 vccd1 vccd1 _07885_/B sky130_fd_sc_hd__inv_2
X_06835_ _06839_/A _08772_/A vssd1 vssd1 vccd1 vccd1 _08830_/B sky130_fd_sc_hd__nand2_1
X_09623_ _10112_/A input19/X _10108_/B input20/X vssd1 vssd1 vccd1 vccd1 _09624_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09554_ _09786_/B _09554_/B vssd1 vssd1 vccd1 vccd1 _09555_/C sky130_fd_sc_hd__nand2_1
X_06766_ _08881_/B _06766_/B _06766_/C vssd1 vssd1 vccd1 vccd1 _08881_/A sky130_fd_sc_hd__nand3_2
X_09485_ _09485_/A vssd1 vssd1 vccd1 vccd1 _09744_/B sky130_fd_sc_hd__inv_2
XFILLER_0_53_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05717_ _06121_/A _06121_/B vssd1 vssd1 vccd1 vccd1 _06120_/A sky130_fd_sc_hd__nand2_1
X_06697_ _06697_/A _06697_/B vssd1 vssd1 vccd1 vccd1 _07274_/B sky130_fd_sc_hd__nand2_1
X_08505_ _08505_/A _08505_/B vssd1 vssd1 vccd1 vccd1 _08521_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08436_ _08556_/A _08555_/A vssd1 vssd1 vccd1 vccd1 _08436_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08157__B _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05648_ _05648_/A _05648_/B vssd1 vssd1 vccd1 vccd1 _05695_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08367_ _08367_/A _08367_/B vssd1 vssd1 vccd1 vccd1 _10511_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05579_ _05709_/C vssd1 vssd1 vccd1 vccd1 _05580_/B sky130_fd_sc_hd__inv_2
X_07318_ _07322_/B _07319_/A vssd1 vssd1 vccd1 vccd1 _07321_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_276 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08298_ _08299_/B _08331_/B vssd1 vssd1 vccd1 vccd1 _08319_/A sky130_fd_sc_hd__or2_1
XFILLER_0_33_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07249_ _07241_/Y _07291_/B _07248_/Y vssd1 vssd1 vccd1 vccd1 _07427_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10260_ _10048_/C _10048_/B _10259_/Y vssd1 vssd1 vccd1 vccd1 _10263_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__06405__B _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10191_ _10191_/A _10191_/B vssd1 vssd1 vccd1 vccd1 _10193_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__06140__B _07897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput37 b_i[13] vssd1 vssd1 vccd1 vccd1 input37/X sky130_fd_sc_hd__clkbuf_4
Xinput26 a_i[3] vssd1 vssd1 vccd1 vccd1 input26/X sky130_fd_sc_hd__buf_1
Xinput15 a_i[22] vssd1 vssd1 vccd1 vccd1 input15/X sky130_fd_sc_hd__clkbuf_1
Xinput48 b_i[23] vssd1 vssd1 vccd1 vccd1 input48/X sky130_fd_sc_hd__clkbuf_1
Xinput59 b_i[4] vssd1 vssd1 vccd1 vccd1 input59/X sky130_fd_sc_hd__buf_1
X_10527_ _10527_/A vssd1 vssd1 vccd1 vccd1 _10529_/A sky130_fd_sc_hd__inv_2
X_10458_ _10542_/A hold43/X _10542_/B vssd1 vssd1 vccd1 vccd1 _10668_/B sky130_fd_sc_hd__nand3_1
X_10389_ _10389_/A _10389_/B vssd1 vssd1 vccd1 vccd1 _10394_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06620_ _06624_/B _06621_/A vssd1 vssd1 vccd1 vccd1 _06623_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09361__B _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06551_ _06553_/A vssd1 vssd1 vccd1 vccd1 _06552_/B sky130_fd_sc_hd__inv_2
X_09270_ _09270_/A _09269_/Y vssd1 vssd1 vccd1 vccd1 _09271_/B sky130_fd_sc_hd__or2b_1
XFILLER_0_59_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06482_ _06603_/C vssd1 vssd1 vccd1 vccd1 _06600_/B sky130_fd_sc_hd__inv_2
X_05502_ _05500_/Y _05387_/B _05501_/Y vssd1 vssd1 vccd1 vccd1 _05894_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_7_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08221_ _08224_/B _08245_/B vssd1 vssd1 vccd1 vccd1 _08362_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05433_ input4/X vssd1 vssd1 vccd1 vccd1 _09677_/A sky130_fd_sc_hd__buf_6
XFILLER_0_74_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08152_ _08280_/A vssd1 vssd1 vccd1 vccd1 _08153_/C sky130_fd_sc_hd__inv_2
X_05364_ _05392_/A _05393_/B vssd1 vssd1 vccd1 vccd1 _05364_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08083_ _08087_/A _08083_/B vssd1 vssd1 vccd1 vccd1 _08085_/A sky130_fd_sc_hd__nand2_1
X_07103_ _07113_/A _07115_/A vssd1 vssd1 vccd1 vccd1 _07103_/Y sky130_fd_sc_hd__nor2_1
X_07034_ _07034_/A _07034_/B _07034_/C vssd1 vssd1 vccd1 vccd1 _07036_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_30_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08985_ _08985_/A _08985_/B vssd1 vssd1 vccd1 vccd1 _08988_/C sky130_fd_sc_hd__nor2_1
X_07936_ _07975_/A _07975_/B _07936_/C vssd1 vssd1 vccd1 vccd1 _07937_/B sky130_fd_sc_hd__nand3_1
X_07867_ _07867_/A vssd1 vssd1 vccd1 vccd1 _07871_/B sky130_fd_sc_hd__inv_2
X_09606_ _09606_/A _10012_/A vssd1 vssd1 vccd1 vccd1 _09607_/B sky130_fd_sc_hd__nand2_1
X_06818_ _06818_/A _06818_/B _06818_/C vssd1 vssd1 vccd1 vccd1 _09036_/C sky130_fd_sc_hd__nand3_1
X_07798_ _07798_/A _07798_/B vssd1 vssd1 vccd1 vccd1 _07942_/A sky130_fd_sc_hd__nand2_2
X_09537_ _09537_/A _09771_/A _09766_/A vssd1 vssd1 vccd1 vccd1 _09542_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_78_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06749_ _08435_/B _06753_/B vssd1 vssd1 vccd1 vccd1 _06751_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10210__B _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09468_ _09474_/A _09692_/A vssd1 vssd1 vccd1 vccd1 _09472_/A sky130_fd_sc_hd__nand2_1
X_08419_ _08420_/B _08420_/A vssd1 vssd1 vccd1 vccd1 _08421_/A sky130_fd_sc_hd__or2_1
X_09399_ _09399_/A vssd1 vssd1 vccd1 vccd1 _09400_/B sky130_fd_sc_hd__inv_2
XFILLER_0_34_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10043__B2 _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__A1 input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10312_ _10314_/B vssd1 vssd1 vccd1 vccd1 _10313_/B sky130_fd_sc_hd__inv_2
XANTENNA__06135__B _07891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10243_ _10243_/A _10243_/B _10243_/C vssd1 vssd1 vccd1 vccd1 _10314_/C sky130_fd_sc_hd__nand3_1
X_10174_ _10176_/B vssd1 vssd1 vccd1 vccd1 _10175_/B sky130_fd_sc_hd__inv_2
XFILLER_0_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06326__A _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07157__A _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08770_ _08832_/B vssd1 vssd1 vccd1 vccd1 _08833_/A sky130_fd_sc_hd__inv_2
X_05982_ _05982_/A _05982_/B vssd1 vssd1 vccd1 vccd1 _05998_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09372__A _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07721_ _08075_/A _07721_/B _07721_/C vssd1 vssd1 vccd1 vccd1 _08384_/A sky130_fd_sc_hd__nand3b_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07652_ _07652_/A _07809_/A vssd1 vssd1 vccd1 vccd1 _07654_/A sky130_fd_sc_hd__nand2_1
X_07583_ _07583_/A _07583_/B vssd1 vssd1 vccd1 vccd1 _07585_/B sky130_fd_sc_hd__nand2_1
X_06603_ _06603_/A _06603_/B _06603_/C vssd1 vssd1 vccd1 vccd1 _06943_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_75_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10030__B _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09322_ _09322_/A _09322_/B vssd1 vssd1 vccd1 vccd1 _10364_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06534_ _06661_/A _06659_/A vssd1 vssd1 vccd1 vccd1 _06534_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_47_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09253_ _10040_/B _10201_/B vssd1 vssd1 vccd1 vccd1 _09254_/A sky130_fd_sc_hd__nand2_1
X_06465_ _06465_/A _06465_/B vssd1 vssd1 vccd1 vccd1 _06469_/B sky130_fd_sc_hd__nand2_1
X_09184_ _09184_/A _09184_/B vssd1 vssd1 vccd1 vccd1 _09221_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10729__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08204_ _08203_/B _08204_/B _08204_/C vssd1 vssd1 vccd1 vccd1 _08207_/B sky130_fd_sc_hd__nand3b_1
X_06396_ _06401_/B _06401_/A vssd1 vssd1 vccd1 vccd1 _06579_/C sky130_fd_sc_hd__nand2_1
X_05416_ _05416_/A vssd1 vssd1 vccd1 vccd1 _05417_/B sky130_fd_sc_hd__inv_2
X_08135_ _08135_/A _08135_/B vssd1 vssd1 vccd1 vccd1 _08135_/Y sky130_fd_sc_hd__nor2_1
X_05347_ _05476_/A vssd1 vssd1 vccd1 vccd1 _05353_/A sky130_fd_sc_hd__inv_2
XFILLER_0_43_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08066_ _08066_/A _08066_/B _08066_/C vssd1 vssd1 vccd1 vccd1 _08076_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_11_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07017_ _07184_/B vssd1 vssd1 vccd1 vccd1 _07183_/A sky130_fd_sc_hd__inv_2
XFILLER_0_59_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08968_ _09025_/B _09025_/C vssd1 vssd1 vccd1 vccd1 _09024_/A sky130_fd_sc_hd__nand2_1
X_08899_ input50/X _10284_/B vssd1 vssd1 vccd1 vccd1 _09100_/C sky130_fd_sc_hd__nand2_1
X_07919_ _07919_/A _07919_/B vssd1 vssd1 vccd1 vccd1 _07946_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05985__A input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10226_ _10226_/A _10226_/B vssd1 vssd1 vccd1 vccd1 _10234_/A sky130_fd_sc_hd__nand2_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
X_10157_ _10157_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _10159_/A sky130_fd_sc_hd__nand2_1
X_10088_ _10090_/B _10089_/A _10089_/B vssd1 vssd1 vccd1 vccd1 _10334_/B sky130_fd_sc_hd__nand3b_4
XFILLER_0_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06250_ _06250_/A vssd1 vssd1 vccd1 vccd1 _06251_/A sky130_fd_sc_hd__inv_2
XANTENNA__10007__B2 _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10007__A1 _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06181_ _09778_/D vssd1 vssd1 vccd1 vccd1 _10284_/B sky130_fd_sc_hd__buf_6
XFILLER_0_52_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09940_ _09996_/B vssd1 vssd1 vccd1 vccd1 _09994_/A sky130_fd_sc_hd__inv_2
XANTENNA__09517__D _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09871_ _09893_/A _09893_/B vssd1 vssd1 vccd1 vccd1 _09892_/A sky130_fd_sc_hd__nand2_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _08822_/A _08822_/B vssd1 vssd1 vccd1 vccd1 _08874_/B sky130_fd_sc_hd__nand2_1
X_08753_ _08753_/A _08753_/B vssd1 vssd1 vccd1 vccd1 _09288_/A sky130_fd_sc_hd__nand2_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05965_ _06013_/A _06013_/B vssd1 vssd1 vccd1 vccd1 _06012_/A sky130_fd_sc_hd__nand2_1
X_07704_ _07734_/B _07735_/A vssd1 vssd1 vccd1 vccd1 _07704_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08684_ _10040_/B _10187_/B vssd1 vssd1 vccd1 vccd1 _08767_/B sky130_fd_sc_hd__nand2_1
X_05896_ _06821_/A vssd1 vssd1 vccd1 vccd1 _05963_/A sky130_fd_sc_hd__inv_2
XFILLER_0_45_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07635_ _08112_/A _07897_/B vssd1 vssd1 vccd1 vccd1 _07778_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07566_ _07566_/A _07566_/B _07566_/C vssd1 vssd1 vccd1 vccd1 _07835_/B sky130_fd_sc_hd__nand3_1
X_09305_ _09081_/Y _08958_/B _09082_/Y vssd1 vssd1 vccd1 vccd1 _09309_/B sky130_fd_sc_hd__a21oi_1
X_06517_ _06640_/C vssd1 vssd1 vccd1 vccd1 _06642_/B sky130_fd_sc_hd__inv_2
XFILLER_0_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09236_ _09236_/A _09236_/B vssd1 vssd1 vccd1 vccd1 _09469_/B sky130_fd_sc_hd__nand2_1
X_07497_ _07496_/B _07497_/B _07497_/C vssd1 vssd1 vccd1 vccd1 _07498_/B sky130_fd_sc_hd__nand3b_1
X_06448_ _06623_/C vssd1 vssd1 vccd1 vccd1 _06625_/B sky130_fd_sc_hd__inv_2
XFILLER_0_50_108 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09167_ _09400_/A _09166_/Y vssd1 vssd1 vccd1 vccd1 _09169_/A sky130_fd_sc_hd__nor2b_1
XFILLER_0_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06379_ _06379_/A _06379_/B vssd1 vssd1 vccd1 vccd1 _06380_/A sky130_fd_sc_hd__nand2_1
X_09098_ _09539_/A _09539_/B _09103_/C vssd1 vssd1 vccd1 vccd1 _09105_/A sky130_fd_sc_hd__a21o_1
X_08118_ _08118_/A _08118_/B _08118_/C vssd1 vssd1 vccd1 vccd1 _08185_/B sky130_fd_sc_hd__nand3_1
X_08049_ _08148_/A _08148_/B _08049_/C vssd1 vssd1 vccd1 vccd1 _08212_/B sky130_fd_sc_hd__nand3_1
X_10011_ _10184_/A _10019_/B vssd1 vssd1 vccd1 vccd1 _10018_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07525__A _07756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10209_ _10209_/A _10209_/B vssd1 vssd1 vccd1 vccd1 _10216_/C sky130_fd_sc_hd__nand2_1
X_05750_ input27/X vssd1 vssd1 vccd1 vccd1 _09517_/C sky130_fd_sc_hd__buf_12
XFILLER_0_82_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06993__B _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05681_ _05683_/A _05681_/B vssd1 vssd1 vccd1 vccd1 _05682_/B sky130_fd_sc_hd__nand2_1
X_07420_ _07432_/A _07437_/B vssd1 vssd1 vccd1 vccd1 _07420_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07351_ _07351_/A _07351_/B _07351_/C vssd1 vssd1 vccd1 vccd1 _07357_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_72_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06302_ _06302_/A _06302_/B vssd1 vssd1 vccd1 vccd1 _06302_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_17_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07282_ _07284_/B _07284_/A vssd1 vssd1 vccd1 vccd1 _07282_/Y sky130_fd_sc_hd__nand2_1
X_09021_ _09021_/A _09021_/B _09021_/C vssd1 vssd1 vccd1 vccd1 _09053_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_60_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06233_ _06233_/A _06233_/B vssd1 vssd1 vccd1 vccd1 _06237_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06164_ _06166_/A vssd1 vssd1 vccd1 vccd1 _06165_/B sky130_fd_sc_hd__inv_2
XFILLER_0_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06095_ _06095_/A _06095_/B vssd1 vssd1 vccd1 vccd1 _06096_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_13_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09923_ _09923_/A vssd1 vssd1 vccd1 vccd1 _09927_/A sky130_fd_sc_hd__inv_2
X_09854_ _10255_/A _09854_/B _09854_/C vssd1 vssd1 vccd1 vccd1 _10265_/B sky130_fd_sc_hd__nand3_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _08805_/A _08805_/B vssd1 vssd1 vccd1 vccd1 _08827_/B sky130_fd_sc_hd__nand2_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ _09786_/B _09786_/A vssd1 vssd1 vccd1 vccd1 _09888_/B sky130_fd_sc_hd__or2_1
X_06997_ _07008_/A _07008_/B vssd1 vssd1 vccd1 vccd1 _06998_/C sky130_fd_sc_hd__nand2_1
X_08736_ _10210_/A _09517_/D vssd1 vssd1 vccd1 vccd1 _08737_/A sky130_fd_sc_hd__nand2_1
X_05948_ _05948_/A _05948_/B vssd1 vssd1 vccd1 vccd1 _05948_/Y sky130_fd_sc_hd__nor2_1
X_08667_ _08667_/A _08668_/A _09134_/A vssd1 vssd1 vccd1 vccd1 _09133_/B sky130_fd_sc_hd__nand3_2
X_05879_ _06202_/B _06199_/A vssd1 vssd1 vccd1 vccd1 _06188_/B sky130_fd_sc_hd__nand2_1
X_07618_ _07618_/A _07618_/B vssd1 vssd1 vccd1 vccd1 _07644_/B sky130_fd_sc_hd__nand2_1
X_08598_ _08602_/B _09156_/A vssd1 vssd1 vccd1 vccd1 _08600_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08176__A _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07549_ _07664_/C vssd1 vssd1 vccd1 vccd1 _07663_/B sky130_fd_sc_hd__inv_2
XFILLER_0_36_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10560_ _10560_/A _10560_/B vssd1 vssd1 vccd1 vccd1 _10562_/A sky130_fd_sc_hd__nand2_1
X_09219_ _09219_/A _09219_/B vssd1 vssd1 vccd1 vccd1 _09220_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10491_ _10493_/C vssd1 vssd1 vccd1 vccd1 _10492_/B sky130_fd_sc_hd__inv_2
XFILLER_0_63_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09454__B _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07874__A2 _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10689_ _10689_/A vssd1 vssd1 vccd1 vccd1 _10724_/D sky130_fd_sc_hd__clkbuf_1
XANTENNA__06334__A _08672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06053__B _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07149__B _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09645__A _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06920_ _06925_/B _06925_/C vssd1 vssd1 vccd1 vccd1 _09324_/B sky130_fd_sc_hd__nand2_1
X_06851_ _06881_/B _06881_/C vssd1 vssd1 vccd1 vccd1 _06880_/A sky130_fd_sc_hd__nand2_1
X_09570_ _09570_/A _09570_/B _09810_/B vssd1 vssd1 vccd1 vccd1 _09810_/A sky130_fd_sc_hd__nand3_2
X_06782_ _06782_/A _08769_/A vssd1 vssd1 vccd1 vccd1 _06801_/C sky130_fd_sc_hd__nand2_1
X_05802_ _05802_/A _05802_/B vssd1 vssd1 vccd1 vccd1 _05836_/B sky130_fd_sc_hd__nand2_1
X_08521_ _08521_/A _08521_/B _08601_/B vssd1 vssd1 vccd1 vccd1 _08601_/A sky130_fd_sc_hd__nand3_1
X_05733_ input28/X vssd1 vssd1 vccd1 vccd1 _08739_/A sky130_fd_sc_hd__buf_6
XFILLER_0_77_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08452_ input4/X vssd1 vssd1 vccd1 vccd1 _10202_/A sky130_fd_sc_hd__inv_2
X_07403_ _07403_/A _07403_/B vssd1 vssd1 vccd1 vccd1 _07407_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05664_ _05664_/A _05664_/B vssd1 vssd1 vccd1 vccd1 _06124_/B sky130_fd_sc_hd__nand2_1
X_05595_ _10212_/B _10156_/A vssd1 vssd1 vccd1 vccd1 _05597_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08383_ _10472_/C _08383_/B vssd1 vssd1 vccd1 vccd1 _10467_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_18_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06228__B _06228_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08724__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07334_ _07353_/A vssd1 vssd1 vccd1 vccd1 _07337_/A sky130_fd_sc_hd__inv_2
X_07265_ _07265_/A _07265_/B vssd1 vssd1 vccd1 vccd1 _07270_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09004_ _09018_/B _09009_/C vssd1 vssd1 vccd1 vccd1 _09008_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06216_ _06216_/A _06216_/B vssd1 vssd1 vccd1 vccd1 _06376_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_60_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07196_ _07196_/A _07206_/A vssd1 vssd1 vccd1 vccd1 _07308_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_13_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06147_ _06233_/A _06234_/A vssd1 vssd1 vccd1 vccd1 _06147_/Y sky130_fd_sc_hd__nand2_1
X_06078_ _06078_/A _06078_/B vssd1 vssd1 vccd1 vccd1 _06078_/Y sky130_fd_sc_hd__nor2_1
X_09906_ _09906_/A _09906_/B vssd1 vssd1 vccd1 vccd1 _10320_/A sky130_fd_sc_hd__nand2_1
X_09837_ _09837_/A vssd1 vssd1 vccd1 vccd1 _10080_/B sky130_fd_sc_hd__inv_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ _09763_/Y _09768_/B _09768_/C vssd1 vssd1 vccd1 vccd1 _09775_/B sky130_fd_sc_hd__nand3b_1
X_08719_ _10248_/B _10202_/C _08722_/C vssd1 vssd1 vccd1 vccd1 _08781_/C sky130_fd_sc_hd__o21ai_2
X_09699_ _09699_/A _10027_/A _10202_/C _10202_/D vssd1 vssd1 vccd1 vccd1 _10035_/B
+ sky130_fd_sc_hd__or4_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10612_ _10616_/A vssd1 vssd1 vccd1 vccd1 _10615_/A sky130_fd_sc_hd__inv_2
X_10543_ hold43/X vssd1 vssd1 vccd1 vccd1 _10544_/B sky130_fd_sc_hd__inv_2
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10474_ hold57/A vssd1 vssd1 vccd1 vccd1 _10475_/B sky130_fd_sc_hd__inv_2
XFILLER_0_63_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08528__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06329__A _08453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06048__B _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05380_ input60/X vssd1 vssd1 vccd1 vccd1 _08101_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_105 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07050_ _09840_/B _10157_/A vssd1 vssd1 vccd1 vccd1 _07212_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_27_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06064__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06001_ _06001_/A _06001_/B vssd1 vssd1 vccd1 vccd1 _06001_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_2_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07952_ _07952_/A _07952_/B vssd1 vssd1 vccd1 vccd1 _07953_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06511__B _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06903_ _06901_/Y _06088_/B _06902_/Y vssd1 vssd1 vccd1 vccd1 _09062_/A sky130_fd_sc_hd__a21oi_2
X_07883_ _07883_/A vssd1 vssd1 vccd1 vccd1 _07885_/A sky130_fd_sc_hd__inv_2
X_06834_ _06833_/B _08772_/B _06834_/C vssd1 vssd1 vccd1 vccd1 _08772_/A sky130_fd_sc_hd__nand3b_1
X_09622_ _10112_/A _10108_/B input19/X input20/X vssd1 vssd1 vccd1 vccd1 _09622_/X
+ sky130_fd_sc_hd__and4_1
X_09553_ _09553_/A _09786_/B _09554_/B vssd1 vssd1 vccd1 vccd1 _09800_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_77_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06765_ _06769_/C vssd1 vssd1 vccd1 vccd1 _06766_/C sky130_fd_sc_hd__inv_2
X_08504_ _08506_/A vssd1 vssd1 vccd1 vccd1 _08505_/B sky130_fd_sc_hd__inv_2
XFILLER_0_77_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09484_ _09486_/B _09486_/A vssd1 vssd1 vccd1 vccd1 _09485_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_65_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05716_ _05547_/Y _05716_/B _05716_/C vssd1 vssd1 vccd1 vccd1 _06121_/B sky130_fd_sc_hd__nand3b_1
X_06696_ _06696_/A _06696_/B vssd1 vssd1 vccd1 vccd1 _06697_/A sky130_fd_sc_hd__nand2_1
X_08435_ _08435_/A _08435_/B vssd1 vssd1 vccd1 vccd1 _08558_/B sky130_fd_sc_hd__nand2_1
X_05647_ _05647_/A vssd1 vssd1 vccd1 vccd1 _05648_/B sky130_fd_sc_hd__inv_2
X_08366_ _08369_/B _08366_/B vssd1 vssd1 vccd1 vccd1 _08367_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05578_ _05578_/A _05578_/B vssd1 vssd1 vccd1 vccd1 _05709_/C sky130_fd_sc_hd__nand2_1
X_07317_ _07320_/B vssd1 vssd1 vccd1 vccd1 _07322_/B sky130_fd_sc_hd__inv_2
XFILLER_0_18_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08297_ _08269_/Y _08297_/B vssd1 vssd1 vccd1 vccd1 _08331_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07248_ _07287_/A _07289_/A vssd1 vssd1 vccd1 vccd1 _07248_/Y sky130_fd_sc_hd__nor2_1
X_07179_ _07351_/C vssd1 vssd1 vccd1 vccd1 _07181_/B sky130_fd_sc_hd__inv_2
X_10190_ _10190_/A _10190_/B vssd1 vssd1 vccd1 vccd1 _10191_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06149__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput27 a_i[4] vssd1 vssd1 vccd1 vccd1 input27/X sky130_fd_sc_hd__buf_1
Xinput16 a_i[23] vssd1 vssd1 vccd1 vccd1 input16/X sky130_fd_sc_hd__clkbuf_1
Xinput49 b_i[24] vssd1 vssd1 vccd1 vccd1 input49/X sky130_fd_sc_hd__buf_4
Xinput38 b_i[14] vssd1 vssd1 vccd1 vccd1 input38/X sky130_fd_sc_hd__buf_2
X_10526_ _10526_/A _10532_/A vssd1 vssd1 vccd1 vccd1 _10527_/A sky130_fd_sc_hd__nand2_1
X_10457_ _10449_/A _10457_/B vssd1 vssd1 vccd1 vccd1 _10542_/A sky130_fd_sc_hd__nand2b_1
XANTENNA__09754__A2 _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10388_ _10390_/B _10390_/C vssd1 vssd1 vccd1 vccd1 _10389_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06550_ _06553_/B _06553_/C vssd1 vssd1 vccd1 vccd1 _06552_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06481_ _06481_/A _06481_/B vssd1 vssd1 vccd1 vccd1 _06603_/C sky130_fd_sc_hd__nand2_1
X_05501_ _05501_/A _05501_/B vssd1 vssd1 vccd1 vccd1 _05501_/Y sky130_fd_sc_hd__nor2_1
X_05432_ input63/X vssd1 vssd1 vccd1 vccd1 _07897_/B sky130_fd_sc_hd__buf_4
X_08220_ _08222_/B _08225_/A vssd1 vssd1 vccd1 vccd1 _08224_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08151_ _08151_/A _08280_/A vssd1 vssd1 vccd1 vccd1 _08245_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05363_ _05394_/C vssd1 vssd1 vccd1 vccd1 _05396_/B sky130_fd_sc_hd__inv_2
X_08082_ _08084_/A _08384_/A vssd1 vssd1 vccd1 vccd1 _08087_/A sky130_fd_sc_hd__nand2_1
X_07102_ _07118_/C vssd1 vssd1 vccd1 vccd1 _07117_/B sky130_fd_sc_hd__inv_2
X_07033_ _07031_/Y _07024_/B _07032_/Y vssd1 vssd1 vccd1 vccd1 _07075_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_11_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08984_ _08984_/A vssd1 vssd1 vccd1 vccd1 _08985_/B sky130_fd_sc_hd__inv_2
XFILLER_0_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07935_ _07935_/A _07975_/C vssd1 vssd1 vccd1 vccd1 _07937_/A sky130_fd_sc_hd__nand2_1
X_09605_ _10151_/A _10148_/B _10150_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _10012_/A
+ sky130_fd_sc_hd__a22o_1
X_07866_ _07871_/A _07867_/A vssd1 vssd1 vccd1 vccd1 _07870_/A sky130_fd_sc_hd__nand2_1
X_06817_ _06817_/A _08881_/A _06817_/C vssd1 vssd1 vccd1 vccd1 _06818_/B sky130_fd_sc_hd__nand3_1
X_07797_ _07797_/A _07797_/B _07797_/C vssd1 vssd1 vccd1 vccd1 _07798_/B sky130_fd_sc_hd__nand3_1
X_09536_ _09536_/A vssd1 vssd1 vccd1 vccd1 _09771_/A sky130_fd_sc_hd__inv_2
XFILLER_0_78_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06748_ _09971_/A _08633_/B _06744_/Y vssd1 vssd1 vccd1 vccd1 _06753_/B sky130_fd_sc_hd__o21ai_1
X_09467_ _09466_/B _09467_/B _09692_/B vssd1 vssd1 vccd1 vccd1 _09692_/A sky130_fd_sc_hd__nand3b_1
X_08418_ _08418_/A vssd1 vssd1 vccd1 vccd1 _08420_/B sky130_fd_sc_hd__inv_2
X_06679_ _06679_/A _06679_/B _06679_/C vssd1 vssd1 vccd1 vccd1 _06938_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09398_ _09611_/B _09403_/C vssd1 vssd1 vccd1 vccd1 _09401_/A sky130_fd_sc_hd__nand2_1
X_08349_ _08349_/A _08349_/B _08355_/B vssd1 vssd1 vccd1 vccd1 _08354_/A sky130_fd_sc_hd__nand3_1
XANTENNA__10043__A2 _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10311_ _10311_/A _10311_/B vssd1 vssd1 vccd1 vccd1 _10314_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10242_ _10242_/A _10242_/B vssd1 vssd1 vccd1 vccd1 _10314_/A sky130_fd_sc_hd__nand2_1
X_10173_ _10173_/A _10173_/B vssd1 vssd1 vccd1 vccd1 _10176_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10129__A _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06326__B _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10509_ _10649_/B _10652_/A _10652_/B vssd1 vssd1 vccd1 vccd1 _10510_/B sky130_fd_sc_hd__nand3_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07157__B _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05981_ _05598_/B _05598_/C _05966_/B vssd1 vssd1 vccd1 vccd1 _05982_/B sky130_fd_sc_hd__a21boi_1
X_07720_ _07842_/B _08075_/A vssd1 vssd1 vccd1 vccd1 _08084_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07651_ _07653_/C vssd1 vssd1 vccd1 vccd1 _07809_/A sky130_fd_sc_hd__inv_2
XANTENNA__07173__A _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07582_ _07582_/A _07582_/B vssd1 vssd1 vccd1 vccd1 _07594_/B sky130_fd_sc_hd__nand2_1
X_06602_ _06602_/A _06602_/B _06602_/C vssd1 vssd1 vccd1 vccd1 _06603_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10030__C _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09321_ _09587_/A _09321_/B _09351_/A vssd1 vssd1 vccd1 vccd1 _09322_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_47_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06533_ _06653_/B _06653_/C _06532_/Y vssd1 vssd1 vccd1 vccd1 _06659_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09252_ _09278_/A _09278_/C vssd1 vssd1 vccd1 vccd1 _09277_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06464_ _06466_/A vssd1 vssd1 vccd1 vccd1 _06465_/B sky130_fd_sc_hd__inv_2
XFILLER_0_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09183_ _08623_/C _08623_/A _09185_/B vssd1 vssd1 vccd1 vccd1 _09184_/B sky130_fd_sc_hd__a21boi_1
X_08203_ _08203_/A _08203_/B vssd1 vssd1 vccd1 vccd1 _08207_/A sky130_fd_sc_hd__nand2_1
X_06395_ _06557_/C _06557_/B _06394_/Y vssd1 vssd1 vccd1 vccd1 _06401_/A sky130_fd_sc_hd__a21oi_1
X_05415_ _05415_/A _05416_/A vssd1 vssd1 vccd1 vccd1 _05418_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08134_ _08155_/B _08134_/B vssd1 vssd1 vccd1 vccd1 _08203_/B sky130_fd_sc_hd__and2_1
X_05346_ _05353_/B _05476_/A vssd1 vssd1 vccd1 vccd1 _05352_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08065_ _07815_/Y _07967_/B _07816_/Y vssd1 vssd1 vccd1 vccd1 _08066_/A sky130_fd_sc_hd__a21o_1
X_07016_ _10040_/B _07891_/B vssd1 vssd1 vccd1 vccd1 _07184_/B sky130_fd_sc_hd__nand2_1
X_08967_ _08967_/A _08967_/B _08967_/C vssd1 vssd1 vccd1 vccd1 _09025_/C sky130_fd_sc_hd__nand3_1
X_08898_ _08898_/A vssd1 vssd1 vccd1 vccd1 _08903_/B sky130_fd_sc_hd__inv_2
X_07918_ _07918_/A _07918_/B vssd1 vssd1 vccd1 vccd1 _07919_/A sky130_fd_sc_hd__nand2_1
X_07849_ _07849_/A _07852_/A _07849_/C vssd1 vssd1 vccd1 vccd1 _07849_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09519_ input49/X _09840_/B input50/X _09749_/B vssd1 vssd1 vccd1 vccd1 _09520_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10225_ _10227_/C vssd1 vssd1 vccd1 vccd1 _10226_/B sky130_fd_sc_hd__inv_2
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08393__A1 _09201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10156_ _10156_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _10160_/A sky130_fd_sc_hd__nand2_1
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ _10087_/A _10087_/B _10087_/C vssd1 vssd1 vccd1 vccd1 _10089_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_55_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_106 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10007__A2 _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06180_ _06221_/B _06221_/C vssd1 vssd1 vccd1 vccd1 _06220_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09870_ _09870_/A _09870_/B _10305_/A vssd1 vssd1 vccd1 vccd1 _09893_/B sky130_fd_sc_hd__nand3_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _08871_/A _08872_/C vssd1 vssd1 vccd1 vccd1 _08821_/Y sky130_fd_sc_hd__nand2_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08752_ _08754_/B vssd1 vssd1 vccd1 vccd1 _08753_/B sky130_fd_sc_hd__inv_2
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05964_ _06821_/A _05964_/B _05964_/C vssd1 vssd1 vccd1 vccd1 _06013_/B sky130_fd_sc_hd__nand3_1
X_08683_ _08683_/A _08683_/B vssd1 vssd1 vccd1 vccd1 _08763_/A sky130_fd_sc_hd__nand2_1
X_07703_ _07736_/B vssd1 vssd1 vccd1 vccd1 _07733_/B sky130_fd_sc_hd__inv_2
X_05895_ _05530_/C _05530_/B _05894_/Y vssd1 vssd1 vccd1 vccd1 _06821_/A sky130_fd_sc_hd__a21oi_2
X_07634_ _07637_/A _07637_/B vssd1 vssd1 vccd1 vccd1 _07777_/A sky130_fd_sc_hd__or2_1
XFILLER_0_75_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07565_ _07565_/A _07565_/B vssd1 vssd1 vccd1 vccd1 _07835_/A sky130_fd_sc_hd__nand2_1
X_09304_ _09309_/A _09572_/A vssd1 vssd1 vccd1 vccd1 _09308_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ _07496_/A _07496_/B vssd1 vssd1 vccd1 vccd1 _07498_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06516_ _10212_/B _10101_/A vssd1 vssd1 vccd1 vccd1 _06640_/C sky130_fd_sc_hd__nand2_1
X_09235_ _09236_/B _09236_/A vssd1 vssd1 vccd1 vccd1 _09469_/A sky130_fd_sc_hd__or2_1
X_06447_ _08114_/B _10187_/A vssd1 vssd1 vccd1 vccd1 _06623_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_16_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09166_ _09971_/A _09912_/B _09165_/C vssd1 vssd1 vccd1 vccd1 _09166_/Y sky130_fd_sc_hd__o21ai_1
X_06378_ _06380_/B _06379_/B _06379_/A vssd1 vssd1 vccd1 vccd1 _06489_/B sky130_fd_sc_hd__nand3b_1
X_09097_ _08742_/Y _08745_/B _08743_/A vssd1 vssd1 vccd1 vccd1 _09103_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_9_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08117_ _08167_/B _08169_/B _08116_/Y vssd1 vssd1 vccd1 vccd1 _08118_/C sky130_fd_sc_hd__a21oi_1
X_08048_ _08048_/A _08048_/B vssd1 vssd1 vccd1 vccd1 _08148_/A sky130_fd_sc_hd__nand2_1
X_10010_ _10010_/A _10010_/B vssd1 vssd1 vccd1 vccd1 _10019_/B sky130_fd_sc_hd__nand2_1
X_09999_ _10001_/A vssd1 vssd1 vccd1 vccd1 _10000_/B sky130_fd_sc_hd__inv_2
XFILLER_0_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10208_ _10208_/A vssd1 vssd1 vccd1 vccd1 _10208_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_66_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10139_ _10140_/B _10140_/A vssd1 vssd1 vccd1 vccd1 _10141_/A sky130_fd_sc_hd__or2_1
XFILLER_0_82_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05680_ _05680_/A vssd1 vssd1 vccd1 vccd1 _05683_/A sky130_fd_sc_hd__inv_2
X_07350_ _07350_/A _07350_/B vssd1 vssd1 vccd1 vccd1 _07351_/B sky130_fd_sc_hd__nand2_1
X_06301_ _06302_/B _06302_/A vssd1 vssd1 vccd1 vccd1 _06310_/B sky130_fd_sc_hd__nor2_1
X_09020_ _09020_/A _09020_/B vssd1 vssd1 vccd1 vccd1 _09053_/B sky130_fd_sc_hd__nand2_1
X_07281_ _10406_/B _10409_/A _10404_/A vssd1 vssd1 vccd1 vccd1 _07286_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_72_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06232_ _06234_/A vssd1 vssd1 vccd1 vccd1 _06233_/B sky130_fd_sc_hd__inv_2
XFILLER_0_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_183 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06163_ _06166_/B _06166_/C vssd1 vssd1 vccd1 vccd1 _06165_/A sky130_fd_sc_hd__nand2_1
X_06094_ _06927_/B vssd1 vssd1 vccd1 vccd1 _06928_/C sky130_fd_sc_hd__inv_2
XFILLER_0_40_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09922_ _10148_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _09923_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09853_ _09853_/A _09853_/B vssd1 vssd1 vccd1 vccd1 _09855_/A sky130_fd_sc_hd__nand2_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _09873_/A _09784_/B vssd1 vssd1 vccd1 vccd1 _09786_/A sky130_fd_sc_hd__nand2_1
X_08804_ _08815_/A vssd1 vssd1 vccd1 vccd1 _08805_/B sky130_fd_sc_hd__inv_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08735_ _08750_/C vssd1 vssd1 vccd1 vccd1 _08735_/Y sky130_fd_sc_hd__inv_2
XANTENNA__09841__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _06996_/A vssd1 vssd1 vccd1 vccd1 _06998_/B sky130_fd_sc_hd__inv_2
X_05947_ _05952_/A _06760_/A vssd1 vssd1 vccd1 vccd1 _06804_/B sky130_fd_sc_hd__nand2_1
X_08666_ _09134_/B _08666_/B _08666_/C vssd1 vssd1 vccd1 vccd1 _09134_/A sky130_fd_sc_hd__nand3_2
X_05878_ _06200_/B _06199_/A _06199_/B vssd1 vssd1 vccd1 vccd1 _06202_/B sky130_fd_sc_hd__nand3b_1
X_08597_ _09156_/B _08597_/B _08597_/C vssd1 vssd1 vccd1 vccd1 _09156_/A sky130_fd_sc_hd__nand3_1
X_07617_ _07617_/A _07617_/B vssd1 vssd1 vccd1 vccd1 _07618_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07548_ _07548_/A _07548_/B vssd1 vssd1 vccd1 vccd1 _07664_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08176__B _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07479_ _10292_/B _10151_/A vssd1 vssd1 vccd1 vccd1 _07618_/B sky130_fd_sc_hd__nand2_1
X_09218_ _09217_/B _09218_/B _09218_/C vssd1 vssd1 vccd1 vccd1 _09219_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_51_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10713__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10490_ _10490_/A _10490_/B vssd1 vssd1 vccd1 vccd1 _10493_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_8_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09149_ _09393_/C _09149_/B vssd1 vssd1 vccd1 vccd1 _09151_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09454__C _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10688_ _10688_/A _10690_/A vssd1 vssd1 vccd1 vccd1 _10689_/A sky130_fd_sc_hd__and2_1
XFILLER_0_2_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06334__B _07785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09645__B _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06850_ _06850_/A _06850_/B _08983_/A vssd1 vssd1 vccd1 vccd1 _06881_/C sky130_fd_sc_hd__nand3_1
X_05801_ _05801_/A _05801_/B vssd1 vssd1 vccd1 vccd1 _05802_/B sky130_fd_sc_hd__nand2_1
X_06781_ _06780_/B _08769_/B _06781_/C vssd1 vssd1 vccd1 vccd1 _08769_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_77_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05732_ _05738_/C vssd1 vssd1 vccd1 vccd1 _05732_/Y sky130_fd_sc_hd__inv_2
X_08520_ _08520_/A vssd1 vssd1 vccd1 vccd1 _08521_/A sky130_fd_sc_hd__inv_2
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08451_ _08817_/B _08817_/C vssd1 vssd1 vccd1 vccd1 _08463_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05663_ _05663_/A _05663_/B vssd1 vssd1 vccd1 vccd1 _06124_/A sky130_fd_sc_hd__nand2_1
X_07402_ _07400_/Y _07368_/B _07401_/Y vssd1 vssd1 vccd1 vccd1 _07403_/B sky130_fd_sc_hd__a21o_1
X_05594_ _08672_/A vssd1 vssd1 vccd1 vccd1 _10212_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08382_ _08382_/A _08382_/B vssd1 vssd1 vccd1 vccd1 _08383_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07333_ _10210_/B _10103_/B vssd1 vssd1 vccd1 vccd1 _07353_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07264_ _07264_/A vssd1 vssd1 vccd1 vccd1 _07265_/B sky130_fd_sc_hd__inv_2
X_09003_ _09003_/A _09003_/B vssd1 vssd1 vccd1 vccd1 _09009_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_26_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06215_ _06217_/A vssd1 vssd1 vccd1 vccd1 _06216_/B sky130_fd_sc_hd__inv_2
XFILLER_0_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07195_ _07206_/B _07195_/B _07195_/C vssd1 vssd1 vccd1 vccd1 _07206_/A sky130_fd_sc_hd__nand3_1
XANTENNA__08740__A _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06146_ _06255_/B _06255_/C _06145_/Y vssd1 vssd1 vccd1 vccd1 _06234_/A sky130_fd_sc_hd__a21oi_2
X_06077_ _06078_/B _06078_/A vssd1 vssd1 vccd1 vccd1 _06077_/Y sky130_fd_sc_hd__nand2_1
X_09905_ _09907_/B vssd1 vssd1 vccd1 vccd1 _09906_/B sky130_fd_sc_hd__inv_2
X_09836_ _09836_/A _09836_/B vssd1 vssd1 vccd1 vccd1 _09837_/A sky130_fd_sc_hd__nand2_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ _09763_/Y _09765_/Y _09768_/B vssd1 vssd1 vccd1 vccd1 _09775_/A sky130_fd_sc_hd__o21bai_1
X_06979_ _10108_/B _10201_/A vssd1 vssd1 vccd1 vccd1 _07143_/A sky130_fd_sc_hd__nand2_1
X_08718_ _09710_/B _09698_/A vssd1 vssd1 vccd1 vccd1 _08722_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09698_ _09698_/A vssd1 vssd1 vccd1 vccd1 _10202_/D sky130_fd_sc_hd__inv_2
XFILLER_0_68_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08649_ _09201_/A _10006_/A _08648_/C vssd1 vssd1 vccd1 vccd1 _08650_/A sky130_fd_sc_hd__o21ai_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _10611_/A hold20/X vssd1 vssd1 vccd1 vccd1 _10616_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10542_ _10542_/A _10542_/B vssd1 vssd1 vccd1 vccd1 _10544_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_51_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10473_ _10476_/A _10476_/C vssd1 vssd1 vccd1 vccd1 _10475_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08097__A _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05514__A _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06329__B _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06048__C _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06064__B _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06000_ _06001_/B _06001_/A vssd1 vssd1 vccd1 vccd1 _06000_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_2_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_167 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07951_ _07951_/A _07951_/B _07951_/C vssd1 vssd1 vccd1 vccd1 _07952_/B sky130_fd_sc_hd__nand3_1
X_06902_ _06902_/A _06902_/B vssd1 vssd1 vccd1 vccd1 _06902_/Y sky130_fd_sc_hd__nor2_1
X_07882_ _07883_/A _07884_/A vssd1 vssd1 vccd1 vccd1 _07913_/C sky130_fd_sc_hd__nand2_1
X_06833_ _06833_/A _06833_/B vssd1 vssd1 vccd1 vccd1 _06839_/A sky130_fd_sc_hd__nand2_1
X_09621_ _10115_/A input21/X vssd1 vssd1 vccd1 vccd1 _09626_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_37_83 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09552_ input52/X _10284_/B input53/X _10292_/B vssd1 vssd1 vccd1 vccd1 _09554_/B
+ sky130_fd_sc_hd__a22o_1
X_06764_ _06764_/A _08819_/A vssd1 vssd1 vccd1 vccd1 _06769_/C sky130_fd_sc_hd__nand2_1
X_05715_ _05547_/Y _05714_/Y _05546_/A vssd1 vssd1 vccd1 vccd1 _06121_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__05424__A _07891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08503_ _08476_/B _08476_/A _08474_/A vssd1 vssd1 vccd1 vccd1 _08506_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09483_ _09705_/A _09483_/B vssd1 vssd1 vccd1 vccd1 _09486_/A sky130_fd_sc_hd__nand2_1
X_06695_ _07274_/C vssd1 vssd1 vccd1 vccd1 _07273_/B sky130_fd_sc_hd__inv_2
XFILLER_0_65_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08434_ _08555_/A _08556_/A vssd1 vssd1 vccd1 vccd1 _08434_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05646_ _05646_/A vssd1 vssd1 vccd1 vccd1 _05648_/A sky130_fd_sc_hd__inv_2
X_05577_ _05577_/A _05577_/B _05577_/C vssd1 vssd1 vccd1 vccd1 _05578_/B sky130_fd_sc_hd__nand3_1
X_08365_ _08365_/A _08376_/B vssd1 vssd1 vccd1 vccd1 _08369_/B sky130_fd_sc_hd__and2_1
XFILLER_0_18_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08454__B _09201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07316_ _07500_/B _07500_/C vssd1 vssd1 vccd1 vccd1 _07502_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08296_ _08296_/A vssd1 vssd1 vccd1 vccd1 _08356_/A sky130_fd_sc_hd__inv_2
X_07247_ _07429_/B _07293_/B vssd1 vssd1 vccd1 vccd1 _07291_/B sky130_fd_sc_hd__nor2b_1
XFILLER_0_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07178_ _10247_/B _10128_/A vssd1 vssd1 vccd1 vccd1 _07351_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08470__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06129_ _06280_/A _06281_/B vssd1 vssd1 vccd1 vccd1 _06284_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07086__A _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09819_ _09818_/B _09819_/B _09835_/B vssd1 vssd1 vccd1 vccd1 _09835_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__08645__A _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput28 a_i[5] vssd1 vssd1 vccd1 vccd1 input28/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xinput17 a_i[24] vssd1 vssd1 vccd1 vccd1 input17/X sky130_fd_sc_hd__buf_2
Xinput39 b_i[15] vssd1 vssd1 vccd1 vccd1 input39/X sky130_fd_sc_hd__clkbuf_2
X_10525_ _10525_/A _10525_/B vssd1 vssd1 vccd1 vccd1 _10532_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09476__A _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10456_ _10456_/A _10456_/B vssd1 vssd1 vccd1 vccd1 _10667_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09754__A3 _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10387_ _10390_/B hold28/X _10387_/C vssd1 vssd1 vccd1 vccd1 _10690_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10150__A _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06480_ _06480_/A _06480_/B vssd1 vssd1 vccd1 vccd1 _06481_/B sky130_fd_sc_hd__nand2_1
X_05500_ _05501_/B _05501_/A vssd1 vssd1 vccd1 vccd1 _05500_/Y sky130_fd_sc_hd__nand2_1
X_05431_ _05524_/B _05437_/C vssd1 vssd1 vccd1 vccd1 _05435_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08150_ _08211_/A _08212_/B _08212_/A vssd1 vssd1 vccd1 vccd1 _08280_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_15_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07101_ _07101_/A _07106_/A vssd1 vssd1 vccd1 vccd1 _07118_/C sky130_fd_sc_hd__nand2_1
X_05362_ _08114_/B _10150_/B vssd1 vssd1 vccd1 vccd1 _05394_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08081_ _08081_/A _08238_/A _08238_/B vssd1 vssd1 vccd1 vccd1 _10493_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_15_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09386__A _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07032_ _07032_/A _07032_/B vssd1 vssd1 vccd1 vccd1 _07032_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_70_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08983_ _08983_/A _08983_/B vssd1 vssd1 vccd1 vccd1 _08985_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07934_ _07936_/C vssd1 vssd1 vccd1 vccd1 _07975_/C sky130_fd_sc_hd__inv_2
X_07865_ _07868_/B vssd1 vssd1 vccd1 vccd1 _07871_/A sky130_fd_sc_hd__inv_2
X_09604_ _09604_/A vssd1 vssd1 vccd1 vccd1 _09606_/A sky130_fd_sc_hd__inv_2
XFILLER_0_3_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06816_ _06816_/A _06816_/B vssd1 vssd1 vccd1 vccd1 _06818_/A sky130_fd_sc_hd__nand2_1
X_07796_ _07796_/A vssd1 vssd1 vccd1 vccd1 _07797_/C sky130_fd_sc_hd__inv_2
X_09535_ _09771_/B _09536_/A vssd1 vssd1 vccd1 vccd1 _09542_/B sky130_fd_sc_hd__nand2_1
X_06747_ _10148_/B vssd1 vssd1 vccd1 vccd1 _08633_/B sky130_fd_sc_hd__inv_2
X_09466_ _09466_/A _09466_/B vssd1 vssd1 vccd1 vccd1 _09474_/A sky130_fd_sc_hd__nand2_1
X_06678_ _06678_/A _06678_/B vssd1 vssd1 vccd1 vccd1 _06938_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08417_ _08421_/B _08660_/B _08417_/C vssd1 vssd1 vccd1 vccd1 _08660_/A sky130_fd_sc_hd__nand3b_1
X_05629_ _06016_/B _05629_/B _05629_/C vssd1 vssd1 vccd1 vccd1 _06106_/B sky130_fd_sc_hd__nand3_2
XANTENNA__10028__B1 _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09397_ _09397_/A _09397_/B _09397_/C vssd1 vssd1 vccd1 vccd1 _09403_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_46_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08348_ _08349_/B _08355_/B _08349_/A vssd1 vssd1 vccd1 vccd1 _08356_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08279_ _08324_/B _08324_/A vssd1 vssd1 vccd1 vccd1 _08282_/A sky130_fd_sc_hd__nor2_1
X_10310_ _10310_/A _10310_/B _10310_/C vssd1 vssd1 vccd1 vccd1 _10311_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10241_ _10243_/A vssd1 vssd1 vccd1 vccd1 _10242_/B sky130_fd_sc_hd__inv_2
X_10172_ _10171_/B _10172_/B _10172_/C vssd1 vssd1 vccd1 vccd1 _10173_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_69_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10508_ _10508_/A vssd1 vssd1 vccd1 vccd1 _10649_/B sky130_fd_sc_hd__inv_2
XFILLER_0_12_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10439_ hold25/X vssd1 vssd1 vccd1 vccd1 _10440_/B sky130_fd_sc_hd__inv_2
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05980_ _05980_/A _06796_/A vssd1 vssd1 vccd1 vccd1 _05982_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07650_ _07875_/A _07808_/A vssd1 vssd1 vccd1 vccd1 _07653_/C sky130_fd_sc_hd__nor2_1
XANTENNA__07173__B _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ _07250_/Y _07429_/B _07251_/Y vssd1 vssd1 vccd1 vccd1 _07582_/B sky130_fd_sc_hd__a21o_1
X_06601_ _06601_/A _06601_/B vssd1 vssd1 vccd1 vccd1 _06603_/A sky130_fd_sc_hd__nand2_1
X_09320_ _09351_/B _09320_/B vssd1 vssd1 vccd1 vccd1 _09322_/A sky130_fd_sc_hd__nand2_1
X_06532_ _06650_/A _06649_/A vssd1 vssd1 vccd1 vccd1 _06532_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_34_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09251_ _09471_/A _09251_/B _09251_/C vssd1 vssd1 vccd1 vccd1 _09278_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08202_ _08204_/B _08204_/C vssd1 vssd1 vccd1 vccd1 _08203_/A sky130_fd_sc_hd__nand2_1
X_06463_ _06610_/A _06605_/A vssd1 vssd1 vccd1 vccd1 _06463_/Y sky130_fd_sc_hd__nand2_1
X_09182_ _09186_/B _09409_/A vssd1 vssd1 vccd1 vccd1 _09184_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06394_ _06394_/A _06394_/B vssd1 vssd1 vccd1 vccd1 _06394_/Y sky130_fd_sc_hd__nor2_1
X_05414_ _08101_/B input6/X vssd1 vssd1 vccd1 vccd1 _05416_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08133_ _08133_/A _08133_/B vssd1 vssd1 vccd1 vccd1 _08134_/B sky130_fd_sc_hd__nand2_1
X_05345_ _08573_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _05476_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_70_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08064_ _08064_/A _08064_/B vssd1 vssd1 vccd1 vccd1 _08233_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_70_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07015_ _07183_/B vssd1 vssd1 vccd1 vccd1 _07184_/A sky130_fd_sc_hd__inv_2
XANTENNA__10738__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ _08966_/A _08966_/B vssd1 vssd1 vccd1 vccd1 _09025_/B sky130_fd_sc_hd__nand2_1
X_08897_ input51/X _08897_/B vssd1 vssd1 vccd1 vccd1 _08898_/A sky130_fd_sc_hd__nand2_1
X_07917_ _07917_/A vssd1 vssd1 vccd1 vccd1 _07918_/B sky130_fd_sc_hd__inv_2
X_07848_ _07848_/A _07850_/B _07848_/C vssd1 vssd1 vccd1 vccd1 _07849_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ _09518_/A vssd1 vssd1 vccd1 vccd1 _09759_/B sky130_fd_sc_hd__inv_2
XANTENNA__10249__B1 input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07811__B _07811_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ _07783_/A _07783_/C vssd1 vssd1 vccd1 vccd1 _07781_/A sky130_fd_sc_hd__nand2_1
X_09449_ _09449_/A _09449_/B vssd1 vssd1 vccd1 vccd1 _09450_/B sky130_fd_sc_hd__and2_1
XFILLER_0_38_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06443__A _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10224_ _10222_/Y _09936_/Y _10223_/Y vssd1 vssd1 vccd1 vccd1 _10227_/C sky130_fd_sc_hd__a21oi_1
X_10155_ _10155_/A _10155_/B vssd1 vssd1 vccd1 vccd1 _10161_/A sky130_fd_sc_hd__and2_1
X_10086_ _10086_/A vssd1 vssd1 vccd1 vccd1 _10087_/B sky130_fd_sc_hd__inv_2
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _08871_/B vssd1 vssd1 vccd1 vccd1 _08872_/C sky130_fd_sc_hd__inv_2
XFILLER_0_0_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08751_ _08751_/A _08751_/B vssd1 vssd1 vccd1 vccd1 _08754_/B sky130_fd_sc_hd__nand2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05963_ _05963_/A _06821_/B vssd1 vssd1 vccd1 vccd1 _06013_/A sky130_fd_sc_hd__nand2_1
X_08682_ _08692_/C vssd1 vssd1 vccd1 vccd1 _08683_/B sky130_fd_sc_hd__inv_2
X_05894_ _05894_/A _05894_/B vssd1 vssd1 vccd1 vccd1 _05894_/Y sky130_fd_sc_hd__nor2_1
X_07702_ _07702_/A _07702_/B vssd1 vssd1 vccd1 vccd1 _07736_/B sky130_fd_sc_hd__nand2_1
X_07633_ _09749_/B _10129_/A vssd1 vssd1 vccd1 vccd1 _07637_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07564_ _07566_/A vssd1 vssd1 vccd1 vccd1 _07565_/B sky130_fd_sc_hd__inv_2
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09303_ _09308_/B _09572_/A _09309_/A vssd1 vssd1 vccd1 vccd1 _09583_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07495_ _07644_/C _07617_/B vssd1 vssd1 vccd1 vccd1 _07496_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06515_ _08101_/B vssd1 vssd1 vccd1 vccd1 _10101_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09234_ _09234_/A _09234_/B vssd1 vssd1 vccd1 vccd1 _09236_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_63_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06446_ _06621_/A _06622_/B vssd1 vssd1 vccd1 vccd1 _06625_/C sky130_fd_sc_hd__nand2_1
X_09165_ _09971_/A _09912_/B _09165_/C vssd1 vssd1 vccd1 vccd1 _09400_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08116_ _08164_/A _08165_/A vssd1 vssd1 vccd1 vccd1 _08116_/Y sky130_fd_sc_hd__nor2_1
X_06377_ _06377_/A _06377_/B vssd1 vssd1 vccd1 vccd1 _06379_/A sky130_fd_sc_hd__nand2_1
X_09096_ _09096_/A _09096_/B vssd1 vssd1 vccd1 vccd1 _09539_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07359__A _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08047_ _08047_/A _08047_/B vssd1 vssd1 vccd1 vccd1 _08048_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09998_ _09998_/A _09998_/B vssd1 vssd1 vccd1 vccd1 _10001_/A sky130_fd_sc_hd__nand2_1
X_08949_ _08949_/A _08949_/B vssd1 vssd1 vccd1 vccd1 _08950_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05607__A input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09627__A2 _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09749__A input51/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10207_ _10209_/B _10209_/A vssd1 vssd1 vccd1 vccd1 _10208_/A sky130_fd_sc_hd__nor2_1
X_10138_ _10125_/Y _10126_/X _10141_/B vssd1 vssd1 vccd1 vccd1 _10146_/A sky130_fd_sc_hd__o21bai_1
X_10069_ _10073_/B _10073_/C vssd1 vssd1 vccd1 vccd1 _10072_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_82_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06348__A _08725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06300_ _06300_/A _06300_/B vssd1 vssd1 vccd1 vccd1 _06302_/A sky130_fd_sc_hd__and2_1
X_07280_ _10431_/C _07276_/Y _07859_/A vssd1 vssd1 vccd1 vccd1 _10404_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06231_ _06315_/B _06315_/C vssd1 vssd1 vccd1 vccd1 _06314_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06162_ _06162_/A _06162_/B _06162_/C vssd1 vssd1 vccd1 vccd1 _06166_/C sky130_fd_sc_hd__nand3_1
X_06093_ _06095_/B _06095_/A vssd1 vssd1 vccd1 vccd1 _06927_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_13_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_195 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09921_ _09921_/A _09921_/B vssd1 vssd1 vccd1 vccd1 _09930_/C sky130_fd_sc_hd__nand2_1
X_09852_ _09855_/B _09852_/B _09852_/C vssd1 vssd1 vccd1 vccd1 _09862_/B sky130_fd_sc_hd__nand3b_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08803_ _08803_/A _08803_/B vssd1 vssd1 vccd1 vccd1 _08815_/A sky130_fd_sc_hd__nand2_1
X_09783_ _09782_/A _09782_/B _09782_/C vssd1 vssd1 vccd1 vccd1 _09784_/B sky130_fd_sc_hd__o21ai_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05427__A _07785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _08734_/A _08734_/B vssd1 vssd1 vccd1 vccd1 _08750_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_56_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ _06995_/A _06995_/B vssd1 vssd1 vccd1 vccd1 _06998_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08738__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05946_ _05945_/B _06760_/B _05946_/C vssd1 vssd1 vccd1 vccd1 _06760_/A sky130_fd_sc_hd__nand3b_1
X_08665_ _08665_/A vssd1 vssd1 vccd1 vccd1 _08666_/B sky130_fd_sc_hd__inv_2
X_05877_ _05877_/A _05877_/B vssd1 vssd1 vccd1 vccd1 _06199_/B sky130_fd_sc_hd__nand2_1
X_08596_ _08596_/A vssd1 vssd1 vccd1 vccd1 _08597_/B sky130_fd_sc_hd__inv_2
X_07616_ _07714_/A _07616_/B vssd1 vssd1 vccd1 vccd1 _07823_/B sky130_fd_sc_hd__nand2_1
X_07547_ _07547_/A _07547_/B _07547_/C vssd1 vssd1 vccd1 vccd1 _07548_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08223__A_N _08363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07478_ _07497_/B _07497_/C vssd1 vssd1 vccd1 vccd1 _07496_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09217_ _09217_/A _09217_/B vssd1 vssd1 vccd1 vccd1 _09219_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_395 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06429_ _06602_/B _06602_/C vssd1 vssd1 vccd1 vccd1 _06601_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07089__A _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ _10103_/A input20/X vssd1 vssd1 vccd1 vccd1 _09149_/B sky130_fd_sc_hd__nand2_1
X_09079_ _09079_/A vssd1 vssd1 vccd1 vccd1 _10370_/A sky130_fd_sc_hd__inv_2
XFILLER_0_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09454__D _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08648__A _09201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10687_ _10687_/A _10687_/B vssd1 vssd1 vccd1 vccd1 _10690_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06631__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05800_ _05800_/A vssd1 vssd1 vccd1 vccd1 _05802_/A sky130_fd_sc_hd__inv_2
X_06780_ _06780_/A _06780_/B vssd1 vssd1 vccd1 vccd1 _06782_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05731_ _05731_/A _05731_/B vssd1 vssd1 vccd1 vccd1 _05738_/C sky130_fd_sc_hd__nand2_1
X_08450_ _08450_/A _08450_/B _08450_/C vssd1 vssd1 vccd1 vccd1 _08817_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05662_ _05664_/B vssd1 vssd1 vccd1 vccd1 _05663_/B sky130_fd_sc_hd__inv_2
XFILLER_0_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07401_ _07401_/A _07401_/B vssd1 vssd1 vccd1 vccd1 _07401_/Y sky130_fd_sc_hd__nor2_1
X_08381_ _08381_/A vssd1 vssd1 vccd1 vccd1 _10472_/C sky130_fd_sc_hd__inv_4
XFILLER_0_73_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05593_ _05966_/B _05598_/C vssd1 vssd1 vccd1 vccd1 _05596_/A sky130_fd_sc_hd__nand2_1
X_07332_ _07508_/A _07509_/A vssd1 vssd1 vccd1 vccd1 _07332_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_18_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07263_ _07263_/A _07263_/B vssd1 vssd1 vccd1 vccd1 _07265_/A sky130_fd_sc_hd__nand2_1
X_09002_ _09002_/A _09002_/B vssd1 vssd1 vccd1 vccd1 _09003_/A sky130_fd_sc_hd__nand2_1
X_07194_ _07201_/B _07201_/A vssd1 vssd1 vccd1 vccd1 _07195_/B sky130_fd_sc_hd__nand2_1
X_06214_ _06567_/C _06382_/A vssd1 vssd1 vccd1 vccd1 _06217_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06145_ _06250_/A _06145_/B vssd1 vssd1 vccd1 vccd1 _06145_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__08740__B _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06076_ _06891_/A _06082_/C vssd1 vssd1 vccd1 vccd1 _06081_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09904_ _09904_/A _09904_/B vssd1 vssd1 vccd1 vccd1 _09907_/B sky130_fd_sc_hd__nor2_1
X_09835_ _09835_/A _09835_/B vssd1 vssd1 vccd1 vccd1 _10090_/B sky130_fd_sc_hd__and2_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _09766_/A _09766_/B vssd1 vssd1 vccd1 vccd1 _09768_/B sky130_fd_sc_hd__nand2_1
X_06978_ _07138_/B _07138_/C vssd1 vssd1 vccd1 vccd1 _07137_/A sky130_fd_sc_hd__nand2_1
X_08717_ _08725_/A vssd1 vssd1 vccd1 vccd1 _10248_/B sky130_fd_sc_hd__inv_2
X_09697_ _10211_/B _10201_/B vssd1 vssd1 vccd1 vccd1 _09703_/B sky130_fd_sc_hd__nand2_1
X_05929_ _06755_/B _05929_/B _05929_/C vssd1 vssd1 vccd1 vccd1 _06755_/A sky130_fd_sc_hd__nand3_1
X_08648_ _09201_/A _10006_/A _08648_/C vssd1 vssd1 vccd1 vccd1 _08651_/A sky130_fd_sc_hd__nor3_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08579_ _08579_/A _08579_/B vssd1 vssd1 vccd1 vccd1 _08581_/B sky130_fd_sc_hd__nand2_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ hold20/X _10611_/A vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__nor2_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06716__A _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10541_ _10541_/A _10541_/B vssd1 vssd1 vccd1 vccd1 _10664_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_24_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10472_ _10479_/A _10472_/B _10472_/C vssd1 vssd1 vccd1 vccd1 _10476_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_32_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08097__B _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05514__B _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10739_ _10741_/CLK hold3/X fanout98/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10148__A _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07950_ _07950_/A _07950_/B vssd1 vssd1 vccd1 vccd1 _07952_/A sky130_fd_sc_hd__nand2_1
X_06901_ _06902_/B _06902_/A vssd1 vssd1 vccd1 vccd1 _06901_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_10_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07881_ _08724_/A input33/X vssd1 vssd1 vccd1 vccd1 _07884_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06832_ _09710_/B _10187_/B vssd1 vssd1 vccd1 vccd1 _06833_/B sky130_fd_sc_hd__nand2_1
X_09620_ _09620_/A _09620_/B vssd1 vssd1 vccd1 vccd1 _09664_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09551_ _10276_/A _10276_/C _09551_/C _09782_/B vssd1 vssd1 vccd1 vccd1 _09786_/B
+ sky130_fd_sc_hd__or4_2
X_06763_ _06763_/A _08819_/B _06763_/C vssd1 vssd1 vccd1 vccd1 _08819_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05714_ _05716_/C vssd1 vssd1 vccd1 vccd1 _05714_/Y sky130_fd_sc_hd__inv_2
XANTENNA__05424__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08502_ _08571_/A _08506_/C vssd1 vssd1 vccd1 vccd1 _08505_/A sky130_fd_sc_hd__nand2_1
X_09482_ _09482_/A _09482_/B vssd1 vssd1 vccd1 vccd1 _09483_/B sky130_fd_sc_hd__nand2_1
X_06694_ _07264_/A _07263_/A _07263_/B vssd1 vssd1 vccd1 vccd1 _07274_/C sky130_fd_sc_hd__nand3_2
X_08433_ _08555_/B vssd1 vssd1 vccd1 vccd1 _08556_/A sky130_fd_sc_hd__inv_2
X_05645_ _05646_/A _05647_/A vssd1 vssd1 vccd1 vccd1 _05695_/B sky130_fd_sc_hd__nand2_1
X_05576_ _05576_/A vssd1 vssd1 vccd1 vccd1 _05577_/B sky130_fd_sc_hd__inv_2
X_08364_ _08365_/A _08376_/B _08366_/B vssd1 vssd1 vccd1 vccd1 _08367_/A sky130_fd_sc_hd__a21o_1
XANTENNA__06536__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07315_ _07315_/A _07315_/B _07315_/C vssd1 vssd1 vccd1 vccd1 _07500_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08295_ _08295_/A _08324_/B vssd1 vssd1 vccd1 vccd1 _08296_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07246_ _07246_/A _07246_/B vssd1 vssd1 vccd1 vccd1 _07293_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07177_ _07350_/A _07349_/A vssd1 vssd1 vccd1 vccd1 _07182_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08470__B _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06271__A _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06128_ _08337_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _06281_/B sky130_fd_sc_hd__nand2_1
X_06059_ _06059_/A vssd1 vssd1 vccd1 vccd1 _06060_/A sky130_fd_sc_hd__inv_2
XANTENNA__07086__B _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09818_ _09818_/A _09818_/B vssd1 vssd1 vccd1 vccd1 _09824_/B sky130_fd_sc_hd__nand2_2
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09749_ input51/X _09749_/B vssd1 vssd1 vccd1 vccd1 _09752_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_68_102 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08645__B _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput18 a_i[25] vssd1 vssd1 vccd1 vccd1 input18/X sky130_fd_sc_hd__buf_2
X_10524_ _10525_/B _10525_/A vssd1 vssd1 vccd1 vccd1 _10526_/A sky130_fd_sc_hd__or2_1
Xinput29 a_i[6] vssd1 vssd1 vccd1 vccd1 input29/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__09476__B _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10455_ hold59/X vssd1 vssd1 vccd1 vccd1 _10456_/B sky130_fd_sc_hd__inv_2
XANTENNA__06181__A _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10386_ _10386_/A _10386_/B _10386_/C vssd1 vssd1 vccd1 vccd1 _10387_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_20_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10150__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09427__B1 _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05430_ _05430_/A _05430_/B vssd1 vssd1 vccd1 vccd1 _05437_/C sky130_fd_sc_hd__nand2_1
X_05361_ _05392_/A _05393_/B vssd1 vssd1 vccd1 vccd1 _05396_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_55_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07100_ _07243_/A _07106_/B _07100_/C vssd1 vssd1 vccd1 vccd1 _07106_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_70_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08080_ _08080_/A _08080_/B _08087_/B vssd1 vssd1 vccd1 vccd1 _08238_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_70_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09386__B _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07031_ _07032_/B _07032_/A vssd1 vssd1 vccd1 vccd1 _07031_/Y sky130_fd_sc_hd__nand2_1
X_08982_ _08988_/A _08988_/B vssd1 vssd1 vccd1 vccd1 _08987_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07933_ _07938_/B _07938_/A vssd1 vssd1 vccd1 vccd1 _08046_/B sky130_fd_sc_hd__nand2_1
X_07864_ _07864_/A vssd1 vssd1 vccd1 vccd1 _08387_/A sky130_fd_sc_hd__inv_2
X_09603_ _10151_/A _10150_/A _09922_/B _10148_/B vssd1 vssd1 vccd1 vccd1 _09604_/A
+ sky130_fd_sc_hd__and4_1
X_06815_ _08972_/B _06815_/B _06815_/C vssd1 vssd1 vccd1 vccd1 _09036_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07795_ _07795_/A _07796_/A vssd1 vssd1 vccd1 vccd1 _07798_/A sky130_fd_sc_hd__nand2_1
X_09534_ _09534_/A _09534_/B vssd1 vssd1 vccd1 vccd1 _09536_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06746_ _07785_/B vssd1 vssd1 vccd1 vccd1 _09971_/A sky130_fd_sc_hd__inv_2
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09465_ _09234_/A _09234_/B _09469_/B vssd1 vssd1 vccd1 vccd1 _09466_/B sky130_fd_sc_hd__o21a_1
X_06677_ _06679_/A _06679_/B vssd1 vssd1 vccd1 vccd1 _06678_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08416_ _08420_/A _08418_/A vssd1 vssd1 vccd1 vccd1 _08417_/C sky130_fd_sc_hd__nand2_1
X_05628_ _05632_/C vssd1 vssd1 vccd1 vccd1 _05629_/C sky130_fd_sc_hd__inv_2
XFILLER_0_80_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10028__B2 _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10028__A1 _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09418__B1 _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09396_ _09397_/A _09395_/Y vssd1 vssd1 vccd1 vccd1 _09611_/B sky130_fd_sc_hd__or2b_1
XFILLER_0_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05559_ _05559_/A vssd1 vssd1 vccd1 vccd1 _05560_/B sky130_fd_sc_hd__inv_2
X_08347_ _08347_/A _08347_/B vssd1 vssd1 vccd1 vccd1 _08349_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08481__A _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08278_ _08289_/B _08289_/C vssd1 vssd1 vccd1 vccd1 _08324_/A sky130_fd_sc_hd__nand2_1
X_07229_ _07229_/A _07229_/B vssd1 vssd1 vccd1 vccd1 _07230_/A sky130_fd_sc_hd__nand2_1
X_10240_ _10068_/A _10068_/B _10068_/C vssd1 vssd1 vccd1 vccd1 _10243_/A sky130_fd_sc_hd__a21boi_1
X_10171_ _10171_/A _10171_/B vssd1 vssd1 vccd1 vccd1 _10173_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05345__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09487__A _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__A _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10507_ _10507_/A _10653_/B vssd1 vssd1 vccd1 vccd1 _10508_/A sky130_fd_sc_hd__nand2_1
X_10438_ _10438_/A _10438_/B vssd1 vssd1 vccd1 vccd1 _10440_/A sky130_fd_sc_hd__nand2_1
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10369_ _10369_/A _10369_/B hold31/X vssd1 vssd1 vccd1 vccd1 _10558_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_79_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09648__B1 _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07580_ _07580_/A _07580_/B vssd1 vssd1 vccd1 vccd1 _07582_/A sky130_fd_sc_hd__nand2_1
X_06600_ _06600_/A _06600_/B _06600_/C vssd1 vssd1 vccd1 vccd1 _06943_/B sky130_fd_sc_hd__nand3_1
X_06531_ _07012_/C _06531_/B vssd1 vssd1 vccd1 vccd1 _06653_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_75_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09250_ _09250_/A _09250_/B vssd1 vssd1 vccd1 vccd1 _09278_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08201_ _08201_/A _08201_/B vssd1 vssd1 vccd1 vccd1 _08204_/C sky130_fd_sc_hd__nand2_1
X_06462_ _06608_/B _06608_/C _06461_/Y vssd1 vssd1 vccd1 vccd1 _06605_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09181_ _09181_/A _09181_/B _09409_/B vssd1 vssd1 vccd1 vccd1 _09409_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_50_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06393_ _06393_/A vssd1 vssd1 vccd1 vccd1 _06557_/B sky130_fd_sc_hd__inv_2
X_05413_ _05417_/A _05417_/C vssd1 vssd1 vccd1 vccd1 _05415_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_55_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08132_ _08146_/C vssd1 vssd1 vccd1 vccd1 _08155_/B sky130_fd_sc_hd__inv_2
XFILLER_0_7_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05344_ input10/X vssd1 vssd1 vccd1 vccd1 _10150_/B sky130_fd_sc_hd__buf_6
XFILLER_0_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08063_ _08225_/A vssd1 vssd1 vccd1 vccd1 _08064_/B sky130_fd_sc_hd__inv_2
XFILLER_0_3_452 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07014_ _10210_/B _10130_/A vssd1 vssd1 vccd1 vccd1 _07183_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_3_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08965_ _08967_/A _08967_/B vssd1 vssd1 vccd1 vccd1 _08966_/A sky130_fd_sc_hd__nand2_1
X_07916_ _07916_/A vssd1 vssd1 vccd1 vccd1 _07918_/A sky130_fd_sc_hd__inv_2
XFILLER_0_75_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08896_ _08946_/A vssd1 vssd1 vccd1 vccd1 _08945_/A sky130_fd_sc_hd__inv_2
X_07847_ _07850_/A _07847_/B vssd1 vssd1 vccd1 vccd1 _07849_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07778_ _07778_/A _07778_/B vssd1 vssd1 vccd1 vccd1 _07783_/A sky130_fd_sc_hd__nand2_1
X_09517_ input49/X input50/X _09517_/C _09517_/D vssd1 vssd1 vccd1 vccd1 _09518_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__10249__A1 input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10249__B2 _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06729_ _08478_/B _06732_/C vssd1 vssd1 vccd1 vccd1 _06731_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07380__A _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_38_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09448_ _09451_/B _09670_/A vssd1 vssd1 vccd1 vccd1 _09450_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09379_ _09379_/A _09641_/B _09379_/C vssd1 vssd1 vccd1 vccd1 _09641_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_19_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06443__B _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10223_ _10223_/A _10223_/B vssd1 vssd1 vccd1 vccd1 _10223_/Y sky130_fd_sc_hd__nor2_1
X_10154_ _10154_/A vssd1 vssd1 vccd1 vccd1 _10165_/B sky130_fd_sc_hd__inv_2
X_10085_ _10085_/A _10086_/A vssd1 vssd1 vccd1 vccd1 _10089_/A sky130_fd_sc_hd__nand2_1
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10156__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07465__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _08750_/A _08750_/B _08750_/C vssd1 vssd1 vccd1 vccd1 _08751_/B sky130_fd_sc_hd__nand3_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05962_ _05964_/B _05964_/C vssd1 vssd1 vccd1 vccd1 _06821_/B sky130_fd_sc_hd__nand2_1
X_08681_ _08681_/A _08681_/B vssd1 vssd1 vccd1 vccd1 _08692_/C sky130_fd_sc_hd__nand2_1
X_05893_ _05629_/B _05629_/C _05892_/Y vssd1 vssd1 vccd1 vccd1 _06902_/A sky130_fd_sc_hd__a21oi_2
X_07701_ _07701_/A _07701_/B _07701_/C vssd1 vssd1 vccd1 vccd1 _07702_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_45_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07632_ _09840_/B _10130_/A vssd1 vssd1 vccd1 vccd1 _07637_/A sky130_fd_sc_hd__nand2_1
X_09302_ _09302_/A _09302_/B vssd1 vssd1 vccd1 vccd1 _09309_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_48_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07563_ _07560_/Y _07607_/A _07562_/Y vssd1 vssd1 vccd1 vccd1 _07839_/B sky130_fd_sc_hd__a21oi_1
X_07494_ _07618_/B _07617_/A _07617_/B vssd1 vssd1 vccd1 vccd1 _07644_/C sky130_fd_sc_hd__nand3b_2
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06514_ _06638_/A _06639_/B vssd1 vssd1 vccd1 vccd1 _06642_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09233_ _09677_/A _09678_/C vssd1 vssd1 vccd1 vccd1 _09234_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_63_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06445_ _10112_/A _09677_/A vssd1 vssd1 vccd1 vccd1 _06622_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_28_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09164_ _10129_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _09165_/C sky130_fd_sc_hd__nand2_1
X_08115_ _08168_/B vssd1 vssd1 vccd1 vccd1 _08169_/B sky130_fd_sc_hd__inv_2
X_06376_ _06376_/A _06376_/B vssd1 vssd1 vccd1 vccd1 _06377_/A sky130_fd_sc_hd__nand2_1
X_09095_ _09096_/B _09096_/A vssd1 vssd1 vccd1 vccd1 _09539_/A sky130_fd_sc_hd__or2_1
XFILLER_0_71_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07359__B _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08046_ _08046_/A _08046_/B _08046_/C vssd1 vssd1 vccd1 vccd1 _08047_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09997_ _10001_/B _10001_/C vssd1 vssd1 vccd1 vccd1 _10000_/A sky130_fd_sc_hd__nand2_1
X_08948_ _08939_/B _08938_/C _08938_/B vssd1 vssd1 vccd1 vccd1 _08998_/A sky130_fd_sc_hd__a21o_1
XANTENNA__09590__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08879_ _08879_/A _08879_/B vssd1 vssd1 vccd1 vccd1 _08884_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_39_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08934__A input49/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09749__B _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10206_ _10206_/A _10206_/B vssd1 vssd1 vccd1 vccd1 _10209_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10137_ _10137_/A _10137_/B vssd1 vssd1 vccd1 vccd1 _10141_/B sky130_fd_sc_hd__nand2_1
X_10068_ _10068_/A _10068_/B _10068_/C vssd1 vssd1 vccd1 vccd1 _10073_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06230_ _06230_/A _06230_/B _06230_/C vssd1 vssd1 vccd1 vccd1 _06315_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_60_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06161_ _06161_/A _06161_/B vssd1 vssd1 vccd1 vccd1 _06162_/A sky130_fd_sc_hd__nand2_1
X_06092_ _05842_/A _05843_/A _05888_/A vssd1 vssd1 vccd1 vccd1 _06095_/A sky130_fd_sc_hd__o21a_1
X_09920_ _09921_/B _09921_/A vssd1 vssd1 vccd1 vccd1 _10170_/B sky130_fd_sc_hd__or2_1
XFILLER_0_40_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09851_ _10255_/A _09853_/B _09854_/B vssd1 vssd1 vccd1 vccd1 _09852_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _08802_/A _08802_/B _08802_/C vssd1 vssd1 vccd1 vccd1 _08803_/B sky130_fd_sc_hd__nand3_1
X_09782_ _09782_/A _09782_/B _09782_/C vssd1 vssd1 vccd1 vccd1 _09873_/A sky130_fd_sc_hd__or3_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06994_ _06994_/A _06994_/B _06996_/A vssd1 vssd1 vccd1 vccd1 _06999_/A sky130_fd_sc_hd__nand3_1
XANTENNA__05427__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08733_ _08734_/B _08734_/A vssd1 vssd1 vccd1 vccd1 _08748_/A sky130_fd_sc_hd__nor2_1
X_05945_ _05945_/A _05945_/B vssd1 vssd1 vccd1 vccd1 _05952_/A sky130_fd_sc_hd__nand2_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07923__A _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08664_ _08664_/A _08665_/A vssd1 vssd1 vccd1 vccd1 _08668_/A sky130_fd_sc_hd__nand2_1
X_05876_ _05876_/A _05876_/B vssd1 vssd1 vccd1 vccd1 _06199_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06539__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08595_ _08595_/A _08596_/A vssd1 vssd1 vccd1 vccd1 _08602_/B sky130_fd_sc_hd__nand2_1
X_07615_ _07615_/A _07615_/B _07615_/C vssd1 vssd1 vccd1 vccd1 _07616_/B sky130_fd_sc_hd__nand3_1
X_07546_ _07546_/A vssd1 vssd1 vccd1 vccd1 _07547_/C sky130_fd_sc_hd__inv_2
XFILLER_0_48_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _09216_/A _09216_/B vssd1 vssd1 vccd1 vccd1 _09217_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07477_ _07477_/A _07477_/B _07477_/C vssd1 vssd1 vccd1 vccd1 _07497_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_51_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06428_ _06428_/A _06428_/B _06428_/C vssd1 vssd1 vccd1 vccd1 _06602_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_44_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07089__B _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06359_ _06359_/A _06359_/B _06359_/C vssd1 vssd1 vccd1 vccd1 _06365_/B sky130_fd_sc_hd__nand3_1
X_09147_ _10103_/B _10128_/B vssd1 vssd1 vccd1 vccd1 _09393_/C sky130_fd_sc_hd__nand2_1
X_09078_ _09078_/A _10365_/C vssd1 vssd1 vccd1 vccd1 _09079_/A sky130_fd_sc_hd__nand2_1
X_08029_ _10292_/B _10158_/A vssd1 vssd1 vccd1 vccd1 _08052_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10722__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10686_ _10687_/B _10687_/A vssd1 vssd1 vccd1 vccd1 _10688_/A sky130_fd_sc_hd__or2_1
XFILLER_0_35_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06631__B _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05730_ _05731_/A _05731_/B vssd1 vssd1 vccd1 vccd1 _05730_/Y sky130_fd_sc_hd__nor2_1
X_05661_ _08453_/A _07891_/B vssd1 vssd1 vccd1 vccd1 _05664_/B sky130_fd_sc_hd__nand2_1
X_07400_ _07401_/B _07401_/A vssd1 vssd1 vccd1 vccd1 _07400_/Y sky130_fd_sc_hd__nand2_1
X_08380_ _10467_/A _10467_/B vssd1 vssd1 vccd1 vccd1 _10466_/A sky130_fd_sc_hd__nand2_1
X_05592_ _05592_/A _05592_/B vssd1 vssd1 vccd1 vccd1 _05598_/C sky130_fd_sc_hd__nand2_1
X_07331_ _07520_/C _07520_/B _07330_/Y vssd1 vssd1 vccd1 vccd1 _07509_/A sky130_fd_sc_hd__a21oi_4
XANTENNA__08574__A _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07262_ _07594_/A _07595_/A vssd1 vssd1 vccd1 vccd1 _07857_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_33_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09001_ _09001_/A _09002_/B _09002_/A vssd1 vssd1 vccd1 vccd1 _09018_/B sky130_fd_sc_hd__nand3_1
X_07193_ _07193_/A _07193_/B _07193_/C vssd1 vssd1 vccd1 vccd1 _07206_/B sky130_fd_sc_hd__nand3_1
X_06213_ _06382_/A _06382_/B _06383_/A vssd1 vssd1 vccd1 vccd1 _06567_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_26_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06144_ _06466_/C _06253_/B vssd1 vssd1 vccd1 vccd1 _06255_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_41_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06075_ _06075_/A _06075_/B _06075_/C vssd1 vssd1 vccd1 vccd1 _06082_/C sky130_fd_sc_hd__nand3_1
X_09903_ _09903_/A vssd1 vssd1 vccd1 vccd1 _09904_/B sky130_fd_sc_hd__inv_2
X_09834_ _10569_/A _10569_/B vssd1 vssd1 vccd1 vccd1 _10096_/A sky130_fd_sc_hd__nand2_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _09768_/C vssd1 vssd1 vccd1 vccd1 _09765_/Y sky130_fd_sc_hd__inv_2
X_06977_ _06977_/A _06977_/B _06977_/C vssd1 vssd1 vccd1 vccd1 _07138_/C sky130_fd_sc_hd__nand3_1
X_08716_ _08754_/A _08754_/C vssd1 vssd1 vccd1 vccd1 _08753_/A sky130_fd_sc_hd__nand2_1
X_09696_ _09722_/A _09722_/C vssd1 vssd1 vccd1 vccd1 _09721_/A sky130_fd_sc_hd__nand2_1
X_05928_ _05928_/A vssd1 vssd1 vccd1 vccd1 _05929_/C sky130_fd_sc_hd__inv_2
X_08647_ _10004_/A _10150_/A vssd1 vssd1 vccd1 vccd1 _08648_/C sky130_fd_sc_hd__nand2_1
X_05859_ _06113_/C _06113_/B vssd1 vssd1 vccd1 vccd1 _06115_/B sky130_fd_sc_hd__nand2_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05901__A input55/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ _08579_/B _08579_/A vssd1 vssd1 vccd1 vccd1 _09135_/A sky130_fd_sc_hd__or2_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07529_ _07666_/A _07667_/A vssd1 vssd1 vccd1 vccd1 _07659_/B sky130_fd_sc_hd__nand2_1
X_10540_ _10540_/A _10649_/A vssd1 vssd1 vccd1 vccd1 _10541_/B sky130_fd_sc_hd__nand2_1
X_10471_ _10471_/A _10471_/B vssd1 vssd1 vccd1 vccd1 _10476_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10738_ _10741_/CLK _10738_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__dfrtp_2
XFILLER_0_15_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10148__B _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10669_ _10669_/A hold44/X vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09953__A _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06900_ _09037_/A _06906_/C vssd1 vssd1 vccd1 vccd1 _09062_/B sky130_fd_sc_hd__nand2_1
X_07880_ _09517_/C input59/X vssd1 vssd1 vccd1 vccd1 _07883_/A sky130_fd_sc_hd__nand2_1
X_06831_ _08772_/B _06834_/C vssd1 vssd1 vccd1 vccd1 _06833_/A sky130_fd_sc_hd__nand2_1
X_09550_ input53/X vssd1 vssd1 vccd1 vccd1 _10276_/C sky130_fd_sc_hd__inv_2
X_06762_ _06762_/A _06762_/B vssd1 vssd1 vccd1 vccd1 _06764_/A sky130_fd_sc_hd__nand2_1
X_09481_ _09482_/B _09482_/A vssd1 vssd1 vccd1 vccd1 _09705_/A sky130_fd_sc_hd__or2_1
X_05713_ _05744_/B _05744_/C vssd1 vssd1 vccd1 vccd1 _05743_/A sky130_fd_sc_hd__nand2_1
X_08501_ _08501_/A _08501_/B vssd1 vssd1 vccd1 vccd1 _08506_/C sky130_fd_sc_hd__nand2_1
X_08432_ _08432_/A _08432_/B vssd1 vssd1 vccd1 vccd1 _08555_/B sky130_fd_sc_hd__nand2_1
X_06693_ _06692_/B _06693_/B _06693_/C vssd1 vssd1 vccd1 vccd1 _07263_/B sky130_fd_sc_hd__nand3b_1
X_05644_ _08337_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _05647_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05575_ _05575_/A _05576_/A vssd1 vssd1 vccd1 vccd1 _05578_/A sky130_fd_sc_hd__nand2_1
X_08363_ _08363_/A _08363_/B vssd1 vssd1 vccd1 vccd1 _08365_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05721__A _08725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08294_ _08294_/A _08321_/A vssd1 vssd1 vccd1 vccd1 _08295_/A sky130_fd_sc_hd__nand2_1
X_07314_ _07314_/A _07314_/B vssd1 vssd1 vccd1 vccd1 _07500_/B sky130_fd_sc_hd__nand2_1
X_07245_ _07246_/B _07246_/A vssd1 vssd1 vccd1 vccd1 _07429_/B sky130_fd_sc_hd__nor2_2
XFILLER_0_5_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07176_ _07350_/B vssd1 vssd1 vccd1 vccd1 _07349_/A sky130_fd_sc_hd__inv_2
XANTENNA__06271__B _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06127_ _08171_/B input5/X vssd1 vssd1 vccd1 vccd1 _06280_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06058_ _06058_/A _06059_/A vssd1 vssd1 vccd1 vccd1 _06071_/A sky130_fd_sc_hd__nand2_1
X_09817_ _09817_/A _09817_/B vssd1 vssd1 vccd1 vccd1 _09818_/B sky130_fd_sc_hd__nor2_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09748_ _09839_/B _09748_/B vssd1 vssd1 vccd1 vccd1 _09752_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09679_ _09679_/A vssd1 vssd1 vccd1 vccd1 _10003_/B sky130_fd_sc_hd__inv_2
XFILLER_0_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10523_ _10523_/A vssd1 vssd1 vccd1 vccd1 _10525_/B sky130_fd_sc_hd__inv_2
Xinput19 a_i[26] vssd1 vssd1 vccd1 vccd1 input19/X sky130_fd_sc_hd__buf_2
X_10454_ _10460_/A _10460_/C vssd1 vssd1 vccd1 vccd1 _10456_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10385_ _10385_/A _10385_/B vssd1 vssd1 vccd1 vccd1 _10390_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08389__A _08453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09427__A1 _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09427__B2 _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05360_ _08574_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _05393_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09386__C _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07468__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07030_ _07123_/A _07124_/A vssd1 vssd1 vccd1 vccd1 _07122_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_2_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08981_ _08995_/B _08981_/B vssd1 vssd1 vccd1 vccd1 _08988_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07932_ _07948_/C _07979_/B _07931_/Y vssd1 vssd1 vccd1 vccd1 _07938_/A sky130_fd_sc_hd__a21oi_1
X_07863_ _07863_/A _07863_/B vssd1 vssd1 vccd1 vccd1 _10386_/A sky130_fd_sc_hd__nor2_1
X_09602_ _10148_/A _09602_/B vssd1 vssd1 vccd1 vccd1 _09607_/A sky130_fd_sc_hd__nand2_1
X_06814_ _06818_/C vssd1 vssd1 vccd1 vccd1 _06815_/C sky130_fd_sc_hd__inv_2
X_09533_ _09537_/A _09766_/A vssd1 vssd1 vccd1 vccd1 _09771_/B sky130_fd_sc_hd__nand2_1
X_07794_ _07889_/C _07794_/B vssd1 vssd1 vccd1 vccd1 _07796_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06745_ _06744_/Y _10130_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _08435_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ _09467_/B _09692_/B vssd1 vssd1 vccd1 vccd1 _09466_/A sky130_fd_sc_hd__nand2_1
X_06676_ _06676_/A _06676_/B _06676_/C vssd1 vssd1 vccd1 vccd1 _06679_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_65_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08415_ _08418_/A _08420_/A vssd1 vssd1 vccd1 vccd1 _08660_/B sky130_fd_sc_hd__or2_1
XANTENNA__09418__A1 _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05627_ _05627_/A _05627_/B vssd1 vssd1 vccd1 vccd1 _05632_/C sky130_fd_sc_hd__nand2_1
X_09395_ _09397_/C _09397_/B vssd1 vssd1 vccd1 vccd1 _09395_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__05451__A _08453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10028__A2 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09418__B2 _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08346_ _08346_/A _08346_/B vssd1 vssd1 vccd1 vccd1 _08347_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05558_ _05558_/A _05559_/A vssd1 vssd1 vccd1 vccd1 _05564_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05489_ _05493_/A _05493_/C vssd1 vssd1 vccd1 vccd1 _05491_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08481__B _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08277_ _08277_/A _08277_/B vssd1 vssd1 vccd1 vccd1 _08289_/C sky130_fd_sc_hd__nand2_1
X_07228_ _07228_/A _07228_/B vssd1 vssd1 vccd1 vccd1 _07229_/A sky130_fd_sc_hd__nand2_1
X_07159_ _10103_/A _10004_/A vssd1 vssd1 vccd1 vccd1 _07187_/B sky130_fd_sc_hd__nand2_1
X_10170_ _10170_/A _10170_/B vssd1 vssd1 vccd1 vccd1 _10171_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08002__A _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05345__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08672__A _08672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09487__B _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08391__B _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10506_ _10506_/A _10506_/B vssd1 vssd1 vccd1 vccd1 _10507_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06192__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10437_ _10675_/B _10676_/A _10443_/B vssd1 vssd1 vccd1 vccd1 _10464_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__09593__B1 _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _10368_/A _10368_/B vssd1 vssd1 vccd1 vccd1 _10558_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _10303_/B _10303_/C vssd1 vssd1 vccd1 vccd1 _10301_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_18_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09648__B2 _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09648__A1 _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06530_ _06531_/B _06530_/B _06530_/C vssd1 vssd1 vccd1 vccd1 _07012_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_34_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08285__C _08363_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06461_ _06616_/A _06615_/A vssd1 vssd1 vccd1 vccd1 _06461_/Y sky130_fd_sc_hd__nor2_1
X_08200_ _08200_/A _08200_/B vssd1 vssd1 vccd1 vccd1 _08201_/B sky130_fd_sc_hd__nand2_1
X_05412_ _05439_/A _05439_/B vssd1 vssd1 vccd1 vccd1 _05417_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09678__A _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09180_ _09180_/A vssd1 vssd1 vccd1 vccd1 _09181_/B sky130_fd_sc_hd__inv_2
X_06392_ _08112_/A _10148_/A vssd1 vssd1 vccd1 vccd1 _06393_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08131_ _08133_/B _08133_/A vssd1 vssd1 vccd1 vccd1 _08146_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05343_ input55/X vssd1 vssd1 vccd1 vccd1 _08573_/A sky130_fd_sc_hd__buf_6
XFILLER_0_50_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08062_ _08218_/A _08217_/A _08217_/B vssd1 vssd1 vccd1 vccd1 _08225_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_3_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07013_ _07025_/B _07025_/C vssd1 vssd1 vccd1 vccd1 _07024_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07926__A _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08964_ _08964_/A _08964_/B _08964_/C vssd1 vssd1 vccd1 vccd1 _08967_/B sky130_fd_sc_hd__nand3_1
X_07915_ _07980_/B vssd1 vssd1 vccd1 vccd1 _07948_/C sky130_fd_sc_hd__inv_2
XFILLER_0_75_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08895_ _08893_/Y _08864_/B _08894_/Y vssd1 vssd1 vccd1 vccd1 _08946_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07846_ _07848_/A _07848_/C vssd1 vssd1 vccd1 vccd1 _07850_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07777_ _07777_/A _07777_/B vssd1 vssd1 vccd1 vccd1 _07778_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09516_ _09269_/Y _09271_/A _09270_/A vssd1 vssd1 vccd1 vccd1 _09528_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__10249__A2 _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07380__B _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06728_ _06728_/A _06728_/B vssd1 vssd1 vccd1 vccd1 _06732_/C sky130_fd_sc_hd__nand2_1
X_09447_ _09447_/A _09447_/B _09670_/B vssd1 vssd1 vccd1 vccd1 _09670_/A sky130_fd_sc_hd__nand3_1
X_06659_ _06659_/A _06659_/B _06659_/C vssd1 vssd1 vccd1 vccd1 _06665_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09378_ _09379_/A _09641_/B _09379_/C vssd1 vssd1 vccd1 vccd1 _09383_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_74_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08329_ _08329_/A _08329_/B vssd1 vssd1 vccd1 vccd1 _08360_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09100__B _09875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10222_ _10223_/B _10223_/A vssd1 vssd1 vccd1 vccd1 _10222_/Y sky130_fd_sc_hd__nand2_1
X_10153_ _10153_/A _10153_/B vssd1 vssd1 vccd1 vccd1 _10154_/A sky130_fd_sc_hd__xor2_1
X_10084_ _10084_/A _10084_/B vssd1 vssd1 vccd1 vccd1 _10086_/A sky130_fd_sc_hd__nor2_1
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_312 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10156__B _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07746__A _10247_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07465__B _07785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05961_ _05961_/A _05961_/B _05961_/C vssd1 vssd1 vccd1 vccd1 _05964_/C sky130_fd_sc_hd__nand3_1
X_07700_ _07638_/B _07777_/B _07777_/A vssd1 vssd1 vccd1 vccd1 _07701_/C sky130_fd_sc_hd__a21boi_1
X_08680_ _08692_/A _08694_/A vssd1 vssd1 vccd1 vccd1 _08683_/A sky130_fd_sc_hd__nand2_1
X_05892_ _05892_/A _05892_/B vssd1 vssd1 vccd1 vccd1 _05892_/Y sky130_fd_sc_hd__nor2_1
X_07631_ _07696_/A _07697_/A vssd1 vssd1 vccd1 vccd1 _07631_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07562_ _07604_/A _07603_/A vssd1 vssd1 vccd1 vccd1 _07562_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_0_10 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09301_ _09572_/B _09301_/B vssd1 vssd1 vccd1 vccd1 _09302_/A sky130_fd_sc_hd__nand2_1
X_06513_ _10103_/A _09602_/B vssd1 vssd1 vccd1 vccd1 _06639_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07493_ _07493_/A _07493_/B _07493_/C vssd1 vssd1 vccd1 vccd1 _07617_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_75_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09232_ _10201_/A _10005_/A vssd1 vssd1 vccd1 vccd1 _09234_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06444_ _08574_/A vssd1 vssd1 vccd1 vccd1 _10112_/A sky130_fd_sc_hd__buf_6
XANTENNA__09201__A _09201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09163_ _10157_/B vssd1 vssd1 vccd1 vccd1 _09912_/B sky130_fd_sc_hd__inv_2
X_06375_ _06346_/Y _06480_/B _06374_/Y vssd1 vssd1 vccd1 vccd1 _06380_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08114_ _09840_/B _08114_/B vssd1 vssd1 vccd1 vccd1 _08168_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09094_ _09094_/A _09094_/B vssd1 vssd1 vccd1 vccd1 _09096_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_9_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08045_ _08045_/A _08045_/B vssd1 vssd1 vccd1 vccd1 _08047_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09996_ _09996_/A _09996_/B vssd1 vssd1 vccd1 vccd1 _10001_/C sky130_fd_sc_hd__nand2_1
X_08947_ _09080_/B _08955_/C vssd1 vssd1 vccd1 vccd1 _08954_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09590__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _08878_/A _08878_/B vssd1 vssd1 vccd1 vccd1 _08879_/A sky130_fd_sc_hd__nand2_1
X_07829_ _07821_/C _07824_/A _07711_/Y vssd1 vssd1 vccd1 vccd1 _07830_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__07391__A _09551_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_204 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08934__B _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_470 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10205_ _10205_/A _10205_/B vssd1 vssd1 vccd1 vccd1 _10209_/B sky130_fd_sc_hd__xnor2_1
X_10136_ _10136_/A _10136_/B vssd1 vssd1 vccd1 vccd1 _10137_/B sky130_fd_sc_hd__nand2_1
X_10067_ _10067_/A vssd1 vssd1 vccd1 vccd1 _10068_/B sky130_fd_sc_hd__inv_2
XANTENNA__08397__A input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_2_3__f_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 _10741_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_212 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06160_ _06160_/A _06160_/B _06160_/C vssd1 vssd1 vccd1 vccd1 _06166_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_80_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06091_ _06091_/A _06091_/B vssd1 vssd1 vccd1 vccd1 _06095_/B sky130_fd_sc_hd__and2_1
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09850_ _09853_/A _09854_/C vssd1 vssd1 vccd1 vccd1 _09852_/B sky130_fd_sc_hd__nand2_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08801_ _08802_/A _08802_/B _08802_/C vssd1 vssd1 vccd1 vccd1 _08803_/A sky130_fd_sc_hd__a21o_1
X_09781_ _09873_/B _09781_/B vssd1 vssd1 vccd1 vccd1 _09782_/C sky130_fd_sc_hd__nand2_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _10211_/B _10101_/A vssd1 vssd1 vccd1 vccd1 _06996_/A sky130_fd_sc_hd__nand2_1
X_08732_ _08732_/A _09261_/A vssd1 vssd1 vccd1 vccd1 _08734_/A sky130_fd_sc_hd__nand2_1
X_05944_ _10128_/A _10187_/A vssd1 vssd1 vccd1 vccd1 _05945_/B sky130_fd_sc_hd__nand2_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07923__B _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08663_ _08663_/A _08663_/B vssd1 vssd1 vccd1 vccd1 _08665_/A sky130_fd_sc_hd__nand2_1
X_05875_ _05877_/B vssd1 vssd1 vccd1 vccd1 _05876_/B sky130_fd_sc_hd__inv_2
XANTENNA__06539__B input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08594_ _08594_/A _08594_/B vssd1 vssd1 vccd1 vccd1 _08596_/A sky130_fd_sc_hd__nand2_1
X_07614_ _07614_/A _07614_/B _07614_/C vssd1 vssd1 vccd1 vccd1 _07615_/B sky130_fd_sc_hd__nand3_1
X_07545_ _07545_/A _07545_/B _07545_/C vssd1 vssd1 vccd1 vccd1 _07547_/B sky130_fd_sc_hd__nand3_1
X_07476_ _07476_/A _07476_/B vssd1 vssd1 vccd1 vccd1 _07497_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_63_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09215_ _09218_/B _09218_/C vssd1 vssd1 vccd1 vccd1 _09217_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06427_ _06427_/A _06427_/B vssd1 vssd1 vccd1 vccd1 _06602_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09146_ _09154_/B _09381_/B vssd1 vssd1 vccd1 vccd1 _09153_/A sky130_fd_sc_hd__nand2_1
X_06358_ _06360_/A _06358_/B vssd1 vssd1 vccd1 vccd1 _06359_/B sky130_fd_sc_hd__nand2_1
X_09077_ _09351_/A _09077_/B _09077_/C vssd1 vssd1 vccd1 vccd1 _10365_/C sky130_fd_sc_hd__nand3_2
XFILLER_0_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06289_ _06424_/A _06425_/A vssd1 vssd1 vccd1 vccd1 _06289_/Y sky130_fd_sc_hd__nand2_1
X_08028_ _08037_/B _08037_/A vssd1 vssd1 vccd1 vccd1 _08148_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_189 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09979_ _09981_/B _09981_/A vssd1 vssd1 vccd1 vccd1 _09980_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_39_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10685_ _10685_/A _10685_/B vssd1 vssd1 vccd1 vccd1 _10687_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10119_ _10120_/B _10120_/A vssd1 vssd1 vccd1 vccd1 _10121_/A sky130_fd_sc_hd__or2_1
X_05660_ _05664_/A vssd1 vssd1 vccd1 vccd1 _05663_/A sky130_fd_sc_hd__inv_2
X_05591_ _05591_/A _05591_/B vssd1 vssd1 vccd1 vccd1 _05966_/B sky130_fd_sc_hd__nand2_1
X_07330_ _07516_/A _07517_/B vssd1 vssd1 vccd1 vccd1 _07330_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_42_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09000_ _09000_/A _09006_/A vssd1 vssd1 vccd1 vccd1 _09002_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07261_ _07583_/B _07583_/A vssd1 vssd1 vccd1 vccd1 _07595_/A sky130_fd_sc_hd__nor2_1
XANTENNA__08590__A _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07192_ _07195_/C _07192_/B _07192_/C vssd1 vssd1 vccd1 vccd1 _07196_/A sky130_fd_sc_hd__nand3b_1
X_06212_ _06388_/B _06386_/A vssd1 vssd1 vccd1 vccd1 _06383_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06143_ _06253_/B _06143_/B _06143_/C vssd1 vssd1 vccd1 vccd1 _06466_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_41_476 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05719__A _07756_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06074_ _06074_/A _06074_/B vssd1 vssd1 vccd1 vccd1 _06891_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09902_ _09902_/A _09902_/B vssd1 vssd1 vccd1 vccd1 _09904_/A sky130_fd_sc_hd__nor2_1
X_09833_ _09833_/A _09833_/B vssd1 vssd1 vccd1 vccd1 _10569_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ _09764_/A _09764_/B vssd1 vssd1 vccd1 vccd1 _09768_/C sky130_fd_sc_hd__nand2_1
X_06976_ _06976_/A _06976_/B vssd1 vssd1 vccd1 vccd1 _06977_/A sky130_fd_sc_hd__nand2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08715_ _08715_/A _09287_/A vssd1 vssd1 vccd1 vccd1 _08754_/C sky130_fd_sc_hd__nand2_1
X_09695_ _10059_/A _09695_/B vssd1 vssd1 vccd1 vccd1 _09722_/C sky130_fd_sc_hd__nand2_1
X_05927_ _05927_/A _05928_/A vssd1 vssd1 vccd1 vccd1 _05930_/A sky130_fd_sc_hd__nand2_1
X_08646_ _10187_/A vssd1 vssd1 vccd1 vccd1 _10006_/A sky130_fd_sc_hd__inv_2
X_05858_ _05858_/A _05858_/B vssd1 vssd1 vccd1 vccd1 _06113_/B sky130_fd_sc_hd__nand2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05789_ _05789_/A _05789_/B vssd1 vssd1 vccd1 vccd1 _05796_/A sky130_fd_sc_hd__nand2_1
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _09135_/B _08577_/B vssd1 vssd1 vccd1 vccd1 _08579_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07528_ _07682_/C _07674_/B _07527_/Y vssd1 vssd1 vccd1 vccd1 _07667_/A sky130_fd_sc_hd__a21oi_2
XANTENNA__05901__B _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07459_ _07534_/B vssd1 vssd1 vccd1 vccd1 _07535_/B sky130_fd_sc_hd__inv_2
XFILLER_0_17_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10470_ _10472_/B vssd1 vssd1 vccd1 vccd1 _10471_/B sky130_fd_sc_hd__inv_2
XFILLER_0_17_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09129_ _09129_/A vssd1 vssd1 vccd1 vccd1 _09130_/C sky130_fd_sc_hd__inv_2
XFILLER_0_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10737_ _10741_/CLK hold14/X fanout98/X vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10668_ _10668_/A _10668_/B vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10599_ _10630_/A hold49/X vssd1 vssd1 vccd1 vccd1 _10600_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05539__A _08672_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07754__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06830_ _06830_/A _06830_/B vssd1 vssd1 vccd1 vccd1 _06834_/C sky130_fd_sc_hd__nand2_1
X_06761_ _06763_/C vssd1 vssd1 vccd1 vccd1 _06762_/B sky130_fd_sc_hd__inv_2
X_09480_ _09705_/B _09480_/B vssd1 vssd1 vccd1 vccd1 _09482_/A sky130_fd_sc_hd__nand2_1
X_05712_ _05839_/A _05712_/B _05712_/C vssd1 vssd1 vccd1 vccd1 _05744_/C sky130_fd_sc_hd__nand3_1
X_06692_ _06692_/A _06692_/B vssd1 vssd1 vccd1 vccd1 _07263_/A sky130_fd_sc_hd__nand2_1
X_08500_ _08501_/B _08501_/A vssd1 vssd1 vccd1 vccd1 _08571_/A sky130_fd_sc_hd__or2_1
X_08431_ _08556_/B _08556_/C vssd1 vssd1 vccd1 vccd1 _08555_/A sky130_fd_sc_hd__nand2_1
X_05643_ _08171_/B input6/X vssd1 vssd1 vccd1 vccd1 _05646_/A sky130_fd_sc_hd__nand2_1
X_05574_ _07675_/A input38/X vssd1 vssd1 vccd1 vccd1 _05576_/A sky130_fd_sc_hd__nand2_1
X_08362_ _08362_/A _08362_/B vssd1 vssd1 vccd1 vccd1 _08363_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05721__B input35/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08293_ _08293_/A vssd1 vssd1 vccd1 vccd1 _08321_/A sky130_fd_sc_hd__inv_2
X_07313_ _07315_/A _07315_/B vssd1 vssd1 vccd1 vccd1 _07314_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_131 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07244_ _07207_/A _07204_/A _07237_/A vssd1 vssd1 vccd1 vccd1 _07246_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_82_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07175_ _09710_/B _10129_/A vssd1 vssd1 vccd1 vccd1 _07350_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_41_284 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06126_ _06251_/C _06251_/B vssd1 vssd1 vccd1 vccd1 _06145_/B sky130_fd_sc_hd__nand2_1
X_06057_ _06057_/A _06057_/B vssd1 vssd1 vccd1 vccd1 _06059_/A sky130_fd_sc_hd__nand2_1
X_09816_ _09816_/A vssd1 vssd1 vccd1 vccd1 _09817_/B sky130_fd_sc_hd__inv_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09747_ input49/X _10247_/B input50/X _09840_/B vssd1 vssd1 vccd1 vccd1 _09748_/B
+ sky130_fd_sc_hd__a22o_1
X_06959_ _06967_/B _06968_/C _06968_/B vssd1 vssd1 vccd1 vccd1 _06961_/B sky130_fd_sc_hd__nand3_1
X_09678_ _10004_/A _10187_/A _09678_/C _10005_/A vssd1 vssd1 vccd1 vccd1 _09679_/A
+ sky130_fd_sc_hd__and4_1
XANTENNA__08495__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08629_ _08630_/B _08630_/A vssd1 vssd1 vccd1 vccd1 _08629_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_49_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10522_ _10532_/B _10522_/B vssd1 vssd1 vccd1 vccd1 _10523_/A sky130_fd_sc_hd__nand2_1
X_10453_ _10542_/B _10453_/B _10453_/C vssd1 vssd1 vccd1 vccd1 _10460_/C sky130_fd_sc_hd__nand3_1
XANTENNA__10203__B1 _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10384_ _10384_/A _10384_/B vssd1 vssd1 vccd1 vccd1 _10596_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08389__B _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09675__A2 _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05822__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09427__A2 _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07749__A _08725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09386__D _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07468__B _07897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08980_ _08980_/A _08980_/B vssd1 vssd1 vccd1 vccd1 _08995_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_48_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07484__A input12/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07931_ _07930_/A _07930_/B _07930_/C vssd1 vssd1 vccd1 vccd1 _07931_/Y sky130_fd_sc_hd__a21oi_1
X_07862_ _10426_/C _07864_/A vssd1 vssd1 vccd1 vccd1 _07863_/B sky130_fd_sc_hd__nor2_1
X_09601_ _09936_/B _09609_/C vssd1 vssd1 vccd1 vccd1 _09608_/A sky130_fd_sc_hd__nand2_1
X_06813_ _08976_/A _06813_/B vssd1 vssd1 vccd1 vccd1 _06818_/C sky130_fd_sc_hd__nand2_1
X_09532_ _09766_/B _09532_/B _09532_/C vssd1 vssd1 vccd1 vccd1 _09766_/A sky130_fd_sc_hd__nand3_1
X_07793_ _07794_/B _07793_/B _07793_/C vssd1 vssd1 vccd1 vccd1 _07889_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06828__A _10210_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06744_ _10129_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _06744_/Y sky130_fd_sc_hd__nand2_1
X_09463_ _09463_/A _09463_/B _09463_/C vssd1 vssd1 vccd1 vccd1 _09692_/B sky130_fd_sc_hd__nand3_1
X_06675_ _06675_/A _06675_/B vssd1 vssd1 vccd1 vccd1 _06679_/A sky130_fd_sc_hd__nand2_1
X_08414_ _08414_/A _08414_/B vssd1 vssd1 vccd1 vccd1 _08420_/A sky130_fd_sc_hd__nand2_1
X_05626_ _05626_/A _05626_/B vssd1 vssd1 vccd1 vccd1 _05627_/B sky130_fd_sc_hd__nand2_1
X_09394_ _09394_/A vssd1 vssd1 vccd1 vccd1 _09397_/B sky130_fd_sc_hd__inv_2
XFILLER_0_80_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09418__A2 _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05557_ _07756_/A _10156_/A vssd1 vssd1 vccd1 vccd1 _05559_/A sky130_fd_sc_hd__nand2_1
X_08345_ _08345_/A _08345_/B vssd1 vssd1 vccd1 vccd1 _08346_/A sky130_fd_sc_hd__or2_1
XFILLER_0_80_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05488_ _05948_/A _05948_/B vssd1 vssd1 vccd1 vccd1 _05493_/C sky130_fd_sc_hd__nand2_1
X_08276_ _08276_/A _08276_/B _08276_/C vssd1 vssd1 vccd1 vccd1 _08289_/B sky130_fd_sc_hd__nand3_1
X_07227_ _07398_/A _07398_/C vssd1 vssd1 vccd1 vccd1 _07232_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_6_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07158_ _07187_/A vssd1 vssd1 vccd1 vccd1 _07161_/A sky130_fd_sc_hd__inv_2
X_06109_ _06111_/A _06111_/B vssd1 vssd1 vccd1 vccd1 _06110_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_14_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07089_ _10275_/B _10151_/A vssd1 vssd1 vccd1 vccd1 _07091_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08002__B _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10505_ hold46/X vssd1 vssd1 vccd1 vccd1 _10506_/B sky130_fd_sc_hd__inv_2
XANTENNA__06192__B _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10436_ _10443_/A _10443_/B vssd1 vssd1 vccd1 vccd1 _10676_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09593__A1 _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09593__B2 _10151_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10367_ hold31/X vssd1 vssd1 vccd1 vccd1 _10368_/B sky130_fd_sc_hd__inv_2
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10298_ _10298_/A _10298_/B _10298_/C vssd1 vssd1 vccd1 vccd1 _10303_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_18_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06460_ _06617_/C vssd1 vssd1 vccd1 vccd1 _06608_/C sky130_fd_sc_hd__inv_2
XFILLER_0_68_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05411_ _05411_/A _05411_/B vssd1 vssd1 vccd1 vccd1 _05417_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09678__B _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08130_ _08130_/A _08130_/B vssd1 vssd1 vccd1 vccd1 _08133_/A sky130_fd_sc_hd__and2_1
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06391_ _06394_/A _06394_/B vssd1 vssd1 vccd1 vccd1 _06557_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07479__A _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05342_ _05476_/B vssd1 vssd1 vccd1 vccd1 _05353_/B sky130_fd_sc_hd__inv_2
XFILLER_0_70_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08061_ _08061_/A _08061_/B _08061_/C vssd1 vssd1 vccd1 vccd1 _08217_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_31_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07012_ _07032_/A _07012_/B _07012_/C vssd1 vssd1 vccd1 vccd1 _07025_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07926__B _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ _08963_/A _08963_/B vssd1 vssd1 vccd1 vccd1 _08967_/A sky130_fd_sc_hd__nand2_1
X_07914_ _07914_/A _07914_/B vssd1 vssd1 vccd1 vccd1 _07980_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08894_ _08894_/A _08894_/B vssd1 vssd1 vccd1 vccd1 _08894_/Y sky130_fd_sc_hd__nor2_1
X_07845_ _08382_/B _08382_/A vssd1 vssd1 vccd1 vccd1 _08381_/A sky130_fd_sc_hd__nor2_1
X_07776_ _07776_/A _07776_/B vssd1 vssd1 vccd1 vccd1 _07943_/B sky130_fd_sc_hd__nand2_2
X_09515_ _09570_/B _09810_/B vssd1 vssd1 vccd1 vccd1 _09568_/A sky130_fd_sc_hd__nand2_1
X_06727_ _06728_/A _06728_/B vssd1 vssd1 vccd1 vccd1 _08478_/B sky130_fd_sc_hd__or2_1
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09446_ _09446_/A vssd1 vssd1 vccd1 vccd1 _09447_/A sky130_fd_sc_hd__inv_2
X_06658_ _06953_/A _06954_/A vssd1 vssd1 vccd1 vccd1 _06952_/C sky130_fd_sc_hd__nand2_1
X_05609_ _05611_/A _05611_/B vssd1 vssd1 vccd1 vccd1 _05610_/A sky130_fd_sc_hd__nor2_1
X_09377_ _09377_/A vssd1 vssd1 vccd1 vccd1 _09379_/C sky130_fd_sc_hd__inv_2
X_06589_ _06589_/A _06589_/B vssd1 vssd1 vccd1 vccd1 _07060_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07389__A input36/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08328_ _08330_/A vssd1 vssd1 vccd1 vccd1 _08329_/B sky130_fd_sc_hd__inv_2
XFILLER_0_61_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08259_ _10284_/B _10292_/B _10112_/A _10108_/B vssd1 vssd1 vccd1 vccd1 _08304_/B
+ sky130_fd_sc_hd__and4_1
XANTENNA__10716__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10221_ _10227_/A _10227_/B vssd1 vssd1 vccd1 vccd1 _10226_/A sky130_fd_sc_hd__nand2_1
X_10152_ _10152_/A _10152_/B vssd1 vssd1 vccd1 vccd1 _10153_/B sky130_fd_sc_hd__xnor2_1
X_10083_ _10083_/A vssd1 vssd1 vccd1 vccd1 _10084_/B sky130_fd_sc_hd__inv_2
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_298 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_424 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07746__B _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10419_ _10419_/A hold62/X _10419_/C vssd1 vssd1 vccd1 vccd1 _10681_/B sky130_fd_sc_hd__nand3_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_87 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05960_ _05960_/A _05960_/B vssd1 vssd1 vccd1 vccd1 _05964_/B sky130_fd_sc_hd__nand2_1
X_05891_ _05749_/Y _06110_/B _05890_/Y vssd1 vssd1 vccd1 vccd1 _06102_/B sky130_fd_sc_hd__a21o_1
X_07630_ _07687_/C _07686_/B _07684_/A vssd1 vssd1 vccd1 vccd1 _07697_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_45_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07561_ _07561_/A _07561_/B vssd1 vssd1 vccd1 vccd1 _07607_/A sky130_fd_sc_hd__nor2_1
X_09300_ _09300_/A _09572_/B _09301_/B vssd1 vssd1 vccd1 vccd1 _09572_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_0_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06512_ _08337_/A vssd1 vssd1 vccd1 vccd1 _10103_/A sky130_fd_sc_hd__buf_6
XFILLER_0_48_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07492_ _07492_/A vssd1 vssd1 vccd1 vccd1 _07493_/C sky130_fd_sc_hd__inv_2
X_09231_ _09231_/A vssd1 vssd1 vccd1 vccd1 _09236_/B sky130_fd_sc_hd__inv_2
XFILLER_0_0_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06443_ _10108_/B _10004_/A vssd1 vssd1 vccd1 vccd1 _06621_/A sky130_fd_sc_hd__nand2_1
X_09162_ _09162_/A vssd1 vssd1 vccd1 vccd1 _09169_/B sky130_fd_sc_hd__inv_2
XFILLER_0_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06374_ _06477_/A _06476_/A vssd1 vssd1 vccd1 vccd1 _06374_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_43_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08113_ _08164_/A _08165_/A vssd1 vssd1 vccd1 vccd1 _08167_/B sky130_fd_sc_hd__nand2_1
X_09093_ input49/X _09749_/B vssd1 vssd1 vccd1 vccd1 _09094_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_31_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08044_ _08142_/C _08141_/B _08026_/Y vssd1 vssd1 vccd1 vccd1 _08048_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_3_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09995_ _09995_/A _09995_/B vssd1 vssd1 vccd1 vccd1 _09996_/A sky130_fd_sc_hd__nand2_1
X_08946_ _08946_/A _08946_/B vssd1 vssd1 vccd1 vccd1 _08955_/C sky130_fd_sc_hd__nand2_1
X_08877_ _08970_/B vssd1 vssd1 vccd1 vccd1 _08961_/A sky130_fd_sc_hd__inv_2
X_07828_ _07828_/A _07828_/B vssd1 vssd1 vccd1 vccd1 _07830_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07391__B _09201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ _07759_/A _07759_/B vssd1 vssd1 vccd1 vccd1 _07764_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_39_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09429_ _10187_/A _10148_/A vssd1 vssd1 vccd1 vccd1 _09431_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10204_ _10204_/A _10204_/B vssd1 vssd1 vccd1 vccd1 _10205_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10135_ _10136_/B _10136_/A vssd1 vssd1 vccd1 vccd1 _10137_/A sky130_fd_sc_hd__or2_1
X_10066_ _10066_/A _10067_/A vssd1 vssd1 vccd1 vccd1 _10073_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05830__A input46/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06090_ _06102_/B _06103_/B _06103_/C vssd1 vssd1 vccd1 vccd1 _06101_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_40_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08800_ _08800_/A vssd1 vssd1 vccd1 vccd1 _08802_/C sky130_fd_sc_hd__inv_2
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ input52/X _10275_/B input53/X _10284_/B vssd1 vssd1 vccd1 vccd1 _09781_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ _06995_/A _07008_/B vssd1 vssd1 vccd1 vccd1 _06994_/B sky130_fd_sc_hd__nand2_1
X_08731_ _08729_/Y _09261_/B _08731_/C vssd1 vssd1 vccd1 vccd1 _09261_/A sky130_fd_sc_hd__nand3b_1
XFILLER_0_56_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05943_ _06760_/B _05946_/C vssd1 vssd1 vccd1 vccd1 _05945_/A sky130_fd_sc_hd__nand2_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08662_ _08661_/B _08662_/B _08662_/C vssd1 vssd1 vccd1 vccd1 _08663_/B sky130_fd_sc_hd__nand3b_1
X_05874_ _08112_/A input40/X vssd1 vssd1 vccd1 vccd1 _05877_/B sky130_fd_sc_hd__nand2_1
X_07613_ _07613_/A _07613_/B vssd1 vssd1 vccd1 vccd1 _07615_/A sky130_fd_sc_hd__nand2_1
X_08593_ _08587_/Y _08593_/B _08593_/C vssd1 vssd1 vccd1 vccd1 _08594_/B sky130_fd_sc_hd__nand3b_1
X_07544_ _07544_/A _07544_/B vssd1 vssd1 vccd1 vccd1 _07547_/A sky130_fd_sc_hd__nand2_1
X_07475_ _07477_/A vssd1 vssd1 vccd1 vccd1 _07476_/B sky130_fd_sc_hd__inv_2
XFILLER_0_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09214_ _09214_/A _09441_/A _09214_/C vssd1 vssd1 vccd1 vccd1 _09218_/C sky130_fd_sc_hd__nand3_1
X_06426_ _06428_/A _06428_/B vssd1 vssd1 vccd1 vccd1 _06427_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06357_ _06357_/A vssd1 vssd1 vccd1 vccd1 _06360_/A sky130_fd_sc_hd__inv_2
X_09145_ _09145_/A _09145_/B _09145_/C vssd1 vssd1 vccd1 vccd1 _09381_/B sky130_fd_sc_hd__nand3_1
X_09076_ _09076_/A _09076_/B vssd1 vssd1 vccd1 vccd1 _09078_/A sky130_fd_sc_hd__nand2_1
X_06288_ _06422_/B _06422_/C _06287_/Y vssd1 vssd1 vccd1 vccd1 _06425_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08027_ _08142_/C _08141_/B _08026_/Y vssd1 vssd1 vccd1 vccd1 _08037_/A sky130_fd_sc_hd__a21oi_1
X_09978_ _09636_/A _09636_/B _09635_/A vssd1 vssd1 vccd1 vccd1 _09981_/A sky130_fd_sc_hd__o21a_1
X_08929_ _08930_/B _08930_/A vssd1 vssd1 vccd1 vccd1 _08929_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06746__A _07785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10731__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10684_ _10684_/A _10678_/A vssd1 vssd1 vccd1 vccd1 _10685_/A sky130_fd_sc_hd__or2b_1
XFILLER_0_35_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10118_ _10118_/A _10118_/B vssd1 vssd1 vccd1 vccd1 _10120_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_26_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10049_ _10049_/A _10049_/B vssd1 vssd1 vccd1 vccd1 _10052_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05590_ _05592_/B vssd1 vssd1 vccd1 vccd1 _05591_/B sky130_fd_sc_hd__inv_2
XFILLER_0_42_32 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07260_ _07260_/A _07260_/B vssd1 vssd1 vccd1 vccd1 _07583_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_53_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07191_ _07201_/A _07193_/C _07193_/B vssd1 vssd1 vccd1 vccd1 _07192_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06211_ _06387_/B _06386_/A _06386_/B vssd1 vssd1 vccd1 vccd1 _06388_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__08590__B _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07487__A _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06142_ _06322_/B _06323_/B vssd1 vssd1 vccd1 vccd1 _06143_/C sky130_fd_sc_hd__nand2_1
X_06073_ _06075_/C vssd1 vssd1 vccd1 vccd1 _06074_/B sky130_fd_sc_hd__inv_2
X_09901_ _09907_/A _09907_/C vssd1 vssd1 vccd1 vccd1 _09906_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05719__B input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09832_ _10353_/C _10353_/B vssd1 vssd1 vccd1 vccd1 _09833_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_67_73 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _09764_/B _09764_/A vssd1 vssd1 vccd1 vccd1 _09763_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__05735__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08714_ _08714_/A _08714_/B vssd1 vssd1 vccd1 vccd1 _09287_/A sky130_fd_sc_hd__nand2_1
X_06975_ _06975_/A _06975_/B _06975_/C vssd1 vssd1 vccd1 vccd1 _07138_/B sky130_fd_sc_hd__nand3_1
XANTENNA__08111__A _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09694_ _10059_/A _10059_/B vssd1 vssd1 vccd1 vccd1 _09722_/A sky130_fd_sc_hd__nand2b_1
X_05926_ _08101_/B _10148_/B vssd1 vssd1 vccd1 vccd1 _05928_/A sky130_fd_sc_hd__nand2_1
X_08645_ _09677_/A _10148_/A vssd1 vssd1 vccd1 vccd1 _09237_/A sky130_fd_sc_hd__nand2_1
X_05857_ _05857_/A _05857_/B vssd1 vssd1 vccd1 vccd1 _05858_/A sky130_fd_sc_hd__nand2_1
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08576_ _08576_/A _08576_/B vssd1 vssd1 vccd1 vccd1 _08577_/B sky130_fd_sc_hd__nand2_1
X_05788_ _06040_/B _05788_/B vssd1 vssd1 vccd1 vccd1 _05789_/A sky130_fd_sc_hd__nand2_1
X_07527_ _07670_/A _07671_/A vssd1 vssd1 vccd1 vccd1 _07527_/Y sky130_fd_sc_hd__nor2_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07458_ _07675_/A _08101_/B vssd1 vssd1 vccd1 vccd1 _07534_/B sky130_fd_sc_hd__nand2_1
X_07389_ input36/X vssd1 vssd1 vccd1 vccd1 _09201_/A sky130_fd_sc_hd__clkinv_4
XFILLER_0_51_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06409_ _06409_/A _06409_/B vssd1 vssd1 vccd1 vccd1 _06411_/A sky130_fd_sc_hd__nand2_1
X_09128_ _09128_/A _09129_/A vssd1 vssd1 vccd1 vccd1 _09131_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09059_ _09058_/B _09059_/B _09059_/C vssd1 vssd1 vccd1 vccd1 _09328_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08021__A _09551_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10736_ _10741_/CLK hold22/X fanout98/X vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10667_ _10667_/A _10667_/B vssd1 vssd1 vccd1 vccd1 _10669_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10598_ hold49/X _10630_/A vssd1 vssd1 vccd1 vccd1 _10600_/A sky130_fd_sc_hd__or2_1
XANTENNA__05539__B input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07754__B _08171_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput90 hold4/A vssd1 vssd1 vccd1 vccd1 y_o[31] sky130_fd_sc_hd__buf_12
XFILLER_0_37_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06760_ _06760_/A _06760_/B vssd1 vssd1 vccd1 vccd1 _06763_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_77_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05711_ _05711_/A _05839_/B vssd1 vssd1 vccd1 vccd1 _05744_/B sky130_fd_sc_hd__nand2_1
X_06691_ _06693_/B _06693_/C vssd1 vssd1 vccd1 vccd1 _06692_/A sky130_fd_sc_hd__nand2_1
X_08430_ _08430_/A _08430_/B vssd1 vssd1 vccd1 vccd1 _08556_/C sky130_fd_sc_hd__nand2_1
X_05642_ _05696_/B vssd1 vssd1 vccd1 vccd1 _05654_/B sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_53_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08361_ _10517_/B _08361_/B vssd1 vssd1 vccd1 vccd1 _10511_/B sky130_fd_sc_hd__nand2_1
X_05573_ input29/X vssd1 vssd1 vccd1 vccd1 _07675_/A sky130_fd_sc_hd__buf_6
XFILLER_0_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09697__A _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07312_ _07312_/A _07312_/B _07312_/C vssd1 vssd1 vccd1 vccd1 _07315_/B sky130_fd_sc_hd__nand3_1
X_08292_ _08292_/A _08292_/B vssd1 vssd1 vccd1 vccd1 _08294_/A sky130_fd_sc_hd__nand2_1
X_07243_ _07243_/A _07243_/B vssd1 vssd1 vccd1 vccd1 _07246_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_143 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07174_ _07349_/B vssd1 vssd1 vccd1 vccd1 _07350_/A sky130_fd_sc_hd__inv_2
XFILLER_0_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06125_ _06125_/A _06125_/B vssd1 vssd1 vccd1 vccd1 _06251_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06056_ _06060_/B _06869_/A vssd1 vssd1 vccd1 vccd1 _06058_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09815_ _09815_/A _09815_/B vssd1 vssd1 vccd1 vccd1 _09817_/A sky130_fd_sc_hd__nor2_1
XANTENNA__05465__A _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09746_ _09746_/A vssd1 vssd1 vccd1 vccd1 _09839_/B sky130_fd_sc_hd__inv_2
X_06958_ _06977_/C _06977_/B _06633_/Y vssd1 vssd1 vccd1 vccd1 _06967_/B sky130_fd_sc_hd__a21o_1
X_09677_ _09677_/A _10187_/B vssd1 vssd1 vccd1 vccd1 _09683_/B sky130_fd_sc_hd__nand2_1
X_05909_ _05909_/A _05910_/A vssd1 vssd1 vccd1 vccd1 _05917_/A sky130_fd_sc_hd__nand2_1
X_08628_ _09134_/B _08666_/C vssd1 vssd1 vccd1 vccd1 _08664_/A sky130_fd_sc_hd__nand2_1
X_06889_ _06895_/A _06895_/B vssd1 vssd1 vccd1 vccd1 _06894_/A sky130_fd_sc_hd__nand2_1
X_08559_ _08558_/B _08559_/B _08559_/C vssd1 vssd1 vccd1 vccd1 _08560_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10521_ _10641_/A _10519_/Y _10641_/B vssd1 vssd1 vccd1 vccd1 _10644_/A sky130_fd_sc_hd__a21boi_1
XFILLER_0_64_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10203__A1 _09677_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10452_ _10452_/A vssd1 vssd1 vccd1 vccd1 _10453_/C sky130_fd_sc_hd__inv_2
XANTENNA__10203__B2 _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10383_ _10383_/A _10383_/B vssd1 vssd1 vccd1 vccd1 _10384_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_20_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05375__A _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__A _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09675__A3 _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05822__B _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10719_ _10724_/CLK hold45/X fanout99/X vssd1 vssd1 vccd1 vccd1 hold59/A sky130_fd_sc_hd__dfrtp_1
XANTENNA__07749__B _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07930_ _07930_/A _07930_/B _07930_/C vssd1 vssd1 vccd1 vccd1 _07979_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07484__B _07646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ _10406_/B _10409_/A _10403_/B vssd1 vssd1 vccd1 vccd1 _07864_/A sky130_fd_sc_hd__nand3_1
X_06812_ _06811_/B _06812_/B _06812_/C vssd1 vssd1 vccd1 vccd1 _06813_/B sky130_fd_sc_hd__nand3b_1
X_09600_ _09600_/A _09600_/B vssd1 vssd1 vccd1 vccd1 _09609_/C sky130_fd_sc_hd__nand2_1
X_07792_ _07792_/A _07792_/B vssd1 vssd1 vccd1 vccd1 _07793_/C sky130_fd_sc_hd__nand2_1
X_09531_ _09766_/B _09532_/C _09532_/B vssd1 vssd1 vccd1 vccd1 _09537_/A sky130_fd_sc_hd__a21o_1
XFILLER_0_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06743_ _06767_/A _06768_/A vssd1 vssd1 vccd1 vccd1 _06766_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06828__B _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ _09463_/A _09463_/B _09463_/C vssd1 vssd1 vccd1 vccd1 _09467_/B sky130_fd_sc_hd__a21o_1
X_06674_ _06676_/A vssd1 vssd1 vccd1 vccd1 _06675_/B sky130_fd_sc_hd__inv_2
XFILLER_0_65_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08413_ _08407_/Y _08413_/B _08413_/C vssd1 vssd1 vccd1 vccd1 _08414_/B sky130_fd_sc_hd__nand3b_1
X_05625_ _05625_/A _05625_/B vssd1 vssd1 vccd1 vccd1 _05626_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09393_ _09393_/A _09393_/B _09393_/C vssd1 vssd1 vccd1 vccd1 _09394_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_80_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05556_ input35/X vssd1 vssd1 vccd1 vccd1 _10156_/A sky130_fd_sc_hd__clkbuf_8
X_08344_ _08353_/B _08344_/B vssd1 vssd1 vccd1 vccd1 _08347_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_46_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_196 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05487_ _05487_/A _05487_/B vssd1 vssd1 vccd1 vccd1 _05493_/A sky130_fd_sc_hd__nand2_1
X_08275_ _08292_/B _08275_/B vssd1 vssd1 vccd1 vccd1 _08276_/A sky130_fd_sc_hd__nand2_1
X_07226_ _07233_/A _07226_/B _07226_/C vssd1 vssd1 vccd1 vccd1 _07398_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_14_230 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07157_ _10211_/B _10103_/B vssd1 vssd1 vccd1 vccd1 _07187_/A sky130_fd_sc_hd__nand2_1
X_06108_ _06108_/A _06108_/B vssd1 vssd1 vccd1 vccd1 _06111_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07675__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07088_ _09778_/D _10150_/A vssd1 vssd1 vccd1 vccd1 _07091_/A sky130_fd_sc_hd__nand2_1
X_06039_ _06042_/B _06042_/C vssd1 vssd1 vccd1 vccd1 _06041_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_10_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09729_ _10060_/A _09729_/B _09896_/A vssd1 vssd1 vccd1 vccd1 _09733_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_56_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10504_ _10504_/A _10504_/B vssd1 vssd1 vccd1 vccd1 _10506_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10435_ _10435_/A _10435_/B hold63/X vssd1 vssd1 vccd1 vccd1 _10443_/B sky130_fd_sc_hd__nand3_1
XANTENNA__09593__A2 _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10366_ _10369_/A _10369_/B vssd1 vssd1 vccd1 vccd1 _10368_/A sky130_fd_sc_hd__nand2_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ _10297_/A _10297_/B vssd1 vssd1 vccd1 vccd1 _10303_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05410_ _05439_/B vssd1 vssd1 vccd1 vccd1 _05411_/B sky130_fd_sc_hd__inv_2
XANTENNA__09678__C _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06390_ _09517_/C _10151_/A vssd1 vssd1 vccd1 vccd1 _06394_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_50_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07479__B _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05341_ _08574_/A _10148_/B vssd1 vssd1 vccd1 vccd1 _05476_/B sky130_fd_sc_hd__nand2_1
X_08060_ _08060_/A _08060_/B vssd1 vssd1 vccd1 vccd1 _08061_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_70_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07011_ _07032_/B _07011_/B vssd1 vssd1 vccd1 vccd1 _07025_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_51_380 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_74 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08962_ _09031_/B _08969_/B vssd1 vssd1 vccd1 vccd1 _08963_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08893_ _08894_/B _08894_/A vssd1 vssd1 vccd1 vccd1 _08893_/Y sky130_fd_sc_hd__nand2_1
X_07913_ _07913_/A _07913_/B _07913_/C vssd1 vssd1 vccd1 vccd1 _07914_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_75_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07844_ _07844_/A _07852_/A vssd1 vssd1 vccd1 vccd1 _08382_/A sky130_fd_sc_hd__nand2_1
X_07775_ _07775_/A _07775_/B vssd1 vssd1 vccd1 vccd1 _07776_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_78_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09514_ _09513_/B _09514_/B _09739_/A vssd1 vssd1 vccd1 vccd1 _09810_/B sky130_fd_sc_hd__nand3b_2
X_06726_ _10112_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _06728_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_66_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09445_ _09445_/A _09446_/A vssd1 vssd1 vccd1 vccd1 _09451_/B sky130_fd_sc_hd__nand2_1
X_06657_ _06647_/Y _06964_/B _06656_/Y vssd1 vssd1 vccd1 vccd1 _06954_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05608_ _07756_/A _10151_/A vssd1 vssd1 vccd1 vccd1 _05611_/B sky130_fd_sc_hd__nand2_1
X_09376_ _09376_/A _09376_/B vssd1 vssd1 vccd1 vccd1 _09377_/A sky130_fd_sc_hd__xor2_1
X_06588_ _06590_/B vssd1 vssd1 vccd1 vccd1 _06589_/B sky130_fd_sc_hd__inv_2
XFILLER_0_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_05539_ _08672_/A input64/X vssd1 vssd1 vccd1 vccd1 _05547_/A sky130_fd_sc_hd__nand2_1
X_08327_ _08359_/A _08326_/Y vssd1 vssd1 vccd1 vccd1 _08330_/A sky130_fd_sc_hd__nor2b_1
XFILLER_0_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08258_ _08304_/A vssd1 vssd1 vccd1 vccd1 _08258_/Y sky130_fd_sc_hd__inv_2
XFILLER_0_34_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07209_ _07212_/B vssd1 vssd1 vccd1 vccd1 _07214_/B sky130_fd_sc_hd__inv_2
X_10220_ _10220_/A _10220_/B _10220_/C vssd1 vssd1 vccd1 vccd1 _10227_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_61_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08189_ _08176_/Y _08177_/A _08175_/A vssd1 vssd1 vccd1 vccd1 _08192_/A sky130_fd_sc_hd__o21a_1
X_10151_ _10151_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _10152_/B sky130_fd_sc_hd__nand2_1
X_10082_ _10082_/A _10082_/B vssd1 vssd1 vccd1 vccd1 _10084_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_69_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10418_ _10682_/B vssd1 vssd1 vccd1 vccd1 _10418_/Y sky130_fd_sc_hd__inv_2
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ _10376_/A _10376_/B hold61/X vssd1 vssd1 vccd1 vccd1 _10705_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05890_ _06106_/A _06108_/A vssd1 vssd1 vccd1 vccd1 _05890_/Y sky130_fd_sc_hd__nor2_1
X_07560_ _07603_/A _07604_/A vssd1 vssd1 vccd1 vccd1 _07560_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_48_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06511_ _10201_/A _10103_/B vssd1 vssd1 vccd1 vccd1 _06638_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09230_ _10212_/B _10187_/B vssd1 vssd1 vccd1 vccd1 _09231_/A sky130_fd_sc_hd__nand2_1
X_07491_ _07491_/A _07492_/A vssd1 vssd1 vccd1 vccd1 _07617_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_75_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06442_ _08573_/A vssd1 vssd1 vccd1 vccd1 _10108_/B sky130_fd_sc_hd__buf_6
XFILLER_0_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09161_ _10128_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _09162_/A sky130_fd_sc_hd__nand2_1
X_06373_ _06365_/A _06364_/A _06659_/B vssd1 vssd1 vccd1 vccd1 _06480_/B sky130_fd_sc_hd__o21ai_1
X_09092_ input50/X _10275_/B vssd1 vssd1 vccd1 vccd1 _09094_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08112_ _08112_/A _08574_/A vssd1 vssd1 vccd1 vccd1 _08165_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08043_ _08043_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08051_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_16_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08114__A _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09994_ _09994_/A _09995_/A _09995_/B vssd1 vssd1 vccd1 vccd1 _10001_/B sky130_fd_sc_hd__nand3_1
X_08945_ _08945_/A _08945_/B vssd1 vssd1 vccd1 vccd1 _09080_/B sky130_fd_sc_hd__nand2_1
X_08876_ _08876_/A _08876_/B vssd1 vssd1 vccd1 vccd1 _08970_/B sky130_fd_sc_hd__nand2_1
X_07827_ _08067_/B _08067_/A vssd1 vssd1 vccd1 vccd1 _07831_/A sky130_fd_sc_hd__nor2_1
X_07758_ _07758_/A _07758_/B vssd1 vssd1 vccd1 vccd1 _07782_/B sky130_fd_sc_hd__nand2_1
XANTENNA__08784__A _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06709_ _05960_/B _06707_/Y _06708_/Y vssd1 vssd1 vccd1 vccd1 _06816_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07689_ _07689_/A _07689_/B vssd1 vssd1 vccd1 vccd1 _07691_/A sky130_fd_sc_hd__nand2_1
X_09428_ _09426_/X _09428_/B vssd1 vssd1 vccd1 vccd1 _09430_/A sky130_fd_sc_hd__and2b_1
X_09359_ _10348_/A _10348_/B vssd1 vssd1 vccd1 vccd1 _10347_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_22_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10203_ _09677_/A _09698_/A _10004_/A _09477_/C vssd1 vssd1 vccd1 vccd1 _10204_/B
+ sky130_fd_sc_hd__a22o_1
X_10134_ _10134_/A _10134_/B vssd1 vssd1 vccd1 vccd1 _10136_/A sky130_fd_sc_hd__xor2_1
X_10065_ _10065_/A _10300_/A vssd1 vssd1 vccd1 vccd1 _10067_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_57_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05830__B _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ _07008_/A vssd1 vssd1 vccd1 vccd1 _06995_/A sky130_fd_sc_hd__inv_2
X_08730_ _09261_/B _08731_/C _08729_/Y vssd1 vssd1 vccd1 vccd1 _08732_/A sky130_fd_sc_hd__a21bo_1
X_05942_ _05942_/A _05942_/B vssd1 vssd1 vccd1 vccd1 _05946_/C sky130_fd_sc_hd__nand2_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06389__A _09517_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08661_ _08661_/A _08661_/B vssd1 vssd1 vccd1 vccd1 _08663_/A sky130_fd_sc_hd__nand2_1
X_05873_ _05877_/A vssd1 vssd1 vccd1 vccd1 _05876_/A sky130_fd_sc_hd__inv_2
X_07612_ _07714_/B _07612_/B _07612_/C vssd1 vssd1 vccd1 vccd1 _07714_/A sky130_fd_sc_hd__nand3_1
X_08592_ _08592_/A vssd1 vssd1 vccd1 vccd1 _08593_/B sky130_fd_sc_hd__inv_2
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07543_ _07543_/A _07543_/B _07546_/A vssd1 vssd1 vccd1 vccd1 _07548_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_48_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07474_ _07543_/B _07546_/A _07473_/Y vssd1 vssd1 vccd1 vccd1 _07477_/A sky130_fd_sc_hd__a21oi_2
X_09213_ _09213_/A _09213_/B vssd1 vssd1 vccd1 vccd1 _09218_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_8_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06425_ _06425_/A _06425_/B _06425_/C vssd1 vssd1 vccd1 vccd1 _06428_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_56_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09144_ _09145_/A _09144_/B vssd1 vssd1 vccd1 vccd1 _09154_/B sky130_fd_sc_hd__nand2b_1
XANTENNA__06852__A _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06356_ _06360_/B _06357_/A vssd1 vssd1 vccd1 vccd1 _06359_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_71_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09075_ _09077_/B vssd1 vssd1 vccd1 vccd1 _09076_/B sky130_fd_sc_hd__inv_2
X_06287_ _06431_/A _06430_/A vssd1 vssd1 vccd1 vccd1 _06287_/Y sky130_fd_sc_hd__nor2_1
X_08026_ _08026_/A _08026_/B vssd1 vssd1 vccd1 vccd1 _08026_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10093__B _10334_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09977_ _10127_/A _09977_/B vssd1 vssd1 vccd1 vccd1 _09981_/B sky130_fd_sc_hd__nand2_1
X_08928_ _08928_/A _08928_/B vssd1 vssd1 vccd1 vccd1 _08937_/B sky130_fd_sc_hd__nand2_1
X_08859_ _08859_/A _08859_/B _08859_/C vssd1 vssd1 vccd1 vccd1 _08860_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_79_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10683_ _10683_/A hold37/X vssd1 vssd1 vccd1 vccd1 hold38/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10117_ _10115_/Y _10117_/B _10117_/C vssd1 vssd1 vccd1 vccd1 _10118_/B sky130_fd_sc_hd__nand3b_1
X_10048_ _10048_/A _10048_/B _10048_/C vssd1 vssd1 vccd1 vccd1 _10049_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_26_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06210_ _06210_/A _06210_/B vssd1 vssd1 vccd1 vccd1 _06386_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07190_ _07167_/C _07167_/B _07187_/Y vssd1 vssd1 vccd1 vccd1 _07201_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07487__B _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06141_ _06324_/C vssd1 vssd1 vccd1 vccd1 _06143_/B sky130_fd_sc_hd__inv_2
X_06072_ _06072_/A _06072_/B vssd1 vssd1 vccd1 vccd1 _06075_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_41_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09900_ _10306_/A _09900_/B _10319_/A vssd1 vssd1 vccd1 vccd1 _09907_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_6_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09831_ _09831_/A _09831_/B vssd1 vssd1 vccd1 vccd1 _09833_/A sky130_fd_sc_hd__nor2_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ _09762_/A _09859_/A vssd1 vssd1 vccd1 vccd1 _09764_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_67_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05735__B _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06974_ _06976_/A _06974_/B vssd1 vssd1 vccd1 vccd1 _06975_/B sky130_fd_sc_hd__nand2_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _08777_/C _08763_/B vssd1 vssd1 vccd1 vccd1 _08715_/A sky130_fd_sc_hd__nand2_1
X_05925_ _06755_/B _05929_/B vssd1 vssd1 vccd1 vccd1 _05927_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08111__B _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09693_ _09695_/B vssd1 vssd1 vccd1 vccd1 _10059_/B sky130_fd_sc_hd__inv_2
X_08644_ _08654_/B _09216_/B vssd1 vssd1 vccd1 vccd1 _08653_/A sky130_fd_sc_hd__nand2_1
X_05856_ _05858_/B _05857_/B _05857_/A vssd1 vssd1 vccd1 vccd1 _06113_/C sky130_fd_sc_hd__nand3b_1
X_05787_ _05789_/B _06040_/B _05788_/B vssd1 vssd1 vccd1 vccd1 _06040_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__05751__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08575_ _08576_/A _08576_/B vssd1 vssd1 vccd1 vccd1 _09135_/B sky130_fd_sc_hd__or2_1
X_07526_ _07682_/B vssd1 vssd1 vccd1 vccd1 _07674_/B sky130_fd_sc_hd__inv_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07457_ _07530_/A _07531_/A vssd1 vssd1 vccd1 vccd1 _07535_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_44_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07388_ _07449_/A _07449_/B _07448_/B vssd1 vssd1 vccd1 vccd1 _07397_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07678__A _08724_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06582__A _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06408_ _06403_/Y _06569_/B _06407_/Y vssd1 vssd1 vccd1 vccd1 _06409_/B sky130_fd_sc_hd__a21oi_1
X_09127_ _09130_/A _09576_/B vssd1 vssd1 vccd1 vccd1 _09128_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06339_ _10210_/B _07897_/B vssd1 vssd1 vccd1 vccd1 _06508_/C sky130_fd_sc_hd__nand2_1
X_09058_ _09058_/A _09058_/B vssd1 vssd1 vccd1 vccd1 _09328_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08009_ _08009_/A vssd1 vssd1 vccd1 vccd1 _08010_/A sky130_fd_sc_hd__inv_2
XANTENNA__05926__A _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08021__B _09971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05661__A _08453_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10735_ _10741_/CLK hold19/X fanout98/X vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10666_ _10666_/A vssd1 vssd1 vccd1 vccd1 _10718_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10597_ _10597_/A _10605_/B _10605_/A vssd1 vssd1 vccd1 vccd1 _10630_/A sky130_fd_sc_hd__nand3_2
XFILLER_0_2_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput80 hold15/A vssd1 vssd1 vccd1 vccd1 y_o[22] sky130_fd_sc_hd__buf_12
Xoutput91 hold58/A vssd1 vssd1 vccd1 vccd1 y_o[3] sky130_fd_sc_hd__buf_12
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05710_ _05712_/B _05712_/C vssd1 vssd1 vccd1 vccd1 _05839_/B sky130_fd_sc_hd__nand2_1
X_06690_ _06690_/A _06690_/B vssd1 vssd1 vccd1 vccd1 _06693_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_77_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08350__A1 _09875_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05641_ _08101_/B input5/X vssd1 vssd1 vccd1 vccd1 _05696_/B sky130_fd_sc_hd__nand2_1
X_08360_ _08360_/A _08361_/B _08360_/C vssd1 vssd1 vccd1 vccd1 _10517_/B sky130_fd_sc_hd__nand3_1
X_05572_ _05577_/A _05577_/C vssd1 vssd1 vccd1 vccd1 _05575_/A sky130_fd_sc_hd__nand2_1
X_07311_ _07311_/A _07311_/B vssd1 vssd1 vccd1 vccd1 _07315_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09697__B _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08291_ _08291_/A _08291_/B vssd1 vssd1 vccd1 vccd1 _08359_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07242_ _07242_/A _07415_/A vssd1 vssd1 vccd1 vccd1 _07243_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_73_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07173_ _10040_/B _10130_/A vssd1 vssd1 vccd1 vccd1 _07349_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06124_ _06124_/A _06124_/B vssd1 vssd1 vccd1 vccd1 _06125_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_5_199 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06055_ _06054_/B _06869_/B _06055_/C vssd1 vssd1 vccd1 vccd1 _06869_/A sky130_fd_sc_hd__nand3b_2
X_09814_ _09819_/B _09835_/B vssd1 vssd1 vccd1 vccd1 _09818_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05465__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07961__A _08059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09745_ input49/X input50/X _10247_/B _09840_/B vssd1 vssd1 vccd1 vccd1 _09746_/A
+ sky130_fd_sc_hd__and4_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06957_ _06957_/A _06957_/B _06957_/C vssd1 vssd1 vccd1 vccd1 _06965_/A sky130_fd_sc_hd__nand3_1
X_09676_ _09676_/A vssd1 vssd1 vccd1 vccd1 _09687_/B sky130_fd_sc_hd__inv_2
X_06888_ _08984_/A _06888_/B _06888_/C vssd1 vssd1 vccd1 vccd1 _06895_/B sky130_fd_sc_hd__nand3_1
X_05908_ _08114_/B _10157_/B vssd1 vssd1 vccd1 vccd1 _05910_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_68_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08627_ _08627_/A _08627_/B vssd1 vssd1 vccd1 vccd1 _08666_/C sky130_fd_sc_hd__nand2_1
X_05839_ _05839_/A _05839_/B vssd1 vssd1 vccd1 vccd1 _05839_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08558_ _08558_/A _08558_/B vssd1 vssd1 vccd1 vccd1 _08560_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08489_ _08489_/A _08489_/B vssd1 vssd1 vccd1 vccd1 _08550_/B sky130_fd_sc_hd__nand2_1
X_07509_ _07509_/A _07509_/B _07509_/C vssd1 vssd1 vccd1 vccd1 _07512_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_64_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10520_ _10520_/A hold23/X _10520_/C vssd1 vssd1 vccd1 vccd1 _10641_/B sky130_fd_sc_hd__nand3_1
X_10451_ _10451_/A _10452_/A vssd1 vssd1 vccd1 vccd1 _10460_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10203__A2 _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10382_ _10566_/A vssd1 vssd1 vccd1 vccd1 _10383_/B sky130_fd_sc_hd__inv_2
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05375__B _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08686__B _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10718_ _10718_/CLK _10718_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10649_ _10649_/A _10649_/B vssd1 vssd1 vccd1 vccd1 _10653_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07860_ _10426_/B _10431_/B vssd1 vssd1 vccd1 vccd1 _10403_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_64_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06811_ _06811_/A _06811_/B vssd1 vssd1 vccd1 vccd1 _08976_/A sky130_fd_sc_hd__nand2_1
X_07791_ _07791_/A vssd1 vssd1 vccd1 vccd1 _07793_/B sky130_fd_sc_hd__inv_2
X_09530_ _09530_/A vssd1 vssd1 vccd1 vccd1 _09532_/B sky130_fd_sc_hd__inv_2
X_06742_ _06768_/B _08552_/A vssd1 vssd1 vccd1 vccd1 _06767_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_3_78 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06397__A _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09461_ _09461_/A vssd1 vssd1 vccd1 vccd1 _09463_/C sky130_fd_sc_hd__inv_2
XFILLER_0_78_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06673_ _06948_/C _06671_/Y _06672_/Y vssd1 vssd1 vccd1 vccd1 _06939_/B sky130_fd_sc_hd__o21bai_1
X_08412_ _08412_/A vssd1 vssd1 vccd1 vccd1 _08413_/B sky130_fd_sc_hd__inv_2
X_05624_ _05626_/B _05625_/A _05625_/B vssd1 vssd1 vccd1 vccd1 _05627_/A sky130_fd_sc_hd__nand3b_1
X_09392_ input20/X vssd1 vssd1 vccd1 vccd1 _09393_/B sky130_fd_sc_hd__inv_2
XFILLER_0_58_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_05555_ _05560_/A _05560_/C vssd1 vssd1 vccd1 vccd1 _05558_/A sky130_fd_sc_hd__nand2_1
X_08343_ _08352_/A vssd1 vssd1 vccd1 vccd1 _08344_/B sky130_fd_sc_hd__inv_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08274_ _08292_/A _08292_/B _08293_/A vssd1 vssd1 vccd1 vccd1 _08324_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_73_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05486_ _05948_/B vssd1 vssd1 vccd1 vccd1 _05487_/B sky130_fd_sc_hd__inv_2
X_07225_ _07233_/B _07225_/B vssd1 vssd1 vccd1 vccd1 _07398_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_13_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07156_ _07311_/A _07312_/A vssd1 vssd1 vccd1 vccd1 _07156_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07087_ _08897_/B _10148_/A vssd1 vssd1 vccd1 vccd1 _07229_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07675__B _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06107_ _06227_/C _06227_/B _05747_/Y vssd1 vssd1 vccd1 vccd1 _06108_/B sky130_fd_sc_hd__a21o_1
X_06038_ _06038_/A _06841_/A _06846_/A vssd1 vssd1 vccd1 vccd1 _06042_/C sky130_fd_sc_hd__nand3_1
X_09728_ _09896_/B _09728_/B vssd1 vssd1 vccd1 vccd1 _09733_/B sky130_fd_sc_hd__nand2_1
X_07989_ _07989_/A _07990_/A vssd1 vssd1 vccd1 vccd1 _07992_/A sky130_fd_sc_hd__nand2_1
X_09659_ _09659_/A _09932_/A vssd1 vssd1 vccd1 vccd1 _09660_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_291 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10503_ _10503_/A _10503_/B vssd1 vssd1 vccd1 vccd1 _10541_/A sky130_fd_sc_hd__nor2_1
X_10434_ _10434_/A _10434_/B vssd1 vssd1 vccd1 vccd1 _10443_/A sky130_fd_sc_hd__nand2_1
X_10365_ _10364_/B _10560_/B _10365_/C vssd1 vssd1 vccd1 vccd1 _10369_/B sky130_fd_sc_hd__nand3b_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ _10298_/A vssd1 vssd1 vccd1 vccd1 _10297_/B sky130_fd_sc_hd__inv_2
XANTENNA__08697__A _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09678__D _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05340_ input9/X vssd1 vssd1 vccd1 vccd1 _10148_/B sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07010_ _07032_/A vssd1 vssd1 vccd1 vccd1 _07011_/B sky130_fd_sc_hd__inv_2
XFILLER_0_59_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08961_ _08961_/A _08969_/B _08969_/A vssd1 vssd1 vccd1 vccd1 _09031_/B sky130_fd_sc_hd__nand3_1
X_08892_ _08959_/A _08959_/B vssd1 vssd1 vccd1 vccd1 _08958_/A sky130_fd_sc_hd__nand2_1
X_07912_ _07912_/A _07912_/B vssd1 vssd1 vccd1 vccd1 _07914_/A sky130_fd_sc_hd__nand2_1
X_07843_ _07843_/A _07850_/B _07843_/C vssd1 vssd1 vccd1 vccd1 _07852_/A sky130_fd_sc_hd__nand3_1
X_07774_ _07799_/A _07800_/A vssd1 vssd1 vccd1 vccd1 _07775_/A sky130_fd_sc_hd__nand2_1
X_09513_ _09513_/A _09513_/B vssd1 vssd1 vccd1 vccd1 _09570_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07016__A _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06725_ _08573_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _06728_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09444_ _09444_/A _09444_/B vssd1 vssd1 vccd1 vccd1 _09446_/A sky130_fd_sc_hd__nand2_1
X_06656_ _06957_/A _06962_/A vssd1 vssd1 vccd1 vccd1 _06656_/Y sky130_fd_sc_hd__nor2_1
X_05607_ input36/X vssd1 vssd1 vccd1 vccd1 _10151_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09375_ _09373_/Y _09375_/B vssd1 vssd1 vccd1 vccd1 _09376_/B sky130_fd_sc_hd__and2b_1
XFILLER_0_19_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06587_ _09749_/B _10151_/A vssd1 vssd1 vccd1 vccd1 _06590_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08326_ _08357_/B _08357_/A vssd1 vssd1 vccd1 vccd1 _08326_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_19_367 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05538_ input2/X vssd1 vssd1 vccd1 vccd1 _08672_/A sky130_fd_sc_hd__buf_6
XFILLER_0_34_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08257_ _10275_/B _10115_/A vssd1 vssd1 vccd1 vccd1 _08304_/A sky130_fd_sc_hd__nand2_1
X_05469_ _08114_/B _10156_/B vssd1 vssd1 vccd1 vccd1 _05472_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07208_ _07236_/B _07236_/C vssd1 vssd1 vccd1 vccd1 _07235_/A sky130_fd_sc_hd__nand2_1
X_08188_ _08897_/B _10130_/A vssd1 vssd1 vccd1 vccd1 _08192_/B sky130_fd_sc_hd__nand2_1
X_07139_ _07139_/A _07139_/B _07139_/C vssd1 vssd1 vccd1 vccd1 _07303_/C sky130_fd_sc_hd__nand3_1
X_10150_ _10150_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _10152_/A sky130_fd_sc_hd__nand2_1
X_10081_ _10087_/A _10087_/C vssd1 vssd1 vccd1 vccd1 _10085_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10725__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_112 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10417_ _10417_/A hold36/X vssd1 vssd1 vccd1 vccd1 _10682_/B sky130_fd_sc_hd__nand2_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _10348_/A _10348_/B _10348_/C vssd1 vssd1 vccd1 vccd1 _10376_/B sky130_fd_sc_hd__nand3_1
X_10279_ _10279_/A _10279_/B vssd1 vssd1 vccd1 vccd1 _10282_/B sky130_fd_sc_hd__xnor2_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_2_2__f_clk_A clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07490_ _07486_/Y _07488_/Y _07648_/A vssd1 vssd1 vccd1 vccd1 _07492_/A sky130_fd_sc_hd__a21oi_1
X_06510_ _08171_/B vssd1 vssd1 vccd1 vccd1 _10103_/B sky130_fd_sc_hd__buf_6
XFILLER_0_61_43 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06441_ _06616_/B _06616_/C vssd1 vssd1 vccd1 vccd1 _06615_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09160_ _09181_/A _09409_/B vssd1 vssd1 vccd1 vccd1 _09179_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06372_ _06372_/A _06372_/B vssd1 vssd1 vccd1 vccd1 _06659_/B sky130_fd_sc_hd__nand2_1
X_09091_ _09091_/A vssd1 vssd1 vccd1 vccd1 _09096_/B sky130_fd_sc_hd__inv_2
XFILLER_0_9_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08111_ _09749_/B _08573_/A vssd1 vssd1 vccd1 vccd1 _08164_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08042_ _08042_/A _08043_/A _08043_/B vssd1 vssd1 vccd1 vccd1 _08091_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_71_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08114__B _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09993_ _09993_/A _09993_/B _09993_/C vssd1 vssd1 vccd1 vccd1 _09995_/B sky130_fd_sc_hd__nand3_1
X_08944_ _08946_/B vssd1 vssd1 vccd1 vccd1 _08945_/B sky130_fd_sc_hd__inv_2
X_08875_ _08874_/B _08875_/B _08875_/C vssd1 vssd1 vccd1 vccd1 _08876_/B sky130_fd_sc_hd__nand3b_1
X_07826_ _08066_/B _08066_/C vssd1 vssd1 vccd1 vccd1 _08067_/A sky130_fd_sc_hd__nand2_1
X_07757_ _07759_/B vssd1 vssd1 vccd1 vccd1 _07758_/B sky130_fd_sc_hd__inv_2
X_06708_ _06708_/A _06708_/B vssd1 vssd1 vccd1 vccd1 _06708_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_66_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07688_ _07688_/A _07688_/B vssd1 vssd1 vccd1 vccd1 _07799_/B sky130_fd_sc_hd__nand2_2
X_09427_ _10151_/A _09922_/B _10150_/A _09602_/B vssd1 vssd1 vccd1 vccd1 _09428_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06639_ _06641_/A _06639_/B vssd1 vssd1 vccd1 vccd1 _06640_/B sky130_fd_sc_hd__nand2_1
X_09358_ _09358_/A _09358_/B vssd1 vssd1 vccd1 vccd1 _10348_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_47_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08309_ _08351_/A _10292_/B _10108_/B vssd1 vssd1 vccd1 vccd1 _08312_/C sky130_fd_sc_hd__and3_1
XFILLER_0_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09289_ _09289_/A _09289_/B vssd1 vssd1 vccd1 vccd1 _09292_/C sky130_fd_sc_hd__nor2_1
XFILLER_0_22_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10202_ _10202_/A _10202_/B _10202_/C _10202_/D vssd1 vssd1 vccd1 vccd1 _10204_/A
+ sky130_fd_sc_hd__or4_1
X_10133_ _09958_/A _09958_/B _09957_/A vssd1 vssd1 vccd1 vccd1 _10134_/B sky130_fd_sc_hd__o21a_1
X_10064_ _10064_/A _10064_/B _10300_/B vssd1 vssd1 vccd1 vccd1 _10300_/A sky130_fd_sc_hd__nand3_1
XANTENNA__09136__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05574__A _07675_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _06995_/B _07008_/A vssd1 vssd1 vccd1 vccd1 _06994_/A sky130_fd_sc_hd__nand2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05941_ _05942_/A _05942_/B vssd1 vssd1 vccd1 vccd1 _06760_/B sky130_fd_sc_hd__or2_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06389__B input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08660_ _08660_/A _08660_/B vssd1 vssd1 vccd1 vccd1 _08661_/B sky130_fd_sc_hd__nand2_1
X_05872_ _09517_/D _09678_/C vssd1 vssd1 vccd1 vccd1 _05877_/A sky130_fd_sc_hd__nand2_1
X_07611_ _07613_/B _07614_/B _07614_/C vssd1 vssd1 vccd1 vccd1 _07714_/B sky130_fd_sc_hd__nand3_1
X_08591_ _08587_/Y _08589_/Y _08592_/A vssd1 vssd1 vccd1 vccd1 _08594_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_72_64 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07542_ _07544_/B _07545_/B _07545_/A vssd1 vssd1 vccd1 vccd1 _07543_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07473_ _07545_/C _07544_/A vssd1 vssd1 vccd1 vccd1 _07473_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09212_ _09214_/C vssd1 vssd1 vccd1 vccd1 _09213_/B sky130_fd_sc_hd__inv_2
X_06424_ _06424_/A _06424_/B vssd1 vssd1 vccd1 vccd1 _06428_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06355_ _06358_/B vssd1 vssd1 vccd1 vccd1 _06360_/B sky130_fd_sc_hd__inv_2
X_09143_ _09145_/B _09145_/C vssd1 vssd1 vccd1 vccd1 _09144_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06852__B _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09074_ _09336_/A _09335_/A vssd1 vssd1 vccd1 vccd1 _09077_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_44_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06286_ _06432_/C vssd1 vssd1 vccd1 vccd1 _06422_/C sky130_fd_sc_hd__inv_2
X_08025_ _08025_/A _08025_/B vssd1 vssd1 vccd1 vccd1 _08141_/B sky130_fd_sc_hd__nand2_1
XANTENNA__10093__C _10093_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09976_ _09976_/A _09976_/B vssd1 vssd1 vccd1 vccd1 _09977_/B sky130_fd_sc_hd__nand2_1
X_08927_ _08927_/A _08927_/B vssd1 vssd1 vccd1 vccd1 _08928_/B sky130_fd_sc_hd__nand2_1
X_08858_ _08858_/A _08858_/B vssd1 vssd1 vccd1 vccd1 _08860_/A sky130_fd_sc_hd__nand2_1
X_07809_ _07809_/A _07809_/B vssd1 vssd1 vccd1 vccd1 _07811_/A sky130_fd_sc_hd__nand2_1
X_08789_ _08783_/Y _08790_/B _08789_/C vssd1 vssd1 vccd1 vccd1 _08846_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_82_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10682_ _10682_/A _10682_/B vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__nand2_1
XANTENNA__10284__B _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05659__A _07785_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10740__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ _10117_/B _10117_/C _10115_/Y vssd1 vssd1 vccd1 vccd1 _10118_/A sky130_fd_sc_hd__a21bo_1
X_10047_ _10047_/A vssd1 vssd1 vccd1 vccd1 _10048_/B sky130_fd_sc_hd__inv_2
XFILLER_0_26_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06140_ _07756_/A _07897_/B vssd1 vssd1 vccd1 vccd1 _06324_/C sky130_fd_sc_hd__nand2_1
X_06071_ _06071_/A _06071_/B _06071_/C vssd1 vssd1 vccd1 vccd1 _06072_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_6_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09830_ _10347_/A _09830_/B vssd1 vssd1 vccd1 vccd1 _10569_/A sky130_fd_sc_hd__nand2_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _09859_/B _09761_/B _09761_/C vssd1 vssd1 vccd1 vccd1 _09859_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_67_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ _06973_/A vssd1 vssd1 vccd1 vccd1 _06976_/A sky130_fd_sc_hd__inv_2
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _08763_/A _08763_/B _08764_/A vssd1 vssd1 vccd1 vccd1 _08777_/C sky130_fd_sc_hd__nand3_1
X_05924_ _05924_/A _05924_/B vssd1 vssd1 vccd1 vccd1 _05929_/B sky130_fd_sc_hd__nand2_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ _09692_/A _09692_/B vssd1 vssd1 vccd1 vccd1 _09695_/B sky130_fd_sc_hd__nand2_1
X_08643_ _08642_/B _08643_/B _08643_/C vssd1 vssd1 vccd1 vccd1 _09216_/B sky130_fd_sc_hd__nand3b_1
X_05855_ _05855_/A _05855_/B vssd1 vssd1 vccd1 vccd1 _05857_/A sky130_fd_sc_hd__nand2_1
X_05786_ _05786_/A _05786_/B vssd1 vssd1 vccd1 vccd1 _05788_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05751__B input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08574_ _08574_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _08576_/B sky130_fd_sc_hd__nand2_1
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07525_ _07756_/A input44/X vssd1 vssd1 vccd1 vccd1 _07682_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06863__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07456_ _08337_/A _08453_/A vssd1 vssd1 vccd1 vccd1 _07531_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07387_ _07449_/C vssd1 vssd1 vccd1 vccd1 _07448_/B sky130_fd_sc_hd__inv_2
XANTENNA__07678__B _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06582__B _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06407_ _06567_/A _06566_/A vssd1 vssd1 vccd1 vccd1 _06407_/Y sky130_fd_sc_hd__nor2_1
X_09126_ _09126_/A _09126_/B _09564_/A vssd1 vssd1 vccd1 vccd1 _09576_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06338_ _06507_/A _06506_/A vssd1 vssd1 vccd1 vccd1 _06343_/B sky130_fd_sc_hd__nand2_1
X_09057_ _09059_/B _09059_/C vssd1 vssd1 vccd1 vccd1 _09058_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_44_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06269_ _06431_/B _06431_/C vssd1 vssd1 vccd1 vccd1 _06430_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_435 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08008_ _08008_/A _08009_/A vssd1 vssd1 vccd1 vccd1 _08199_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_12_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05926__B _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _09959_/A vssd1 vssd1 vccd1 vccd1 _09961_/B sky130_fd_sc_hd__inv_2
XANTENNA__09414__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05661__B _07891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10734_ _10741_/CLK _10734_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold65/A sky130_fd_sc_hd__dfrtp_2
XFILLER_0_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10665_ _10665_/A _10668_/A vssd1 vssd1 vccd1 vccd1 _10666_/A sky130_fd_sc_hd__and2_1
X_10596_ _10596_/A _10596_/B vssd1 vssd1 vccd1 vccd1 _10605_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput70 hold62/A vssd1 vssd1 vccd1 vccd1 y_o[13] sky130_fd_sc_hd__buf_12
Xoutput81 hold7/A vssd1 vssd1 vccd1 vccd1 y_o[23] sky130_fd_sc_hd__buf_12
Xoutput92 hold46/A vssd1 vssd1 vccd1 vccd1 y_o[4] sky130_fd_sc_hd__buf_12
X_05640_ _05640_/A _05640_/B vssd1 vssd1 vccd1 vccd1 _06229_/B sky130_fd_sc_hd__nand2_2
X_05571_ _05571_/A _05571_/B vssd1 vssd1 vccd1 vccd1 _05577_/C sky130_fd_sc_hd__nand2_1
X_07310_ _07312_/A vssd1 vssd1 vccd1 vccd1 _07311_/B sky130_fd_sc_hd__inv_2
XFILLER_0_73_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08290_ _08290_/A _08325_/A vssd1 vssd1 vccd1 vccd1 _08291_/B sky130_fd_sc_hd__nand2_1
X_07241_ _07289_/A _07287_/A vssd1 vssd1 vccd1 vccd1 _07241_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_26_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07172_ _07305_/B _07303_/A vssd1 vssd1 vccd1 vccd1 _07172_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_14_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06123_ _06234_/B _06234_/C vssd1 vssd1 vccd1 vccd1 _06233_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06054_ _06054_/A _06054_/B vssd1 vssd1 vccd1 vccd1 _06060_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_22_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09813_ _09813_/A _09813_/B _09836_/A vssd1 vssd1 vccd1 vccd1 _09835_/B sky130_fd_sc_hd__nand3_1
XANTENNA__07019__A _09710_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09744_ _09744_/A _09744_/B vssd1 vssd1 vccd1 vccd1 _09764_/B sky130_fd_sc_hd__and2_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06956_ _07113_/B _07113_/C vssd1 vssd1 vccd1 vccd1 _07115_/A sky130_fd_sc_hd__nand2_1
X_09675_ _09428_/B _10187_/A _10148_/A _09426_/X vssd1 vssd1 vccd1 vccd1 _09676_/A
+ sky130_fd_sc_hd__a31o_1
X_06887_ _06887_/A _06887_/B vssd1 vssd1 vccd1 vccd1 _06895_/A sky130_fd_sc_hd__nand2_1
X_05907_ _06734_/B _05911_/C vssd1 vssd1 vccd1 vccd1 _05909_/A sky130_fd_sc_hd__nand2_1
X_08626_ _08547_/A _08547_/C _08570_/B vssd1 vssd1 vccd1 vccd1 _08627_/B sky130_fd_sc_hd__a21boi_1
X_05838_ _05839_/B _05839_/A vssd1 vssd1 vccd1 vccd1 _05838_/Y sky130_fd_sc_hd__nand2_1
X_08557_ _08559_/B _08559_/C vssd1 vssd1 vccd1 vccd1 _08558_/A sky130_fd_sc_hd__nand2_1
X_05769_ _09517_/C _09678_/C vssd1 vssd1 vccd1 vccd1 _05773_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08488_ _08488_/A _08488_/B vssd1 vssd1 vccd1 vccd1 _08489_/B sky130_fd_sc_hd__nand2_1
X_07508_ _07508_/A _07508_/B vssd1 vssd1 vccd1 vccd1 _07512_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07439_ _07439_/A _07439_/B vssd1 vssd1 vccd1 vccd1 _07604_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10450_ _10542_/B _10453_/B vssd1 vssd1 vccd1 vccd1 _10451_/A sky130_fd_sc_hd__nand2_1
X_09109_ _09109_/A _09109_/B vssd1 vssd1 vccd1 vccd1 _09114_/B sky130_fd_sc_hd__nand2_1
X_10381_ _10704_/A _10704_/B _10701_/B vssd1 vssd1 vccd1 vccd1 _10566_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_20_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08313__A _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10717_ _10718_/CLK hold35/X fanout99/X vssd1 vssd1 vccd1 vccd1 hold57/A sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10648_ _10649_/B _10649_/A vssd1 vssd1 vccd1 vccd1 _10650_/A sky130_fd_sc_hd__or2_1
X_10579_ _10707_/B _10707_/A _10603_/A vssd1 vssd1 vccd1 vccd1 _10584_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_23_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06810_ _06810_/A _06810_/B vssd1 vssd1 vccd1 vccd1 _06811_/B sky130_fd_sc_hd__nand2_1
X_07790_ _09778_/D _07897_/B vssd1 vssd1 vccd1 vccd1 _07791_/A sky130_fd_sc_hd__nand2_1
X_06741_ _06767_/B _08552_/A _06768_/B vssd1 vssd1 vccd1 vccd1 _08881_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09460_ _09205_/A _09204_/B _09459_/Y vssd1 vssd1 vccd1 vccd1 _09461_/A sky130_fd_sc_hd__o21a_1
XFILLER_0_78_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08411_ _08407_/Y _08409_/Y _08412_/A vssd1 vssd1 vccd1 vccd1 _08414_/A sky130_fd_sc_hd__o21ai_1
X_06672_ _06943_/A _06945_/A vssd1 vssd1 vccd1 vccd1 _06672_/Y sky130_fd_sc_hd__nor2_1
X_05623_ _06078_/A _05623_/B _05623_/C vssd1 vssd1 vccd1 vccd1 _05625_/B sky130_fd_sc_hd__nand3_1
X_09391_ _09391_/A _09391_/B vssd1 vssd1 vccd1 vccd1 _09397_/A sky130_fd_sc_hd__nand2_1
X_05554_ _05600_/A _05600_/B vssd1 vssd1 vccd1 vccd1 _05560_/C sky130_fd_sc_hd__nand2_1
X_08342_ _09875_/D _09393_/A _08342_/C vssd1 vssd1 vccd1 vccd1 _08352_/A sky130_fd_sc_hd__or3_1
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05485_ _08337_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _05948_/B sky130_fd_sc_hd__nand2_1
X_08273_ _08320_/B _08320_/A vssd1 vssd1 vccd1 vccd1 _08293_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_61_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07224_ _07233_/A vssd1 vssd1 vccd1 vccd1 _07225_/B sky130_fd_sc_hd__inv_2
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07155_ _07323_/C _07323_/B _07154_/Y vssd1 vssd1 vccd1 vccd1 _07312_/A sky130_fd_sc_hd__a21oi_2
X_06106_ _06106_/A _06106_/B _06106_/C vssd1 vssd1 vccd1 vccd1 _06111_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_14_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07086_ _10292_/B _09678_/C vssd1 vssd1 vccd1 vccd1 _07414_/B sky130_fd_sc_hd__nand2_1
X_06037_ _06846_/B _06037_/B vssd1 vssd1 vccd1 vccd1 _06042_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07988_ _08112_/A _08101_/B vssd1 vssd1 vccd1 vccd1 _07990_/A sky130_fd_sc_hd__nand2_1
X_09727_ _09896_/A vssd1 vssd1 vccd1 vccd1 _09728_/B sky130_fd_sc_hd__inv_2
X_06939_ _06939_/A _06939_/B vssd1 vssd1 vccd1 vccd1 _06941_/B sky130_fd_sc_hd__nand2_1
X_09658_ _09932_/B _09658_/B _09658_/C vssd1 vssd1 vccd1 vccd1 _09932_/A sky130_fd_sc_hd__nand3_1
X_09589_ _09589_/A _10353_/C vssd1 vssd1 vccd1 vccd1 _10348_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_49_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08609_ _08609_/A _08609_/B vssd1 vssd1 vccd1 vccd1 _08611_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10502_ _10510_/A _10502_/B vssd1 vssd1 vccd1 vccd1 _10503_/B sky130_fd_sc_hd__nor2_1
X_10433_ hold63/A vssd1 vssd1 vccd1 vccd1 _10434_/B sky130_fd_sc_hd__inv_2
X_10364_ _10364_/A _10364_/B vssd1 vssd1 vccd1 vccd1 _10369_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09139__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10292__B _10292_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10295_ _10295_/A _10295_/B vssd1 vssd1 vccd1 vccd1 _10298_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08697__B _10005_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09602__A _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08218__A _08218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_43_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_59_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08960_ _09016_/B _09016_/C vssd1 vssd1 vccd1 vccd1 _09313_/B sky130_fd_sc_hd__nand2_1
X_08891_ _09082_/A _08891_/B _09133_/A vssd1 vssd1 vccd1 vccd1 _08959_/B sky130_fd_sc_hd__nand3_1
X_07911_ _07913_/A _07913_/C vssd1 vssd1 vccd1 vccd1 _07912_/A sky130_fd_sc_hd__nand2_1
X_07842_ _08075_/A _07842_/B vssd1 vssd1 vccd1 vccd1 _07843_/A sky130_fd_sc_hd__nor2_1
X_09512_ _09512_/A _09512_/B vssd1 vssd1 vccd1 vccd1 _09513_/B sky130_fd_sc_hd__and2_1
X_07773_ _07799_/B vssd1 vssd1 vccd1 vccd1 _07800_/A sky130_fd_sc_hd__inv_2
X_06724_ _06724_/A _08432_/A vssd1 vssd1 vccd1 vccd1 _06740_/B sky130_fd_sc_hd__nand2_1
XANTENNA__07016__B _07891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09443_ _09442_/B _09443_/B _09443_/C vssd1 vssd1 vccd1 vccd1 _09444_/B sky130_fd_sc_hd__nand3b_1
X_06655_ _06965_/C vssd1 vssd1 vccd1 vccd1 _06964_/B sky130_fd_sc_hd__inv_2
X_05606_ _08724_/A input37/X vssd1 vssd1 vccd1 vccd1 _05611_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09374_ _09393_/A _09373_/B _09373_/C vssd1 vssd1 vccd1 vccd1 _09375_/B sky130_fd_sc_hd__o21ai_1
X_06586_ _09517_/D vssd1 vssd1 vccd1 vccd1 _09749_/B sky130_fd_sc_hd__buf_12
X_08325_ _08325_/A _08325_/B vssd1 vssd1 vccd1 vccd1 _08357_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05537_ _05892_/B _05892_/A vssd1 vssd1 vccd1 vccd1 _05629_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_240 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08256_ _10284_/B _10108_/B _10292_/B _10112_/A vssd1 vssd1 vccd1 vccd1 _08303_/A
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05468_ _05471_/A _05913_/B vssd1 vssd1 vccd1 vccd1 _05470_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_6_295 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08187_ _08195_/B _08195_/A vssd1 vssd1 vccd1 vccd1 _08271_/B sky130_fd_sc_hd__nand2_1
X_07207_ _07207_/A _07207_/B vssd1 vssd1 vccd1 vccd1 _07236_/C sky130_fd_sc_hd__nand2_1
X_07138_ _07138_/A _07138_/B _07138_/C vssd1 vssd1 vccd1 vccd1 _07139_/B sky130_fd_sc_hd__nand3_1
X_05399_ input7/X vssd1 vssd1 vccd1 vccd1 _09602_/B sky130_fd_sc_hd__clkbuf_8
X_07069_ _07069_/A _07069_/B vssd1 vssd1 vccd1 vccd1 _07125_/C sky130_fd_sc_hd__nand2_1
X_10080_ _10080_/A _10080_/B vssd1 vssd1 vccd1 vccd1 _10087_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_52_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10416_ _10416_/A vssd1 vssd1 vccd1 vccd1 _10417_/A sky130_fd_sc_hd__inv_2
XFILLER_0_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10347_ _10347_/A _10347_/B vssd1 vssd1 vccd1 vccd1 _10376_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10278_ _10278_/A _10278_/B vssd1 vssd1 vccd1 vccd1 _10279_/B sky130_fd_sc_hd__nand2_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06440_ _06440_/A _06440_/B _06440_/C vssd1 vssd1 vccd1 vccd1 _06616_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_61_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06371_ _06504_/C vssd1 vssd1 vccd1 vccd1 _06372_/B sky130_fd_sc_hd__inv_2
X_09090_ input51/X _10284_/B vssd1 vssd1 vccd1 vccd1 _09091_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07787__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08110_ _08120_/A _08119_/B vssd1 vssd1 vccd1 vccd1 _08118_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_28_176 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08041_ _08041_/A _08041_/B _08041_/C vssd1 vssd1 vccd1 vccd1 _08043_/B sky130_fd_sc_hd__nand3_1
X_09992_ _09992_/A _09992_/B vssd1 vssd1 vccd1 vccd1 _09995_/A sky130_fd_sc_hd__nand2_1
X_08943_ _08943_/A _09129_/A vssd1 vssd1 vccd1 vccd1 _08946_/B sky130_fd_sc_hd__nand2_1
X_08874_ _08874_/A _08874_/B vssd1 vssd1 vccd1 vccd1 _08876_/A sky130_fd_sc_hd__nand2_1
X_07825_ _07825_/A _07825_/B _07825_/C vssd1 vssd1 vccd1 vccd1 _08066_/C sky130_fd_sc_hd__nand3_1
X_07756_ _07756_/A _08337_/A vssd1 vssd1 vccd1 vccd1 _07759_/B sky130_fd_sc_hd__nand2_1
XANTENNA__05770__A input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06707_ _06708_/B _06708_/A vssd1 vssd1 vccd1 vccd1 _06707_/Y sky130_fd_sc_hd__nand2_1
X_09426_ _10151_/A _10150_/A _09602_/B _09922_/B vssd1 vssd1 vccd1 vccd1 _09426_/X
+ sky130_fd_sc_hd__and4_1
X_07687_ _07687_/A _07687_/B _07687_/C vssd1 vssd1 vccd1 vccd1 _07688_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06638_ _06638_/A vssd1 vssd1 vccd1 vccd1 _06641_/A sky130_fd_sc_hd__inv_2
X_09357_ _10361_/B _09357_/B vssd1 vssd1 vccd1 vccd1 _09358_/B sky130_fd_sc_hd__nor2_1
X_06569_ _06569_/A _06569_/B vssd1 vssd1 vccd1 vccd1 _06572_/A sky130_fd_sc_hd__nand2_1
X_09288_ _09288_/A vssd1 vssd1 vccd1 vccd1 _09289_/B sky130_fd_sc_hd__inv_2
XFILLER_0_62_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08308_ _08308_/A vssd1 vssd1 vccd1 vccd1 _08351_/A sky130_fd_sc_hd__inv_2
XFILLER_0_62_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08239_ _08239_/A _08373_/B vssd1 vssd1 vccd1 vccd1 _08240_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10201_ _10201_/A _10201_/B vssd1 vssd1 vccd1 vccd1 _10205_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10132_ _10132_/A _10132_/B vssd1 vssd1 vccd1 vccd1 _10134_/A sky130_fd_sc_hd__xnor2_1
X_10063_ _10063_/A vssd1 vssd1 vccd1 vccd1 _10064_/A sky130_fd_sc_hd__inv_2
XFILLER_0_57_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__05574__B input38/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05940_ _10130_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _05942_/B sky130_fd_sc_hd__nand2_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05871_ _09778_/D _10187_/B vssd1 vssd1 vccd1 vccd1 _06200_/B sky130_fd_sc_hd__nand2_1
X_08590_ _10101_/A _10157_/B vssd1 vssd1 vccd1 vccd1 _08592_/A sky130_fd_sc_hd__nand2_1
X_07610_ _07540_/Y _07663_/B _07550_/Y vssd1 vssd1 vccd1 vccd1 _07613_/B sky130_fd_sc_hd__a21o_1
X_07541_ _07545_/C vssd1 vssd1 vccd1 vccd1 _07544_/B sky130_fd_sc_hd__inv_2
XFILLER_0_72_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07472_ _07697_/C _07472_/B vssd1 vssd1 vccd1 vccd1 _07546_/A sky130_fd_sc_hd__nand2_2
XFILLER_0_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09211_ _09209_/Y _08619_/B _09210_/Y vssd1 vssd1 vccd1 vccd1 _09214_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_8_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06423_ _06605_/B _06423_/B vssd1 vssd1 vccd1 vccd1 _06424_/B sky130_fd_sc_hd__nand2_1
X_06354_ _06549_/C _06549_/B _06353_/Y vssd1 vssd1 vccd1 vccd1 _06365_/A sky130_fd_sc_hd__a21oi_2
X_09142_ _09142_/A _09142_/B vssd1 vssd1 vccd1 vccd1 _09145_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_71_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08406__A _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09073_ _09336_/B _09336_/C vssd1 vssd1 vccd1 vccd1 _09335_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06285_ _06285_/A _06285_/B vssd1 vssd1 vccd1 vccd1 _06432_/C sky130_fd_sc_hd__nand2_1
X_08024_ _08024_/A _08032_/B _08024_/C vssd1 vssd1 vccd1 vccd1 _08025_/B sky130_fd_sc_hd__nand3_1
X_09975_ _09976_/B _09976_/A vssd1 vssd1 vccd1 vccd1 _10127_/A sky130_fd_sc_hd__or2_1
X_08926_ _08942_/A _08942_/C vssd1 vssd1 vccd1 vccd1 _08941_/A sky130_fd_sc_hd__nand2_1
X_08857_ _08859_/B vssd1 vssd1 vccd1 vccd1 _08858_/B sky130_fd_sc_hd__inv_2
X_07808_ _07808_/A _07875_/A vssd1 vssd1 vccd1 vccd1 _07809_/B sky130_fd_sc_hd__nand2_1
X_08788_ _10248_/D _10202_/C _08786_/C vssd1 vssd1 vccd1 vccd1 _08789_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_79_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07739_ _07739_/A _07739_/B vssd1 vssd1 vccd1 vccd1 _07768_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_1_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_219 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09409_ _09409_/A _09409_/B vssd1 vssd1 vccd1 vccd1 _09410_/B sky130_fd_sc_hd__and2_1
X_10681_ _10681_/A _10681_/B vssd1 vssd1 vccd1 vccd1 _10683_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07220__A _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09623__B1 _10108_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05659__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09147__A _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10115_ _10115_/A input24/X vssd1 vssd1 vccd1 vccd1 _10115_/Y sky130_fd_sc_hd__nand2_1
X_10046_ _10046_/A _10047_/A vssd1 vssd1 vccd1 vccd1 _10049_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_38_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06070_ _06070_/A _06070_/B vssd1 vssd1 vccd1 vccd1 _06072_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _09859_/B _09761_/C _09761_/B vssd1 vssd1 vccd1 vccd1 _09762_/A sky130_fd_sc_hd__a21o_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ _06976_/B _06973_/A vssd1 vssd1 vccd1 vccd1 _06975_/A sky130_fd_sc_hd__nand2_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _09287_/B _08714_/A _08714_/B vssd1 vssd1 vccd1 vccd1 _08754_/A sky130_fd_sc_hd__nand3_1
X_09691_ _09691_/A _10022_/A vssd1 vssd1 vccd1 vccd1 _10059_/A sky130_fd_sc_hd__nand2_1
X_05923_ _05923_/A vssd1 vssd1 vccd1 vccd1 _06755_/B sky130_fd_sc_hd__inv_2
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08642_ _08642_/A _08642_/B vssd1 vssd1 vccd1 vccd1 _08654_/B sky130_fd_sc_hd__nand2_1
X_05854_ _05854_/A vssd1 vssd1 vccd1 vccd1 _05855_/B sky130_fd_sc_hd__inv_2
X_05785_ _05785_/A _05785_/B vssd1 vssd1 vccd1 vccd1 _06040_/B sky130_fd_sc_hd__nand2_1
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ _08573_/A input17/X vssd1 vssd1 vccd1 vccd1 _08576_/A sky130_fd_sc_hd__nand2_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07524_ _07670_/A _07671_/A vssd1 vssd1 vccd1 vccd1 _07682_/C sky130_fd_sc_hd__nand2_1
X_07455_ _08725_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _07530_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06863__B _09698_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07959__B _08059_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06406_ _06570_/C vssd1 vssd1 vccd1 vccd1 _06569_/B sky130_fd_sc_hd__inv_2
XANTENNA__09605__B1 _10150_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07386_ _07448_/A _07449_/C vssd1 vssd1 vccd1 vccd1 _07396_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ _09125_/A _09125_/B vssd1 vssd1 vccd1 vccd1 _09130_/A sky130_fd_sc_hd__nand2_1
X_06337_ _06507_/B vssd1 vssd1 vccd1 vccd1 _06506_/A sky130_fd_sc_hd__inv_2
X_09056_ _09056_/A _09056_/B _09056_/C vssd1 vssd1 vccd1 vccd1 _09059_/C sky130_fd_sc_hd__nand3_1
X_06268_ _06268_/A _06268_/B _06268_/C vssd1 vssd1 vccd1 vccd1 _06431_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_32_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08007_ _08109_/B _08120_/B _08107_/A vssd1 vssd1 vccd1 vccd1 _08009_/A sky130_fd_sc_hd__a21oi_1
X_06199_ _06199_/A _06199_/B vssd1 vssd1 vccd1 vccd1 _06200_/A sky130_fd_sc_hd__nand2_1
X_09958_ _09958_/A _09958_/B vssd1 vssd1 vccd1 vccd1 _09959_/A sky130_fd_sc_hd__xnor2_1
X_08909_ _08913_/A _09111_/B vssd1 vssd1 vccd1 vccd1 _08912_/A sky130_fd_sc_hd__nand2_1
X_09889_ _09888_/B _09889_/B _09889_/C vssd1 vssd1 vccd1 vccd1 _10331_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__09414__B _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10733_ _10733_/CLK hold9/X fanout98/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__dfrtp_1
X_10664_ _10664_/A _10664_/B vssd1 vssd1 vccd1 vccd1 _10668_/A sky130_fd_sc_hd__nand2_1
X_10595_ _10595_/A _10603_/C vssd1 vssd1 vccd1 vccd1 _10605_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xoutput82 hold65/A vssd1 vssd1 vccd1 vccd1 y_o[24] sky130_fd_sc_hd__buf_12
Xoutput93 hold60/A vssd1 vssd1 vccd1 vccd1 y_o[5] sky130_fd_sc_hd__buf_12
Xoutput71 hold28/A vssd1 vssd1 vccd1 vccd1 y_o[14] sky130_fd_sc_hd__buf_12
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10029_ _10206_/B _10029_/B vssd1 vssd1 vccd1 vccd1 _10032_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05570_ _05570_/A vssd1 vssd1 vccd1 vccd1 _05577_/A sky130_fd_sc_hd__inv_2
XFILLER_0_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07240_ _07200_/Y _07300_/B _07239_/Y vssd1 vssd1 vccd1 vccd1 _07287_/A sky130_fd_sc_hd__a21oi_1
X_07171_ _07156_/Y _07314_/B _07170_/Y vssd1 vssd1 vccd1 vccd1 _07303_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06122_ _06122_/A _06122_/B _06122_/C vssd1 vssd1 vccd1 vccd1 _06234_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_5_179 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06053_ _08112_/A _10201_/B vssd1 vssd1 vccd1 vccd1 _06054_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06204__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09812_ _09812_/A _09812_/B vssd1 vssd1 vccd1 vccd1 _09819_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07019__B _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09743_ _09808_/B _09836_/B vssd1 vssd1 vccd1 vccd1 _09806_/A sky130_fd_sc_hd__nand2_1
XANTENNA__06858__B _10210_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06955_ _06955_/A _06955_/B _06955_/C vssd1 vssd1 vccd1 vccd1 _07113_/C sky130_fd_sc_hd__nand3_1
X_09674_ _09737_/B _10070_/B vssd1 vssd1 vccd1 vccd1 _09735_/A sky130_fd_sc_hd__nand2_1
X_06886_ _06888_/C vssd1 vssd1 vccd1 vccd1 _06887_/B sky130_fd_sc_hd__inv_2
X_05906_ _05906_/A _05906_/B vssd1 vssd1 vccd1 vccd1 _05911_/C sky130_fd_sc_hd__nand2_1
X_08625_ _08625_/A _09185_/A vssd1 vssd1 vccd1 vccd1 _08627_/A sky130_fd_sc_hd__nand2_1
X_05837_ _05843_/B _05843_/C vssd1 vssd1 vccd1 vccd1 _05842_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_49_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08556_ _08556_/A _08556_/B _08556_/C vssd1 vssd1 vccd1 vccd1 _08559_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_49_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05768_ input39/X vssd1 vssd1 vccd1 vccd1 _09678_/C sky130_fd_sc_hd__clkbuf_8
XFILLER_0_49_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07507_ _07509_/A vssd1 vssd1 vccd1 vccd1 _07508_/B sky130_fd_sc_hd__inv_2
XFILLER_0_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08487_ _08488_/B _08488_/A vssd1 vssd1 vccd1 vccd1 _08489_/A sky130_fd_sc_hd__or2_1
XFILLER_0_9_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_05699_ _06259_/A _06258_/A vssd1 vssd1 vccd1 vccd1 _05699_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07438_ _07442_/A _07442_/B vssd1 vssd1 vccd1 vccd1 _07439_/A sky130_fd_sc_hd__nand2_1
X_07369_ _07368_/B _07369_/B _07369_/C vssd1 vssd1 vccd1 vccd1 _07370_/B sky130_fd_sc_hd__nand3b_1
XFILLER_0_17_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09108_ _09108_/A _09108_/B vssd1 vssd1 vccd1 vccd1 _09109_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_72_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10380_ _10380_/A vssd1 vssd1 vccd1 vccd1 _10701_/B sky130_fd_sc_hd__inv_2
X_09039_ _09055_/A _09056_/A vssd1 vssd1 vccd1 vccd1 _09039_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_4_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08313__B _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10719__RESET_B fanout99/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10716_ _10718_/CLK _10716_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10647_ _10647_/A vssd1 vssd1 vccd1 vccd1 _10713_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10578_ _10603_/A _10578_/B vssd1 vssd1 vccd1 vccd1 hold53/A sky130_fd_sc_hd__xor2_1
XFILLER_0_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05863__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_36 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06740_ _06740_/A _06740_/B vssd1 vssd1 vccd1 vccd1 _06768_/B sky130_fd_sc_hd__nand2_1
X_06671_ _06671_/A vssd1 vssd1 vccd1 vccd1 _06671_/Y sky130_fd_sc_hd__inv_2
X_08410_ _10156_/A _10187_/A vssd1 vssd1 vccd1 vccd1 _08412_/A sky130_fd_sc_hd__nand2_1
X_05622_ _05622_/A _06078_/B vssd1 vssd1 vccd1 vccd1 _05625_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09390_ _09390_/A _09390_/B vssd1 vssd1 vccd1 vccd1 _09391_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05553_ _05553_/A _05553_/B vssd1 vssd1 vccd1 vccd1 _05560_/A sky130_fd_sc_hd__nand2_1
X_08341_ _08341_/A _08341_/B vssd1 vssd1 vccd1 vccd1 _08342_/C sky130_fd_sc_hd__nand2_1
X_08272_ _08272_/A _08272_/B vssd1 vssd1 vccd1 vccd1 _08320_/A sky130_fd_sc_hd__xor2_1
X_05484_ input14/X vssd1 vssd1 vccd1 vccd1 _10157_/B sky130_fd_sc_hd__clkbuf_4
X_07223_ _07377_/C _07377_/B _07222_/Y vssd1 vssd1 vccd1 vccd1 _07233_/A sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07154_ _07319_/A _07320_/B vssd1 vssd1 vccd1 vccd1 _07154_/Y sky130_fd_sc_hd__nor2_1
X_06105_ _06308_/B _06308_/C vssd1 vssd1 vccd1 vccd1 _06705_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07085_ _07106_/B _07100_/C vssd1 vssd1 vccd1 vccd1 _07099_/A sky130_fd_sc_hd__nand2_1
X_06036_ _06846_/A vssd1 vssd1 vccd1 vccd1 _06037_/B sky130_fd_sc_hd__inv_2
X_07987_ _07991_/A _07991_/C vssd1 vssd1 vccd1 vccd1 _07989_/A sky130_fd_sc_hd__nand2_1
X_09726_ _09724_/Y _09442_/B _09725_/Y vssd1 vssd1 vccd1 vccd1 _09896_/A sky130_fd_sc_hd__a21oi_2
X_06938_ _06938_/A _06938_/B _06938_/C vssd1 vssd1 vccd1 vccd1 _06941_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_69_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06869_ _06869_/A _06869_/B vssd1 vssd1 vccd1 vccd1 _06873_/A sky130_fd_sc_hd__nand2_1
X_09657_ _09932_/B _09658_/C _09658_/B vssd1 vssd1 vccd1 vccd1 _09659_/A sky130_fd_sc_hd__a21o_1
X_09588_ _09588_/A _09588_/B _09831_/A vssd1 vssd1 vccd1 vccd1 _10353_/C sky130_fd_sc_hd__nand3_2
X_08608_ _10130_/A _10156_/B vssd1 vssd1 vccd1 vccd1 _08609_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08539_ _08539_/A _08604_/A _08630_/A vssd1 vssd1 vccd1 vccd1 _08543_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_64_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10501_ _10652_/A _10499_/Y _10652_/B vssd1 vssd1 vccd1 vccd1 _10502_/B sky130_fd_sc_hd__a21boi_1
X_10432_ _10435_/A _10435_/B vssd1 vssd1 vccd1 vccd1 _10434_/A sky130_fd_sc_hd__nand2_1
X_10363_ _10560_/B _10365_/C vssd1 vssd1 vccd1 vccd1 _10364_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_236 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10294_ _10293_/B _10294_/B _10294_/C vssd1 vssd1 vccd1 vccd1 _10295_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__06779__A _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09602__B _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_494 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08890_ _09082_/B _08890_/B vssd1 vssd1 vccd1 vccd1 _08959_/A sky130_fd_sc_hd__nand2_1
X_07910_ _07910_/A _07910_/B vssd1 vssd1 vccd1 vccd1 _07938_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07841_ _08384_/B _08384_/A vssd1 vssd1 vccd1 vccd1 _07844_/A sky130_fd_sc_hd__nand2_1
XANTENNA__08369__A_N _08366_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07772_ _07800_/B _07800_/C vssd1 vssd1 vccd1 vccd1 _07799_/A sky130_fd_sc_hd__nand2_1
X_09511_ _09514_/B _09739_/A vssd1 vssd1 vccd1 vccd1 _09513_/A sky130_fd_sc_hd__nand2_1
XANTENNA__10004__A _10004_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06723_ _08432_/B _06723_/B _06723_/C vssd1 vssd1 vccd1 vccd1 _08432_/A sky130_fd_sc_hd__nand3_1
X_09442_ _09442_/A _09442_/B vssd1 vssd1 vccd1 vccd1 _09444_/A sky130_fd_sc_hd__nand2_1
X_06654_ _06654_/A _06660_/A vssd1 vssd1 vccd1 vccd1 _06965_/C sky130_fd_sc_hd__nand2_1
X_05605_ _05620_/A _05620_/B vssd1 vssd1 vccd1 vccd1 _05619_/A sky130_fd_sc_hd__nand2_1
X_09373_ _09393_/A _09373_/B _09373_/C vssd1 vssd1 vccd1 vccd1 _09373_/Y sky130_fd_sc_hd__nor3_1
X_06585_ _06590_/A vssd1 vssd1 vccd1 vccd1 _06589_/A sky130_fd_sc_hd__inv_2
XFILLER_0_74_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08324_ _08324_/A _08324_/B vssd1 vssd1 vccd1 vccd1 _08325_/B sky130_fd_sc_hd__nand2_1
X_05536_ _05422_/Y _05638_/B _05461_/Y vssd1 vssd1 vccd1 vccd1 _05892_/A sky130_fd_sc_hd__a21oi_2
XFILLER_0_74_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08255_ _08255_/A _08255_/B vssd1 vssd1 vccd1 vccd1 _08266_/B sky130_fd_sc_hd__xor2_1
X_05467_ _05913_/A vssd1 vssd1 vccd1 vccd1 _05471_/A sky130_fd_sc_hd__inv_2
XFILLER_0_61_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__05768__A input39/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08186_ _08186_/A _08197_/A vssd1 vssd1 vccd1 vccd1 _08195_/A sky130_fd_sc_hd__nand2_1
X_07206_ _07206_/A _07206_/B vssd1 vssd1 vccd1 vccd1 _07207_/B sky130_fd_sc_hd__nand2_1
X_05398_ _08573_/A _09922_/B vssd1 vssd1 vccd1 vccd1 _05680_/A sky130_fd_sc_hd__nand2_1
X_07137_ _07137_/A _07137_/B vssd1 vssd1 vccd1 vccd1 _07139_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07983__A _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07068_ _07067_/B _07068_/B _07068_/C vssd1 vssd1 vccd1 vccd1 _07069_/B sky130_fd_sc_hd__nand3b_1
X_06019_ _05800_/A _05802_/B _05843_/B vssd1 vssd1 vccd1 vccd1 _06085_/B sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09709_ _09718_/A _09718_/C vssd1 vssd1 vccd1 vccd1 _09716_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_37_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10734__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10415_ _10415_/A _10415_/B vssd1 vssd1 vccd1 vccd1 _10416_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07893__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10346_ _10348_/C vssd1 vssd1 vccd1 vccd1 _10347_/B sky130_fd_sc_hd__inv_2
X_10277_ input52/X _09840_/B input53/X _09749_/B vssd1 vssd1 vccd1 vccd1 _10278_/B
+ sky130_fd_sc_hd__a22o_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06370_ _06370_/A _06370_/B vssd1 vssd1 vccd1 vccd1 _06504_/C sky130_fd_sc_hd__nand2_1
XANTENNA__07787__B _07891_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08040_ _08040_/A _08040_/B vssd1 vssd1 vccd1 vccd1 _08043_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05588__A input64/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08899__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09991_ _09993_/B vssd1 vssd1 vccd1 vccd1 _09992_/B sky130_fd_sc_hd__inv_2
X_08942_ _08942_/A _08942_/B _08942_/C vssd1 vssd1 vccd1 vccd1 _09129_/A sky130_fd_sc_hd__nand3_1
X_08873_ _08875_/B _08875_/C vssd1 vssd1 vccd1 vccd1 _08874_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07824_ _07824_/A vssd1 vssd1 vccd1 vccd1 _07825_/C sky130_fd_sc_hd__inv_2
X_07755_ _07759_/A vssd1 vssd1 vccd1 vccd1 _07758_/A sky130_fd_sc_hd__inv_2
X_06706_ _06704_/Y _06310_/B _06705_/Y vssd1 vssd1 vccd1 vccd1 _06929_/A sky130_fd_sc_hd__a21o_1
X_07686_ _07686_/A _07686_/B vssd1 vssd1 vccd1 vccd1 _07688_/A sky130_fd_sc_hd__nand2_1
X_09425_ _09615_/B _09434_/C vssd1 vssd1 vccd1 vccd1 _09433_/A sky130_fd_sc_hd__nand2_1
X_06637_ _06641_/B _06638_/A vssd1 vssd1 vccd1 vccd1 _06640_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_35_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09356_ _09353_/Y _09354_/Y _09355_/Y vssd1 vssd1 vccd1 vccd1 _10361_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06568_ _06570_/A _06570_/B vssd1 vssd1 vccd1 vccd1 _06569_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_74_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09287_ _09287_/A _09287_/B vssd1 vssd1 vccd1 vccd1 _09289_/A sky130_fd_sc_hd__nor2_1
X_08307_ _10284_/B _10115_/A vssd1 vssd1 vccd1 vccd1 _08308_/A sky130_fd_sc_hd__nand2_1
X_05519_ _05384_/C _05384_/B _05518_/Y vssd1 vssd1 vccd1 vccd1 _06001_/A sky130_fd_sc_hd__a21oi_4
XFILLER_0_34_103 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06499_ _06499_/A _06696_/A _06696_/B vssd1 vssd1 vccd1 vccd1 _07274_/A sky130_fd_sc_hd__nand3_2
X_08238_ _08238_/A _08238_/B vssd1 vssd1 vccd1 vccd1 _08239_/A sky130_fd_sc_hd__nand2_1
X_10200_ _10220_/A _10220_/C vssd1 vssd1 vccd1 vccd1 _10219_/A sky130_fd_sc_hd__nand2_1
X_08169_ _08169_/A _08169_/B vssd1 vssd1 vccd1 vccd1 _08180_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_30_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10131_ _10131_/A _10131_/B vssd1 vssd1 vccd1 vccd1 _10132_/B sky130_fd_sc_hd__xnor2_1
X_10062_ _10062_/A _10063_/A vssd1 vssd1 vccd1 vccd1 _10065_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07218__A _09840_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10329_ _10329_/A _10329_/B _10329_/C vssd1 vssd1 vccd1 vccd1 _10332_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_21_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_05870_ _06185_/A _06186_/C vssd1 vssd1 vccd1 vccd1 _05870_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__05871__A _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07540_ _07661_/A _07656_/A vssd1 vssd1 vccd1 vccd1 _07540_/Y sky130_fd_sc_hd__nand2_1
X_07471_ _07472_/B _07471_/B _07471_/C vssd1 vssd1 vccd1 vccd1 _07697_/C sky130_fd_sc_hd__nand3_1
X_09210_ _09210_/A _09210_/B vssd1 vssd1 vccd1 vccd1 _09210_/Y sky130_fd_sc_hd__nor2_1
X_06422_ _06423_/B _06422_/B _06422_/C vssd1 vssd1 vccd1 vccd1 _06605_/B sky130_fd_sc_hd__nand3_1
X_06353_ _06546_/B _06545_/A vssd1 vssd1 vccd1 vccd1 _06353_/Y sky130_fd_sc_hd__nor2_1
X_09141_ _09142_/B _09142_/A vssd1 vssd1 vccd1 vccd1 _09145_/B sky130_fd_sc_hd__or2_1
X_09072_ _09071_/B _09072_/B _09072_/C vssd1 vssd1 vccd1 vccd1 _09336_/C sky130_fd_sc_hd__nand3b_1
XANTENNA__08406__B _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08023_ _08032_/A _08129_/A vssd1 vssd1 vccd1 vccd1 _08025_/A sky130_fd_sc_hd__nand2_1
X_06284_ _06284_/A _06284_/B _06284_/C vssd1 vssd1 vccd1 vccd1 _06285_/B sky130_fd_sc_hd__nand3_1
XANTENNA__06207__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09974_ _10127_/B _09974_/B vssd1 vssd1 vccd1 vccd1 _09976_/A sky130_fd_sc_hd__nand2_1
X_08925_ _08916_/Y _08925_/B _08925_/C vssd1 vssd1 vccd1 vccd1 _08942_/C sky130_fd_sc_hd__nand3b_1
X_08856_ _08856_/A _08856_/B vssd1 vssd1 vccd1 vccd1 _08859_/B sky130_fd_sc_hd__xor2_1
XANTENNA__09253__A _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__05781__A _08739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ _07797_/A _07796_/A _07797_/B vssd1 vssd1 vccd1 vccd1 _07811_/B sky130_fd_sc_hd__a21boi_2
X_08787_ _08787_/A vssd1 vssd1 vccd1 vccd1 _08790_/B sky130_fd_sc_hd__inv_2
X_05999_ _06005_/B _06810_/A vssd1 vssd1 vccd1 vccd1 _06884_/B sky130_fd_sc_hd__nand2_1
X_07738_ _07744_/B vssd1 vssd1 vccd1 vccd1 _07739_/B sky130_fd_sc_hd__inv_2
X_07669_ _07669_/A _07669_/B vssd1 vssd1 vccd1 vccd1 _07735_/A sky130_fd_sc_hd__nand2_1
X_09408_ _09411_/B _09620_/A vssd1 vssd1 vccd1 vccd1 _09410_/A sky130_fd_sc_hd__nand2_1
X_10680_ _10680_/A vssd1 vssd1 vccd1 vccd1 _10722_/D sky130_fd_sc_hd__clkbuf_1
X_09339_ _09339_/A _09339_/B vssd1 vssd1 vccd1 vccd1 _09340_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07220__B _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09623__A1 _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09387__B1 _10129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ _10108_/B input22/X _10113_/B vssd1 vssd1 vccd1 vccd1 _10117_/C sky130_fd_sc_hd__a21bo_1
X_10045_ _10045_/A _10045_/B vssd1 vssd1 vccd1 vccd1 _10047_/A sky130_fd_sc_hd__xor2_1
XANTENNA__09163__A _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold60 hold60/A vssd1 vssd1 vccd1 vccd1 hold60/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__05866__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ _06974_/B vssd1 vssd1 vccd1 vccd1 _06976_/B sky130_fd_sc_hd__inv_2
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _08710_/A _08710_/B vssd1 vssd1 vccd1 vccd1 _08714_/B sky130_fd_sc_hd__nand2_1
X_09690_ _10022_/B _09690_/B _09690_/C vssd1 vssd1 vccd1 vccd1 _10022_/A sky130_fd_sc_hd__nand3_1
X_05922_ _05924_/A _05924_/B vssd1 vssd1 vccd1 vccd1 _05923_/A sky130_fd_sc_hd__nor2_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08641_ _08413_/C _08413_/B _08407_/Y vssd1 vssd1 vccd1 vccd1 _08642_/B sky130_fd_sc_hd__a21oi_1
X_05853_ _05853_/A _05854_/A _05853_/C vssd1 vssd1 vccd1 vccd1 _05857_/B sky130_fd_sc_hd__nand3_1
X_05784_ _05786_/B vssd1 vssd1 vccd1 vccd1 _05785_/B sky130_fd_sc_hd__inv_2
XFILLER_0_49_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08572_ _10115_/A input18/X vssd1 vssd1 vccd1 vccd1 _08579_/B sky130_fd_sc_hd__nand2_1
X_07523_ _08724_/A input55/X vssd1 vssd1 vccd1 vccd1 _07671_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07454_ _07545_/A _07545_/B vssd1 vssd1 vccd1 vccd1 _07544_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06405_ _10292_/B _09477_/C vssd1 vssd1 vccd1 vccd1 _06570_/C sky130_fd_sc_hd__nand2_1
XANTENNA__09605__B2 _09922_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09605__A1 _10151_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07385_ _07482_/C _07482_/B _07384_/Y vssd1 vssd1 vccd1 vccd1 _07449_/C sky130_fd_sc_hd__a21oi_2
XFILLER_0_17_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09124_ _09126_/B _09564_/A vssd1 vssd1 vccd1 vccd1 _09125_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06336_ _07756_/A _07891_/B vssd1 vssd1 vccd1 vccd1 _06507_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_32_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09055_ _09055_/A _09055_/B vssd1 vssd1 vccd1 vccd1 _09059_/B sky130_fd_sc_hd__nand2_1
X_06267_ _06267_/A _06267_/B vssd1 vssd1 vccd1 vccd1 _06268_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08006_ _08006_/A _08006_/B vssd1 vssd1 vccd1 vccd1 _08107_/A sky130_fd_sc_hd__nor2_1
X_06198_ _06203_/B vssd1 vssd1 vccd1 vccd1 _06201_/A sky130_fd_sc_hd__inv_2
X_09957_ _09957_/A _09957_/B vssd1 vssd1 vccd1 vccd1 _09958_/B sky130_fd_sc_hd__nand2_1
X_08908_ _08907_/B _08908_/B _09101_/A vssd1 vssd1 vccd1 vccd1 _09111_/B sky130_fd_sc_hd__nand3b_1
X_09888_ _09888_/A _09888_/B vssd1 vssd1 vccd1 vccd1 _09890_/A sky130_fd_sc_hd__nand2_1
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08839_ _08839_/A _08839_/B vssd1 vssd1 vccd1 vccd1 _08978_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06400__A _09551_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10732_ _10733_/CLK hold16/X fanout98/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__dfrtp_2
XFILLER_0_82_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10663_ _10663_/A _10663_/B vssd1 vssd1 vccd1 vccd1 _10665_/A sky130_fd_sc_hd__nand2_1
X_10594_ _10594_/A vssd1 vssd1 vccd1 vccd1 _10603_/C sky130_fd_sc_hd__inv_2
XFILLER_0_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05686__A _08573_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08062__A _08218_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput83 hold17/A vssd1 vssd1 vccd1 vccd1 y_o[25] sky130_fd_sc_hd__buf_12
Xoutput72 _10725_/Q vssd1 vssd1 vccd1 vccd1 y_o[15] sky130_fd_sc_hd__buf_12
Xoutput94 hold33/A vssd1 vssd1 vccd1 vccd1 y_o[6] sky130_fd_sc_hd__buf_12
X_10028_ _10201_/A _09698_/A _09677_/A _09477_/C vssd1 vssd1 vccd1 vccd1 _10029_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_68 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09621__A _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07170_ _07312_/A _07311_/A vssd1 vssd1 vccd1 vccd1 _07170_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__06980__A _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06121_ _06121_/A _06121_/B _06121_/C vssd1 vssd1 vccd1 vccd1 _06122_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06052_ _06869_/B _06055_/C vssd1 vssd1 vccd1 vccd1 _06054_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06204__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09811_ _09813_/A vssd1 vssd1 vccd1 vccd1 _09812_/B sky130_fd_sc_hd__inv_2
X_09742_ _09742_/A _09742_/B _10070_/A vssd1 vssd1 vccd1 vccd1 _09836_/B sky130_fd_sc_hd__nand3_2
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06858__C _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06954_ _06954_/A _06954_/B _06954_/C vssd1 vssd1 vccd1 vccd1 _06955_/B sky130_fd_sc_hd__nand3_1
X_09673_ _09673_/A _09998_/A _09673_/C vssd1 vssd1 vccd1 vccd1 _10070_/B sky130_fd_sc_hd__nand3_2
X_06885_ _06883_/Y _06008_/B _06884_/Y vssd1 vssd1 vccd1 vccd1 _06888_/C sky130_fd_sc_hd__a21oi_2
X_05905_ _05905_/A _05905_/B vssd1 vssd1 vccd1 vccd1 _06734_/B sky130_fd_sc_hd__nand2_1
X_08624_ _08624_/A _08625_/A _09185_/A vssd1 vssd1 vccd1 vccd1 _09134_/B sky130_fd_sc_hd__nand3_2
X_05836_ _05836_/A _05836_/B _05836_/C vssd1 vssd1 vccd1 vccd1 _05843_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_27_91 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08555_ _08555_/A _08555_/B vssd1 vssd1 vccd1 vccd1 _08559_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_49_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05767_ _08112_/A _10187_/B vssd1 vssd1 vccd1 vccd1 _05861_/B sky130_fd_sc_hd__nand2_1
X_07506_ _07614_/B _07614_/C vssd1 vssd1 vccd1 vccd1 _07613_/A sky130_fd_sc_hd__nand2_1
X_08486_ _08486_/A _08486_/B vssd1 vssd1 vccd1 vccd1 _08488_/A sky130_fd_sc_hd__nand2_1
X_05698_ _06260_/C vssd1 vssd1 vccd1 vccd1 _06243_/C sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07437_ _07437_/A _07437_/B vssd1 vssd1 vccd1 vccd1 _07442_/B sky130_fd_sc_hd__nand2_1
X_07368_ _07368_/A _07368_/B vssd1 vssd1 vccd1 vccd1 _07370_/A sky130_fd_sc_hd__nand2_1
X_09107_ _09107_/A _09108_/B _09108_/A vssd1 vssd1 vccd1 vccd1 _09544_/B sky130_fd_sc_hd__nand3_2
XFILLER_0_72_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06319_ _06688_/B _06688_/C vssd1 vssd1 vccd1 vccd1 _06690_/B sky130_fd_sc_hd__nand2_1
X_07299_ _07301_/A _07301_/B vssd1 vssd1 vccd1 vccd1 _07300_/A sky130_fd_sc_hd__nand2_1
X_09038_ _09055_/B vssd1 vssd1 vccd1 vccd1 _09056_/A sky130_fd_sc_hd__inv_2
XANTENNA__06130__A _08101_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10715_ _10718_/CLK hold48/X fanout99/X vssd1 vssd1 vccd1 vccd1 hold60/A sky130_fd_sc_hd__dfrtp_1
X_10646_ _10646_/A _10646_/B vssd1 vssd1 vccd1 vccd1 _10647_/A sky130_fd_sc_hd__and2_1
X_10577_ _10708_/B _10580_/A vssd1 vssd1 vccd1 vccd1 _10578_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05863__B input37/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06670_ _06945_/A _06943_/A vssd1 vssd1 vccd1 vccd1 _06671_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_64_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05621_ _05623_/B _05623_/C vssd1 vssd1 vccd1 vccd1 _06078_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_73_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05552_ _05600_/B vssd1 vssd1 vccd1 vccd1 _05553_/B sky130_fd_sc_hd__inv_2
X_08340_ _09782_/B _10113_/A _08308_/A vssd1 vssd1 vccd1 vccd1 _08341_/B sky130_fd_sc_hd__o21ai_1
X_05483_ _05948_/A vssd1 vssd1 vccd1 vccd1 _05487_/A sky130_fd_sc_hd__inv_2
XFILLER_0_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08271_ _08195_/Y _08271_/B vssd1 vssd1 vccd1 vccd1 _08272_/B sky130_fd_sc_hd__nand2b_1
XFILLER_0_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07222_ _07222_/A _07222_/B vssd1 vssd1 vccd1 vccd1 _07222_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_54_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07153_ _07321_/C vssd1 vssd1 vccd1 vccd1 _07323_/B sky130_fd_sc_hd__inv_2
XFILLER_0_6_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06104_ _06104_/A _06104_/B _06104_/C vssd1 vssd1 vccd1 vccd1 _06308_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07084_ _07084_/A _07084_/B vssd1 vssd1 vccd1 vccd1 _07100_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06035_ _05616_/C _05616_/B _05610_/A vssd1 vssd1 vccd1 vccd1 _06846_/A sky130_fd_sc_hd__a21oi_2
X_07986_ _07986_/A _07986_/B vssd1 vssd1 vccd1 vccd1 _07991_/C sky130_fd_sc_hd__nand2_1
X_09725_ _09725_/A _09725_/B vssd1 vssd1 vccd1 vccd1 _09725_/Y sky130_fd_sc_hd__nor2_1
X_06937_ _06937_/A _06937_/B vssd1 vssd1 vccd1 vccd1 _10409_/A sky130_fd_sc_hd__nand2_2
X_09656_ _09388_/B _10128_/A _10156_/B _09386_/X vssd1 vssd1 vccd1 vccd1 _09658_/B
+ sky130_fd_sc_hd__a31o_1
X_06868_ _06870_/B _06870_/A vssd1 vssd1 vccd1 vccd1 _08842_/A sky130_fd_sc_hd__or2_1
X_08607_ _10129_/A _10151_/B vssd1 vssd1 vccd1 vccd1 _08609_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09587_ _09587_/A vssd1 vssd1 vccd1 vccd1 _09588_/B sky130_fd_sc_hd__inv_2
X_05819_ _09778_/D _09698_/A vssd1 vssd1 vccd1 vccd1 _05824_/A sky130_fd_sc_hd__nand2_1
X_06799_ _06799_/A _06799_/B vssd1 vssd1 vccd1 vccd1 _06801_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08538_ _08630_/B _08538_/B vssd1 vssd1 vccd1 vccd1 _08543_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_64_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08469_ _10115_/A _10128_/B vssd1 vssd1 vccd1 vccd1 _08476_/B sky130_fd_sc_hd__nand2_1
X_10500_ _10500_/A hold60/X _10500_/C vssd1 vssd1 vccd1 vccd1 _10652_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_64_178 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08605__A _10128_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10431_ _10438_/A _10431_/B _10431_/C vssd1 vssd1 vccd1 vccd1 _10435_/B sky130_fd_sc_hd__nand3_1
X_10362_ _10370_/B _10370_/A vssd1 vssd1 vccd1 vccd1 _10560_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_20_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10293_ _10293_/A _10293_/B vssd1 vssd1 vccd1 vccd1 _10295_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_20_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06779__B _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10629_ _10629_/A vssd1 vssd1 vccd1 vccd1 _10632_/C sky130_fd_sc_hd__inv_2
XFILLER_0_70_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_362 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05874__A _08112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07840_ _07850_/B _07843_/C vssd1 vssd1 vccd1 vccd1 _08384_/B sky130_fd_sc_hd__nand2_1
X_07771_ _07951_/B _07950_/B _07951_/A vssd1 vssd1 vccd1 vccd1 _07776_/A sky130_fd_sc_hd__a21boi_1
X_09510_ _09510_/A _09510_/B _09739_/B vssd1 vssd1 vccd1 vccd1 _09739_/A sky130_fd_sc_hd__nand3_2
XANTENNA__10004__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06722_ _06722_/A vssd1 vssd1 vccd1 vccd1 _06723_/B sky130_fd_sc_hd__inv_2
X_09441_ _09441_/A _09441_/B vssd1 vssd1 vccd1 vccd1 _09442_/B sky130_fd_sc_hd__nand2_1
X_06653_ _06660_/B _06653_/B _06653_/C vssd1 vssd1 vccd1 vccd1 _06660_/A sky130_fd_sc_hd__nand3_1
X_05604_ _05604_/A _05604_/B _05966_/A vssd1 vssd1 vccd1 vccd1 _05620_/B sky130_fd_sc_hd__nand3_1
X_09372_ _10103_/B input17/X vssd1 vssd1 vccd1 vccd1 _09373_/C sky130_fd_sc_hd__nand2_1
X_06584_ _10275_/B _10150_/A vssd1 vssd1 vccd1 vccd1 _06590_/A sky130_fd_sc_hd__nand2_1
X_05535_ _05631_/B _05631_/C vssd1 vssd1 vccd1 vccd1 _05892_/B sky130_fd_sc_hd__nand2_1
X_08323_ _08356_/A _08323_/B vssd1 vssd1 vccd1 vccd1 _08357_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08425__A _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08254_ _08162_/Y _08254_/B vssd1 vssd1 vccd1 vccd1 _08255_/B sky130_fd_sc_hd__nand2b_1
X_05466_ _05471_/B _05913_/A vssd1 vssd1 vccd1 vccd1 _05470_/A sky130_fd_sc_hd__nand2_1
X_07205_ _07205_/A _07205_/B vssd1 vssd1 vccd1 vccd1 _07207_/A sky130_fd_sc_hd__nand2_1
X_08185_ _08197_/B _08185_/B _08185_/C vssd1 vssd1 vccd1 vccd1 _08197_/A sky130_fd_sc_hd__nand3_1
X_05397_ _05673_/B _05673_/C vssd1 vssd1 vccd1 vccd1 _05672_/A sky130_fd_sc_hd__nand2_1
X_07136_ _07298_/B _07298_/C vssd1 vssd1 vccd1 vccd1 _07297_/A sky130_fd_sc_hd__nand2_1
XANTENNA__07983__B _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07067_ _07067_/A _07067_/B vssd1 vssd1 vccd1 vccd1 _07069_/A sky130_fd_sc_hd__nand2_1
X_06018_ _06089_/A _06089_/B vssd1 vssd1 vccd1 vccd1 _06088_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_2_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09256__A _10211_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08160__A _09749_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09708_ _10035_/A _09708_/B _09708_/C vssd1 vssd1 vccd1 vccd1 _09718_/C sky130_fd_sc_hd__nand3_1
X_07969_ _08069_/A _07971_/A _07971_/B vssd1 vssd1 vccd1 vccd1 _08225_/B sky130_fd_sc_hd__nand3_1
X_09639_ _09642_/A _09963_/A vssd1 vssd1 vccd1 vccd1 _09640_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_77_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09956__B1 _10103_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10414_ _10414_/A _10414_/B _10414_/C vssd1 vssd1 vccd1 vccd1 _10415_/B sky130_fd_sc_hd__nand3_1
X_10345_ _10345_/A vssd1 vssd1 vccd1 vccd1 _10603_/A sky130_fd_sc_hd__inv_2
XANTENNA__07893__B _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10276_ _10276_/A _10276_/B _10276_/C _10276_/D vssd1 vssd1 vccd1 vccd1 _10278_/A
+ sky130_fd_sc_hd__or4_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08899__B _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09990_ _09990_/A _09990_/B vssd1 vssd1 vccd1 vccd1 _09993_/B sky130_fd_sc_hd__nand2_1
X_08941_ _08941_/A _08941_/B vssd1 vssd1 vccd1 vccd1 _08943_/A sky130_fd_sc_hd__nand2_1
X_08872_ _08872_/A _08872_/B _08872_/C vssd1 vssd1 vccd1 vccd1 _08875_/C sky130_fd_sc_hd__nand3_1
X_07823_ _07823_/A _07823_/B vssd1 vssd1 vccd1 vccd1 _07825_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07754_ _08739_/A _08171_/B vssd1 vssd1 vccd1 vccd1 _07759_/A sky130_fd_sc_hd__nand2_1
X_06705_ _06705_/A _06705_/B vssd1 vssd1 vccd1 vccd1 _06705_/Y sky130_fd_sc_hd__nor2_1
X_07685_ _07687_/A _07687_/C vssd1 vssd1 vccd1 vccd1 _07686_/A sky130_fd_sc_hd__nand2_1
X_09424_ _09424_/A _09424_/B vssd1 vssd1 vccd1 vccd1 _09434_/C sky130_fd_sc_hd__nand2_1
X_06636_ _06639_/B vssd1 vssd1 vccd1 vccd1 _06641_/B sky130_fd_sc_hd__inv_2
XFILLER_0_59_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09355_ _09354_/B _09354_/C _09354_/A vssd1 vssd1 vccd1 vccd1 _09355_/Y sky130_fd_sc_hd__a21oi_1
X_06567_ _06567_/A _06567_/B _06567_/C vssd1 vssd1 vccd1 vccd1 _06570_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09286_ _09292_/A _09292_/B vssd1 vssd1 vccd1 vccd1 _09291_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_19_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08306_ _08312_/A _08312_/B vssd1 vssd1 vccd1 vccd1 _08311_/A sky130_fd_sc_hd__nand2_1
X_05518_ _05518_/A _05518_/B vssd1 vssd1 vccd1 vccd1 _05518_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06498_ _06497_/B _06498_/B _06498_/C vssd1 vssd1 vccd1 vccd1 _06696_/B sky130_fd_sc_hd__nand3b_1
X_08237_ _08375_/A _08235_/Y _08236_/Y vssd1 vssd1 vccd1 vccd1 _10487_/B sky130_fd_sc_hd__a21oi_1
X_05449_ _05449_/A _05449_/B vssd1 vssd1 vccd1 vccd1 _05650_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_42_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08168_ _08169_/A _08168_/B vssd1 vssd1 vccd1 vccd1 _08180_/A sky130_fd_sc_hd__nand2b_1
X_08099_ _08099_/A _08099_/B vssd1 vssd1 vccd1 vccd1 _08130_/B sky130_fd_sc_hd__nand2_1
X_07119_ _07427_/B _07427_/C vssd1 vssd1 vccd1 vccd1 _07426_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_30_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10130_ _10130_/A input18/X vssd1 vssd1 vccd1 vccd1 _10131_/B sky130_fd_sc_hd__nand2_1
X_10061_ _10061_/A _10061_/B vssd1 vssd1 vccd1 vccd1 _10063_/A sky130_fd_sc_hd__nor2_1
XANTENNA__09166__A1 _09971_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07218__B _10158_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10328_ _10328_/A _10328_/B vssd1 vssd1 vccd1 vccd1 _10332_/B sky130_fd_sc_hd__nand2_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ _10259_/A _10259_/B vssd1 vssd1 vccd1 vccd1 _10259_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__05871__B _10187_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07470_ _07620_/B _07621_/B vssd1 vssd1 vccd1 vccd1 _07471_/C sky130_fd_sc_hd__nand2_1
X_06421_ _06430_/B _06431_/C _06431_/B vssd1 vssd1 vccd1 vccd1 _06423_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_29_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06352_ _06547_/C vssd1 vssd1 vccd1 vccd1 _06549_/B sky130_fd_sc_hd__inv_2
X_09140_ _09140_/A _09140_/B vssd1 vssd1 vccd1 vccd1 _09142_/A sky130_fd_sc_hd__xor2_1
XFILLER_0_71_232 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09071_ _09071_/A _09071_/B vssd1 vssd1 vccd1 vccd1 _09336_/B sky130_fd_sc_hd__nand2_1
X_06283_ _06283_/A _06283_/B vssd1 vssd1 vccd1 vccd1 _06284_/A sky130_fd_sc_hd__nand2_1
X_08022_ _08032_/B vssd1 vssd1 vccd1 vccd1 _08129_/A sky130_fd_sc_hd__inv_2
XFILLER_0_21_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06207__B _09678_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09973_ _09971_/A _09971_/B _09971_/C vssd1 vssd1 vccd1 vccd1 _09974_/B sky130_fd_sc_hd__o21ai_1
X_08924_ _08924_/A _08928_/A vssd1 vssd1 vccd1 vccd1 _08942_/A sky130_fd_sc_hd__nand2_1
X_08855_ _08855_/A _08855_/B vssd1 vssd1 vccd1 vccd1 _08856_/B sky130_fd_sc_hd__nor2_1
XANTENNA__09253__B _10201_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08786_ _10248_/D _10202_/C _08786_/C vssd1 vssd1 vccd1 vccd1 _08787_/A sky130_fd_sc_hd__nor3_1
XANTENNA__05781__B input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ _07868_/B _07867_/A vssd1 vssd1 vccd1 vccd1 _07872_/C sky130_fd_sc_hd__nand2_1
X_05998_ _05997_/B _06810_/B _05998_/C vssd1 vssd1 vccd1 vccd1 _06810_/A sky130_fd_sc_hd__nand3b_1
X_07737_ _07737_/A _07737_/B vssd1 vssd1 vccd1 vccd1 _07868_/B sky130_fd_sc_hd__nand2_2
XFILLER_0_79_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07668_ _07668_/A _07668_/B _07668_/C vssd1 vssd1 vccd1 vccd1 _07669_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09407_ _09407_/A _09620_/B _09407_/C vssd1 vssd1 vccd1 vccd1 _09620_/A sky130_fd_sc_hd__nand3_1
X_07599_ _07599_/A _07599_/B vssd1 vssd1 vccd1 vccd1 _07600_/A sky130_fd_sc_hd__nand2_1
X_06619_ _06622_/B vssd1 vssd1 vccd1 vccd1 _06624_/B sky130_fd_sc_hd__inv_2
X_09338_ _09354_/A _09338_/B vssd1 vssd1 vccd1 vccd1 _10389_/B sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09269_ _09268_/A _10248_/D _09268_/C vssd1 vssd1 vccd1 vccd1 _09269_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_50_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09387__A1 _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09387__B2 _10157_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ _10113_/A _10113_/B input22/X vssd1 vssd1 vccd1 vccd1 _10117_/B sky130_fd_sc_hd__or3b_1
XFILLER_0_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10044_ _10044_/A _10043_/X vssd1 vssd1 vccd1 vccd1 _10045_/B sky130_fd_sc_hd__or2b_1
Xhold50 hold50/A vssd1 vssd1 vccd1 vccd1 hold50/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 hold61/A vssd1 vssd1 vccd1 vccd1 hold61/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05866__B _10148_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ _07127_/B _07127_/C vssd1 vssd1 vccd1 vccd1 _07132_/A sky130_fd_sc_hd__nand2_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05921_ _08337_/A _10158_/B vssd1 vssd1 vccd1 vccd1 _05924_/B sky130_fd_sc_hd__nand2_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08640_ _08643_/B _08643_/C vssd1 vssd1 vccd1 vccd1 _08642_/A sky130_fd_sc_hd__nand2_1
X_05852_ _06118_/C vssd1 vssd1 vccd1 vccd1 _06117_/B sky130_fd_sc_hd__inv_2
X_05783_ _07675_/A input39/X vssd1 vssd1 vccd1 vccd1 _05786_/B sky130_fd_sc_hd__nand2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08571_ _08571_/A _08571_/B vssd1 vssd1 vccd1 vccd1 _08580_/A sky130_fd_sc_hd__nand2_1
X_07522_ _08725_/A input58/X vssd1 vssd1 vccd1 vccd1 _07670_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07453_ _07453_/A _07453_/B vssd1 vssd1 vccd1 vccd1 _07545_/A sky130_fd_sc_hd__nand2_1
X_06404_ _08897_/B vssd1 vssd1 vccd1 vccd1 _10292_/B sky130_fd_sc_hd__buf_6
X_09123_ _09122_/B _09123_/B _09564_/B vssd1 vssd1 vccd1 vccd1 _09564_/A sky130_fd_sc_hd__nand3b_2
XANTENNA__09605__A2 _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07384_ _07384_/A _07384_/B vssd1 vssd1 vccd1 vccd1 _07384_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06335_ _06506_/B vssd1 vssd1 vccd1 vccd1 _06507_/A sky130_fd_sc_hd__inv_2
X_09054_ _09351_/A _09077_/C vssd1 vssd1 vccd1 vccd1 _09076_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_4_351 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06266_ _06266_/A _06266_/B _06266_/C vssd1 vssd1 vccd1 vccd1 _06431_/B sky130_fd_sc_hd__nand3_1
X_08005_ _08119_/B vssd1 vssd1 vccd1 vccd1 _08120_/B sky130_fd_sc_hd__inv_2
XANTENNA__07049__A _09517_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06197_ _06369_/C _06369_/B _06196_/Y vssd1 vssd1 vccd1 vccd1 _06203_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09956_ _10103_/A input24/X _10103_/B input19/X vssd1 vssd1 vccd1 vccd1 _09957_/B
+ sky130_fd_sc_hd__a22o_1
X_08907_ _08907_/A _08907_/B vssd1 vssd1 vccd1 vccd1 _08913_/A sky130_fd_sc_hd__nand2_1
X_09887_ _09889_/B _09889_/C vssd1 vssd1 vccd1 vccd1 _09888_/A sky130_fd_sc_hd__nand2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _08840_/C vssd1 vssd1 vccd1 vccd1 _08839_/B sky130_fd_sc_hd__inv_2
XANTENNA__06400__B _10188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08769_ _08769_/A _08769_/B vssd1 vssd1 vccd1 vccd1 _08832_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_79_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10731_ _10741_/CLK hold53/X fanout98/X vssd1 vssd1 vccd1 vccd1 hold52/A sky130_fd_sc_hd__dfrtp_2
XANTENNA__08608__A _10130_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10662_ _10664_/A vssd1 vssd1 vccd1 vccd1 _10663_/A sky130_fd_sc_hd__inv_2
XANTENNA__06128__A _08337_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10593_ _10596_/A _10694_/A _10593_/C vssd1 vssd1 vccd1 vccd1 _10597_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__05967__A _07646_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05686__B _09602_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__B2 _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09780__A1 input52/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput84 hold20/A vssd1 vssd1 vccd1 vccd1 y_o[26] sky130_fd_sc_hd__buf_12
Xoutput73 hold54/A vssd1 vssd1 vccd1 vccd1 y_o[16] sky130_fd_sc_hd__buf_12
Xoutput95 hold57/A vssd1 vssd1 vccd1 vccd1 y_o[7] sky130_fd_sc_hd__buf_12
X_10027_ _10027_/A _10202_/A _10202_/C _10202_/D vssd1 vssd1 vccd1 vccd1 _10206_/B
+ sky130_fd_sc_hd__or4_1
XFILLER_0_53_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06980__B _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06120_ _06120_/A _06120_/B vssd1 vssd1 vccd1 vccd1 _06122_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_41_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06051_ _10276_/B _10202_/C _06047_/Y vssd1 vssd1 vccd1 vccd1 _06055_/C sky130_fd_sc_hd__o21ai_1
XFILLER_0_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09810_ _09810_/A _09810_/B vssd1 vssd1 vccd1 vccd1 _09813_/A sky130_fd_sc_hd__nand2_1
X_09741_ _09741_/A _09741_/B vssd1 vssd1 vccd1 vccd1 _09808_/B sky130_fd_sc_hd__nand2_1
X_06953_ _06953_/A _06953_/B vssd1 vssd1 vccd1 vccd1 _06955_/A sky130_fd_sc_hd__nand2_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05904_ _05906_/B vssd1 vssd1 vccd1 vccd1 _05905_/B sky130_fd_sc_hd__inv_2
X_09672_ _09672_/A _09672_/B vssd1 vssd1 vccd1 vccd1 _09737_/B sky130_fd_sc_hd__nand2_1
X_06884_ _06884_/A _06884_/B vssd1 vssd1 vccd1 vccd1 _06884_/Y sky130_fd_sc_hd__nor2_1
X_08623_ _08623_/A _09185_/B _08623_/C vssd1 vssd1 vccd1 vccd1 _09185_/A sky130_fd_sc_hd__nand3_2
X_05835_ _05835_/A _05835_/B vssd1 vssd1 vccd1 vccd1 _05843_/B sky130_fd_sc_hd__nand2_1
X_08554_ _08554_/A _08554_/B vssd1 vssd1 vccd1 vccd1 _08878_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_05766_ input23/X vssd1 vssd1 vccd1 vccd1 _08112_/A sky130_fd_sc_hd__buf_6
XFILLER_0_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07505_ _07505_/A _07505_/B _07505_/C vssd1 vssd1 vccd1 vccd1 _07614_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_76_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05697_ _05697_/A _05697_/B vssd1 vssd1 vccd1 vccd1 _06260_/C sky130_fd_sc_hd__nand2_1
X_08485_ _08485_/A _08485_/B vssd1 vssd1 vccd1 vccd1 _08486_/B sky130_fd_sc_hd__nand2_1
X_07436_ _07713_/B _07436_/B vssd1 vssd1 vccd1 vccd1 _07437_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_17_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07367_ _07545_/B _07452_/A vssd1 vssd1 vccd1 vccd1 _07368_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_17_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ _09102_/A _09102_/B _09105_/Y vssd1 vssd1 vccd1 vccd1 _09108_/A sky130_fd_sc_hd__o21ai_2
XFILLER_0_72_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06318_ _06318_/A _06318_/B _06318_/C vssd1 vssd1 vccd1 vccd1 _06688_/C sky130_fd_sc_hd__nand3_1
X_09037_ _09037_/A _09037_/B vssd1 vssd1 vccd1 vccd1 _09055_/B sky130_fd_sc_hd__nand2_1
X_07298_ _07298_/A _07298_/B _07298_/C vssd1 vssd1 vccd1 vccd1 _07301_/B sky130_fd_sc_hd__nand3_1
X_06249_ _06413_/B _06413_/C vssd1 vssd1 vccd1 vccd1 _06415_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_32_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09939_ _09939_/A _09939_/B vssd1 vssd1 vccd1 vccd1 _09996_/B sky130_fd_sc_hd__nand2_1
XANTENNA__06130__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10728__RESET_B fanout98/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08338__A _08897_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10714_ _10718_/CLK _10714_/D fanout99/X vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10645_ _10539_/B _10538_/C _10538_/A vssd1 vssd1 vccd1 vccd1 _10646_/A sky130_fd_sc_hd__a21o_1
X_10576_ _10707_/B _10707_/A vssd1 vssd1 vccd1 vccd1 _10708_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_23_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10108__A _10112_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09632__A _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_05620_ _05620_/A _05620_/B _05620_/C vssd1 vssd1 vccd1 vccd1 _05623_/C sky130_fd_sc_hd__nand3_1
XANTENNA__07152__A _08114_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_05551_ _08453_/A input64/X vssd1 vssd1 vccd1 vccd1 _05600_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05482_ _08171_/B _10148_/B vssd1 vssd1 vccd1 vccd1 _05948_/A sky130_fd_sc_hd__nand2_1
X_08270_ _08297_/B _08331_/A _08269_/Y vssd1 vssd1 vccd1 vccd1 _08320_/B sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07221_ _07221_/A vssd1 vssd1 vccd1 vccd1 _07377_/B sky130_fd_sc_hd__inv_2
X_07152_ _08114_/B _10201_/A vssd1 vssd1 vccd1 vccd1 _07321_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_54_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06103_ _06921_/A _06103_/B _06103_/C vssd1 vssd1 vccd1 vccd1 _06104_/B sky130_fd_sc_hd__nand3_1
XANTENNA__05400__A _08574_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07083_ _07083_/A _07083_/B vssd1 vssd1 vccd1 vccd1 _07106_/B sky130_fd_sc_hd__nand2_1
X_06034_ _06038_/A _06841_/A vssd1 vssd1 vccd1 vccd1 _06846_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07985_ _07985_/A vssd1 vssd1 vccd1 vccd1 _07991_/A sky130_fd_sc_hd__inv_2
X_09724_ _09725_/B _09725_/A vssd1 vssd1 vccd1 vccd1 _09724_/Y sky130_fd_sc_hd__nand2_1
X_06936_ _09353_/A _06936_/B _07284_/A vssd1 vssd1 vccd1 vccd1 _06937_/B sky130_fd_sc_hd__nand3_1
X_06867_ _08842_/B _06867_/B vssd1 vssd1 vccd1 vccd1 _06870_/A sky130_fd_sc_hd__nand2_1
X_09655_ _09655_/A _09655_/B vssd1 vssd1 vccd1 vccd1 _09658_/C sky130_fd_sc_hd__nand2_1
X_08606_ _08606_/A vssd1 vssd1 vccd1 vccd1 _08611_/B sky130_fd_sc_hd__inv_2
X_05818_ input12/X vssd1 vssd1 vccd1 vccd1 _09778_/D sky130_fd_sc_hd__buf_6
X_09586_ _09586_/A _09587_/A vssd1 vssd1 vccd1 vccd1 _09589_/A sky130_fd_sc_hd__nand2_1
X_06798_ _06801_/C _06798_/B _08822_/B vssd1 vssd1 vccd1 vccd1 _08822_/A sky130_fd_sc_hd__nand3b_1
XANTENNA__08158__A _10284_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08537_ _08630_/A vssd1 vssd1 vccd1 vccd1 _08538_/B sky130_fd_sc_hd__inv_2
X_05749_ _06108_/A _06106_/A vssd1 vssd1 vccd1 vccd1 _05749_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_37_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08468_ _08869_/B vssd1 vssd1 vccd1 vccd1 _08568_/A sky130_fd_sc_hd__inv_2
XANTENNA__09680__B1 _10187_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07419_ _07835_/C _07441_/B vssd1 vssd1 vccd1 vccd1 _07439_/B sky130_fd_sc_hd__nor2b_1
X_08399_ _10157_/A _10187_/A vssd1 vssd1 vccd1 vccd1 _08403_/C sky130_fd_sc_hd__nand2_1
XANTENNA__08605__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10430_ _10430_/A _10430_/B vssd1 vssd1 vccd1 vccd1 _10435_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_33_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10361_ _10361_/A _10361_/B vssd1 vssd1 vccd1 vccd1 _10370_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_5_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10292_ input57/X _10292_/B vssd1 vssd1 vccd1 vccd1 _10293_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_135 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10628_ hold39/A hold1/X vssd1 vssd1 vccd1 vccd1 _10629_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10559_ _10559_/A vssd1 vssd1 vccd1 vccd1 _10698_/A sky130_fd_sc_hd__inv_2
XFILLER_0_59_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__05874__B input40/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ _07770_/A _07770_/B _07770_/C vssd1 vssd1 vccd1 vccd1 _07951_/A sky130_fd_sc_hd__nand3_2
X_06721_ _06721_/A _06722_/A vssd1 vssd1 vccd1 vccd1 _06724_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09440_ _09443_/B _09443_/C vssd1 vssd1 vccd1 vccd1 _09442_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_78_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06652_ _06652_/A _06652_/B _06652_/C vssd1 vssd1 vccd1 vccd1 _06660_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_59_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05603_ _05603_/A _05603_/B vssd1 vssd1 vccd1 vccd1 _05620_/A sky130_fd_sc_hd__nand2_1
X_09371_ input21/X vssd1 vssd1 vccd1 vccd1 _09373_/B sky130_fd_sc_hd__inv_2
X_06583_ _08112_/A vssd1 vssd1 vccd1 vccd1 _10275_/B sky130_fd_sc_hd__buf_8
X_05534_ _05630_/B _05631_/B _05631_/C vssd1 vssd1 vccd1 vccd1 _06016_/B sky130_fd_sc_hd__nand3_1
X_08322_ _08355_/B _08355_/A vssd1 vssd1 vccd1 vccd1 _08323_/B sky130_fd_sc_hd__nor2_1
X_08253_ _08253_/A _08253_/B vssd1 vssd1 vccd1 vccd1 _08269_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08425__B _10150_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07204_ _07204_/A _07205_/A _07205_/B vssd1 vssd1 vccd1 vccd1 _07236_/B sky130_fd_sc_hd__nand3_1
X_05465_ _08574_/A _10150_/B vssd1 vssd1 vccd1 vccd1 _05913_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_54_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08184_ _08184_/A _08184_/B vssd1 vssd1 vccd1 vccd1 _08186_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_05396_ _05396_/A _05396_/B _05396_/C vssd1 vssd1 vccd1 vccd1 _05673_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_42_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07135_ _07135_/A _07135_/B _07135_/C vssd1 vssd1 vccd1 vccd1 _07298_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_30_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07066_ _07205_/A _07066_/B vssd1 vssd1 vccd1 vccd1 _07067_/B sky130_fd_sc_hd__nand2_1
X_06017_ _06902_/B _06017_/B vssd1 vssd1 vccd1 vccd1 _06089_/B sky130_fd_sc_hd__nand2_1
XANTENNA__09256__B _09477_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08160__B _10115_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07968_ _07967_/B _07968_/B _07968_/C vssd1 vssd1 vccd1 vccd1 _07971_/B sky130_fd_sc_hd__nand3b_1
X_09707_ _09707_/A _09707_/B vssd1 vssd1 vccd1 vccd1 _09718_/A sky130_fd_sc_hd__nand2_1
X_06919_ _06919_/A _06919_/B _06919_/C vssd1 vssd1 vccd1 vccd1 _06925_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_69_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07899_ _07900_/B _07899_/B _07899_/C vssd1 vssd1 vccd1 vccd1 _08018_/B sky130_fd_sc_hd__nand3_1
XANTENNA__10211__A _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ _09637_/B _09638_/B _09963_/B vssd1 vssd1 vccd1 vccd1 _09963_/A sky130_fd_sc_hd__nand3b_1
X_09569_ _09569_/A vssd1 vssd1 vccd1 vccd1 _09570_/A sky130_fd_sc_hd__inv_2
XFILLER_0_37_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09956__A1 _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ _10413_/A _10413_/B vssd1 vssd1 vccd1 vccd1 _10681_/A sky130_fd_sc_hd__nand2_1
X_10344_ _10591_/A _10591_/C vssd1 vssd1 vccd1 vccd1 _10345_/A sky130_fd_sc_hd__nand2_1
XANTENNA__05975__A _10201_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10275_ input54/X _10275_/B vssd1 vssd1 vccd1 vccd1 _10279_/A sky130_fd_sc_hd__nand2_1
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09910__A _10156_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_68_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08245__B _08245_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08940_ _08942_/B vssd1 vssd1 vccd1 vccd1 _08941_/B sky130_fd_sc_hd__inv_2
X_08871_ _08871_/A _08871_/B vssd1 vssd1 vccd1 vccd1 _08875_/B sky130_fd_sc_hd__nand2_1
X_07822_ _07822_/A _07822_/B vssd1 vssd1 vccd1 vccd1 _07825_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09092__A input50/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _07753_/A _07753_/B _07767_/A vssd1 vssd1 vccd1 vccd1 _07951_/B sky130_fd_sc_hd__nand3_2
XANTENNA__10031__A _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06704_ _06705_/B _06705_/A vssd1 vssd1 vccd1 vccd1 _06704_/Y sky130_fd_sc_hd__nand2_1
X_07684_ _07684_/A vssd1 vssd1 vccd1 vccd1 _07687_/A sky130_fd_sc_hd__inv_2
XANTENNA__09820__A _09824_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09423_ _09424_/B _09424_/A vssd1 vssd1 vccd1 vccd1 _09615_/B sky130_fd_sc_hd__or2_1
X_06635_ _06967_/A _06968_/A vssd1 vssd1 vccd1 vccd1 _06960_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09354_ _09354_/A _09354_/B _09354_/C vssd1 vssd1 vccd1 vccd1 _09354_/Y sky130_fd_sc_hd__nand3_1
XFILLER_0_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07340__A _10040_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08305_ _08304_/B _08304_/C _08304_/A vssd1 vssd1 vccd1 vccd1 _08312_/B sky130_fd_sc_hd__o21ai_1
X_06566_ _06566_/A _06566_/B vssd1 vssd1 vccd1 vccd1 _06570_/A sky130_fd_sc_hd__nand2_1
X_09285_ _09285_/A _09285_/B _09557_/A vssd1 vssd1 vccd1 vccd1 _09292_/B sky130_fd_sc_hd__nand3_1
XFILLER_0_62_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06497_ _06497_/A _06497_/B vssd1 vssd1 vccd1 vccd1 _06696_/A sky130_fd_sc_hd__nand2_1
X_05517_ _05522_/A _05954_/A vssd1 vssd1 vccd1 vccd1 _06001_/B sky130_fd_sc_hd__nand2_1
X_08236_ _08373_/A _08372_/A vssd1 vssd1 vccd1 vccd1 _08236_/Y sky130_fd_sc_hd__nor2_1
X_05448_ _05454_/B vssd1 vssd1 vccd1 vccd1 _05449_/B sky130_fd_sc_hd__inv_2
XFILLER_0_15_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08167_ _08167_/A _08167_/B vssd1 vssd1 vccd1 vccd1 _08169_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09267__A _10211_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07118_ _07118_/A _07118_/B _07118_/C vssd1 vssd1 vccd1 vccd1 _07427_/C sky130_fd_sc_hd__nand3_1
X_05379_ _05384_/A _05384_/C vssd1 vssd1 vccd1 vccd1 _05382_/A sky130_fd_sc_hd__nand2_1
X_08098_ _08100_/B vssd1 vssd1 vccd1 vccd1 _08099_/B sky130_fd_sc_hd__inv_2
XANTENNA__08171__A _09778_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07049_ _09517_/C vssd1 vssd1 vccd1 vccd1 _09840_/B sky130_fd_sc_hd__buf_8
X_10060_ _10060_/A vssd1 vssd1 vccd1 vccd1 _10061_/B sky130_fd_sc_hd__inv_2
XFILLER_0_65_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10327_ _10329_/B vssd1 vssd1 vccd1 vccd1 _10328_/B sky130_fd_sc_hd__inv_2
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10258_ _10263_/A _10263_/C vssd1 vssd1 vccd1 vccd1 _10262_/A sky130_fd_sc_hd__nand2_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10189_ _09602_/B _10005_/A _09678_/C _09922_/B vssd1 vssd1 vccd1 vccd1 _10190_/B
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06420_ _06431_/A vssd1 vssd1 vccd1 vccd1 _06430_/B sky130_fd_sc_hd__inv_2
XFILLER_0_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06351_ _08739_/A input35/X vssd1 vssd1 vccd1 vccd1 _06547_/C sky130_fd_sc_hd__nand2_1
XFILLER_0_29_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09070_ _09072_/B _09072_/C vssd1 vssd1 vccd1 vccd1 _09071_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06282_ _06282_/A _06282_/B _06282_/C vssd1 vssd1 vccd1 vccd1 _06285_/A sky130_fd_sc_hd__nand3_1
XFILLER_0_71_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08021_ _09551_/C _09971_/A _08021_/C vssd1 vssd1 vccd1 vccd1 _08032_/B sky130_fd_sc_hd__nor3_1
XFILLER_0_12_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09972_ _09972_/A vssd1 vssd1 vccd1 vccd1 _10127_/B sky130_fd_sc_hd__inv_2
X_08923_ _08925_/B vssd1 vssd1 vccd1 vccd1 _08928_/A sky130_fd_sc_hd__inv_2
XFILLER_0_12_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08854_ _08854_/A vssd1 vssd1 vccd1 vccd1 _08855_/B sky130_fd_sc_hd__inv_2
X_08785_ _10247_/B _09698_/A vssd1 vssd1 vccd1 vccd1 _08786_/C sky130_fd_sc_hd__nand2_1
X_05997_ _05997_/A _05997_/B vssd1 vssd1 vccd1 vccd1 _06005_/B sky130_fd_sc_hd__nand2_1
X_07805_ _07943_/B _07942_/A _07943_/C vssd1 vssd1 vccd1 vccd1 _07867_/A sky130_fd_sc_hd__a21boi_4
XANTENNA__07335__A _10103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07736_ _07736_/A _07736_/B _07736_/C vssd1 vssd1 vccd1 vccd1 _07737_/B sky130_fd_sc_hd__nand3_1
X_07667_ _07667_/A _07667_/B _07667_/C vssd1 vssd1 vccd1 vccd1 _07668_/B sky130_fd_sc_hd__nand3_1
X_09406_ _09406_/A vssd1 vssd1 vccd1 vccd1 _09407_/C sky130_fd_sc_hd__inv_2
X_07598_ _07598_/A _07598_/B vssd1 vssd1 vccd1 vccd1 _10452_/A sky130_fd_sc_hd__nand2_1
X_06618_ _06957_/B _06957_/C vssd1 vssd1 vccd1 vccd1 _06962_/A sky130_fd_sc_hd__nand2_1
X_09337_ _09354_/B _09354_/C vssd1 vssd1 vccd1 vccd1 _09338_/B sky130_fd_sc_hd__nand2_1
X_06549_ _06549_/A _06549_/B _06549_/C vssd1 vssd1 vccd1 vccd1 _06553_/C sky130_fd_sc_hd__nand3_1
X_09268_ _09268_/A _10248_/D _09268_/C vssd1 vssd1 vccd1 vccd1 _09270_/A sky130_fd_sc_hd__nor3_1
XFILLER_0_62_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08219_ _08219_/A _08219_/B vssd1 vssd1 vccd1 vccd1 _08222_/B sky130_fd_sc_hd__nand2_1
X_09199_ _10004_/A _10148_/A vssd1 vssd1 vccd1 vccd1 _09205_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09387__A2 _10158_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10112_ _10112_/A input21/X vssd1 vssd1 vccd1 vccd1 _10113_/B sky130_fd_sc_hd__nand2_1
Xhold40 hold40/A vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
X_10043_ input46/X _10211_/B _10211_/A _10210_/B vssd1 vssd1 vccd1 vccd1 _10043_/X
+ sky130_fd_sc_hd__a22o_1
Xhold51 hold51/A vssd1 vssd1 vccd1 vccd1 hold51/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 hold62/A vssd1 vssd1 vccd1 vccd1 hold62/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_05920_ input15/X vssd1 vssd1 vccd1 vccd1 _10158_/B sky130_fd_sc_hd__buf_4
X_05851_ _06302_/B _05851_/B vssd1 vssd1 vccd1 vccd1 _06118_/C sky130_fd_sc_hd__nand2_1
X_08570_ _08570_/A _08570_/B vssd1 vssd1 vccd1 vccd1 _08624_/A sky130_fd_sc_hd__nand2_1
X_05782_ _05786_/A vssd1 vssd1 vccd1 vccd1 _05785_/A sky130_fd_sc_hd__inv_2
XANTENNA__09370__A _10101_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07521_ _07667_/B _07667_/C vssd1 vssd1 vccd1 vccd1 _07666_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_76_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_72 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07452_ _07452_/A _07452_/B vssd1 vssd1 vccd1 vccd1 _07453_/A sky130_fd_sc_hd__nand2_1
X_07383_ _07383_/A vssd1 vssd1 vccd1 vccd1 _07482_/B sky130_fd_sc_hd__inv_2
XFILLER_0_8_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06403_ _06566_/A _06567_/A vssd1 vssd1 vccd1 vccd1 _06403_/Y sky130_fd_sc_hd__nand2_1
X_09122_ _09122_/A _09122_/B vssd1 vssd1 vccd1 vccd1 _09126_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_44_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06334_ _08672_/A _07785_/B vssd1 vssd1 vccd1 vccd1 _06506_/B sky130_fd_sc_hd__nand2_1
X_09053_ _09053_/A _09053_/B _09053_/C vssd1 vssd1 vccd1 vccd1 _09077_/C sky130_fd_sc_hd__nand3_1
XFILLER_0_25_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06265_ _06267_/A _06265_/B vssd1 vssd1 vccd1 vccd1 _06266_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08004_ _10247_/B _08114_/B vssd1 vssd1 vccd1 vccd1 _08119_/B sky130_fd_sc_hd__nand2_1
X_06196_ _06196_/A _06196_/B vssd1 vssd1 vccd1 vccd1 _06196_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_40_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09955_ _09955_/A vssd1 vssd1 vccd1 vccd1 _09957_/A sky130_fd_sc_hd__inv_2
X_08906_ _08797_/A _08905_/Y _08798_/A vssd1 vssd1 vccd1 vccd1 _08907_/B sky130_fd_sc_hd__a21oi_1
X_09886_ _10274_/B _10274_/A vssd1 vssd1 vccd1 vccd1 _09889_/C sky130_fd_sc_hd__nand2_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08837_ _08840_/A _08840_/B vssd1 vssd1 vccd1 vccd1 _08839_/A sky130_fd_sc_hd__nand2_1
X_08768_ _08833_/B _08833_/C vssd1 vssd1 vccd1 vccd1 _08832_/A sky130_fd_sc_hd__nand2_1
X_08699_ _09228_/C _08699_/B vssd1 vssd1 vccd1 vccd1 _08701_/A sky130_fd_sc_hd__xor2_1
X_07719_ _07719_/A _07828_/B _07828_/A vssd1 vssd1 vccd1 vccd1 _08075_/A sky130_fd_sc_hd__nand3_4
X_10730_ _10741_/CLK _10730_/D fanout98/X vssd1 vssd1 vccd1 vccd1 hold64/A sky130_fd_sc_hd__dfrtp_2
XANTENNA__08608__B _10156_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10661_ _10661_/A hold34/X vssd1 vssd1 vccd1 vccd1 hold35/A sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06128__B _10148_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10592_ _10594_/A _10592_/B vssd1 vssd1 vccd1 vccd1 _10596_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_35_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09780__A2 _10275_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput85 hold12/A vssd1 vssd1 vccd1 vccd1 y_o[27] sky130_fd_sc_hd__buf_12
Xoutput74 hold31/A vssd1 vssd1 vccd1 vccd1 y_o[17] sky130_fd_sc_hd__buf_12
Xoutput96 hold43/A vssd1 vssd1 vccd1 vccd1 y_o[8] sky130_fd_sc_hd__buf_12
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10026_ _10052_/B _10052_/C vssd1 vssd1 vccd1 vccd1 _10051_/A sky130_fd_sc_hd__nand2_1
XANTENNA__09190__A _10157_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06050_ _09477_/C vssd1 vssd1 vccd1 vccd1 _10202_/C sky130_fd_sc_hd__inv_2
XFILLER_0_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06989__A _10212_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ _09742_/A vssd1 vssd1 vccd1 vccd1 _09741_/B sky130_fd_sc_hd__inv_2
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06952_ _06952_/A _06952_/B _06952_/C vssd1 vssd1 vccd1 vccd1 _07113_/B sky130_fd_sc_hd__nand3_1
.ends

