magic
tech sky130A
magscale 1 2
timestamp 1759765050
<< obsli1 >>
rect 1104 2159 198812 197489
<< obsm1 >>
rect 934 1232 198982 197520
<< metal2 >>
rect 4894 199200 4950 200000
rect 6090 199200 6146 200000
rect 7286 199200 7342 200000
rect 8482 199200 8538 200000
rect 9678 199200 9734 200000
rect 10874 199200 10930 200000
rect 12070 199200 12126 200000
rect 13266 199200 13322 200000
rect 14462 199200 14518 200000
rect 15658 199200 15714 200000
rect 16854 199200 16910 200000
rect 18050 199200 18106 200000
rect 19246 199200 19302 200000
rect 20442 199200 20498 200000
rect 21638 199200 21694 200000
rect 22834 199200 22890 200000
rect 24030 199200 24086 200000
rect 25226 199200 25282 200000
rect 26422 199200 26478 200000
rect 27618 199200 27674 200000
rect 28814 199200 28870 200000
rect 30010 199200 30066 200000
rect 31206 199200 31262 200000
rect 32402 199200 32458 200000
rect 33598 199200 33654 200000
rect 34794 199200 34850 200000
rect 35990 199200 36046 200000
rect 37186 199200 37242 200000
rect 38382 199200 38438 200000
rect 39578 199200 39634 200000
rect 40774 199200 40830 200000
rect 41970 199200 42026 200000
rect 43166 199200 43222 200000
rect 44362 199200 44418 200000
rect 45558 199200 45614 200000
rect 46754 199200 46810 200000
rect 47950 199200 48006 200000
rect 49146 199200 49202 200000
rect 50342 199200 50398 200000
rect 51538 199200 51594 200000
rect 52734 199200 52790 200000
rect 53930 199200 53986 200000
rect 55126 199200 55182 200000
rect 56322 199200 56378 200000
rect 57518 199200 57574 200000
rect 58714 199200 58770 200000
rect 59910 199200 59966 200000
rect 61106 199200 61162 200000
rect 62302 199200 62358 200000
rect 63498 199200 63554 200000
rect 64694 199200 64750 200000
rect 65890 199200 65946 200000
rect 67086 199200 67142 200000
rect 68282 199200 68338 200000
rect 69478 199200 69534 200000
rect 70674 199200 70730 200000
rect 71870 199200 71926 200000
rect 73066 199200 73122 200000
rect 74262 199200 74318 200000
rect 75458 199200 75514 200000
rect 76654 199200 76710 200000
rect 77850 199200 77906 200000
rect 79046 199200 79102 200000
rect 80242 199200 80298 200000
rect 81438 199200 81494 200000
rect 82634 199200 82690 200000
rect 83830 199200 83886 200000
rect 85026 199200 85082 200000
rect 86222 199200 86278 200000
rect 87418 199200 87474 200000
rect 88614 199200 88670 200000
rect 89810 199200 89866 200000
rect 91006 199200 91062 200000
rect 92202 199200 92258 200000
rect 93398 199200 93454 200000
rect 94594 199200 94650 200000
rect 95790 199200 95846 200000
rect 96986 199200 97042 200000
rect 98182 199200 98238 200000
rect 99378 199200 99434 200000
rect 100574 199200 100630 200000
rect 101770 199200 101826 200000
rect 102966 199200 103022 200000
rect 104162 199200 104218 200000
rect 105358 199200 105414 200000
rect 106554 199200 106610 200000
rect 107750 199200 107806 200000
rect 108946 199200 109002 200000
rect 110142 199200 110198 200000
rect 111338 199200 111394 200000
rect 112534 199200 112590 200000
rect 113730 199200 113786 200000
rect 114926 199200 114982 200000
rect 116122 199200 116178 200000
rect 117318 199200 117374 200000
rect 118514 199200 118570 200000
rect 119710 199200 119766 200000
rect 120906 199200 120962 200000
rect 122102 199200 122158 200000
rect 123298 199200 123354 200000
rect 124494 199200 124550 200000
rect 125690 199200 125746 200000
rect 126886 199200 126942 200000
rect 128082 199200 128138 200000
rect 129278 199200 129334 200000
rect 130474 199200 130530 200000
rect 131670 199200 131726 200000
rect 132866 199200 132922 200000
rect 134062 199200 134118 200000
rect 135258 199200 135314 200000
rect 136454 199200 136510 200000
rect 137650 199200 137706 200000
rect 138846 199200 138902 200000
rect 140042 199200 140098 200000
rect 141238 199200 141294 200000
rect 142434 199200 142490 200000
rect 143630 199200 143686 200000
rect 144826 199200 144882 200000
rect 146022 199200 146078 200000
rect 147218 199200 147274 200000
rect 148414 199200 148470 200000
rect 149610 199200 149666 200000
rect 150806 199200 150862 200000
rect 152002 199200 152058 200000
rect 153198 199200 153254 200000
rect 154394 199200 154450 200000
rect 155590 199200 155646 200000
rect 156786 199200 156842 200000
rect 157982 199200 158038 200000
rect 159178 199200 159234 200000
rect 160374 199200 160430 200000
rect 161570 199200 161626 200000
rect 162766 199200 162822 200000
rect 163962 199200 164018 200000
rect 165158 199200 165214 200000
rect 166354 199200 166410 200000
rect 167550 199200 167606 200000
rect 168746 199200 168802 200000
rect 169942 199200 169998 200000
rect 171138 199200 171194 200000
rect 172334 199200 172390 200000
rect 173530 199200 173586 200000
rect 174726 199200 174782 200000
rect 175922 199200 175978 200000
rect 177118 199200 177174 200000
rect 178314 199200 178370 200000
rect 179510 199200 179566 200000
rect 180706 199200 180762 200000
rect 181902 199200 181958 200000
rect 183098 199200 183154 200000
rect 184294 199200 184350 200000
rect 185490 199200 185546 200000
rect 186686 199200 186742 200000
rect 187882 199200 187938 200000
rect 189078 199200 189134 200000
rect 190274 199200 190330 200000
rect 191470 199200 191526 200000
rect 192666 199200 192722 200000
rect 193862 199200 193918 200000
rect 195058 199200 195114 200000
rect 4894 0 4950 800
rect 6090 0 6146 800
rect 7286 0 7342 800
rect 8482 0 8538 800
rect 9678 0 9734 800
rect 10874 0 10930 800
rect 12070 0 12126 800
rect 13266 0 13322 800
rect 14462 0 14518 800
rect 15658 0 15714 800
rect 16854 0 16910 800
rect 18050 0 18106 800
rect 19246 0 19302 800
rect 20442 0 20498 800
rect 21638 0 21694 800
rect 22834 0 22890 800
rect 24030 0 24086 800
rect 25226 0 25282 800
rect 26422 0 26478 800
rect 27618 0 27674 800
rect 28814 0 28870 800
rect 30010 0 30066 800
rect 31206 0 31262 800
rect 32402 0 32458 800
rect 33598 0 33654 800
rect 34794 0 34850 800
rect 35990 0 36046 800
rect 37186 0 37242 800
rect 38382 0 38438 800
rect 39578 0 39634 800
rect 40774 0 40830 800
rect 41970 0 42026 800
rect 43166 0 43222 800
rect 44362 0 44418 800
rect 45558 0 45614 800
rect 46754 0 46810 800
rect 47950 0 48006 800
rect 49146 0 49202 800
rect 50342 0 50398 800
rect 51538 0 51594 800
rect 52734 0 52790 800
rect 53930 0 53986 800
rect 55126 0 55182 800
rect 56322 0 56378 800
rect 57518 0 57574 800
rect 58714 0 58770 800
rect 59910 0 59966 800
rect 61106 0 61162 800
rect 62302 0 62358 800
rect 63498 0 63554 800
rect 64694 0 64750 800
rect 65890 0 65946 800
rect 67086 0 67142 800
rect 68282 0 68338 800
rect 69478 0 69534 800
rect 70674 0 70730 800
rect 71870 0 71926 800
rect 73066 0 73122 800
rect 74262 0 74318 800
rect 75458 0 75514 800
rect 76654 0 76710 800
rect 77850 0 77906 800
rect 79046 0 79102 800
rect 80242 0 80298 800
rect 81438 0 81494 800
rect 82634 0 82690 800
rect 83830 0 83886 800
rect 85026 0 85082 800
rect 86222 0 86278 800
rect 87418 0 87474 800
rect 88614 0 88670 800
rect 89810 0 89866 800
rect 91006 0 91062 800
rect 92202 0 92258 800
rect 93398 0 93454 800
rect 94594 0 94650 800
rect 95790 0 95846 800
rect 96986 0 97042 800
rect 98182 0 98238 800
rect 99378 0 99434 800
rect 100574 0 100630 800
rect 101770 0 101826 800
rect 102966 0 103022 800
rect 104162 0 104218 800
rect 105358 0 105414 800
rect 106554 0 106610 800
rect 107750 0 107806 800
rect 108946 0 109002 800
rect 110142 0 110198 800
rect 111338 0 111394 800
rect 112534 0 112590 800
rect 113730 0 113786 800
rect 114926 0 114982 800
rect 116122 0 116178 800
rect 117318 0 117374 800
rect 118514 0 118570 800
rect 119710 0 119766 800
rect 120906 0 120962 800
rect 122102 0 122158 800
rect 123298 0 123354 800
rect 124494 0 124550 800
rect 125690 0 125746 800
rect 126886 0 126942 800
rect 128082 0 128138 800
rect 129278 0 129334 800
rect 130474 0 130530 800
rect 131670 0 131726 800
rect 132866 0 132922 800
rect 134062 0 134118 800
rect 135258 0 135314 800
rect 136454 0 136510 800
rect 137650 0 137706 800
rect 138846 0 138902 800
rect 140042 0 140098 800
rect 141238 0 141294 800
rect 142434 0 142490 800
rect 143630 0 143686 800
rect 144826 0 144882 800
rect 146022 0 146078 800
rect 147218 0 147274 800
rect 148414 0 148470 800
rect 149610 0 149666 800
rect 150806 0 150862 800
rect 152002 0 152058 800
rect 153198 0 153254 800
rect 154394 0 154450 800
rect 155590 0 155646 800
rect 156786 0 156842 800
rect 157982 0 158038 800
rect 159178 0 159234 800
rect 160374 0 160430 800
rect 161570 0 161626 800
rect 162766 0 162822 800
rect 163962 0 164018 800
rect 165158 0 165214 800
rect 166354 0 166410 800
rect 167550 0 167606 800
rect 168746 0 168802 800
rect 169942 0 169998 800
rect 171138 0 171194 800
rect 172334 0 172390 800
rect 173530 0 173586 800
rect 174726 0 174782 800
rect 175922 0 175978 800
rect 177118 0 177174 800
rect 178314 0 178370 800
rect 179510 0 179566 800
rect 180706 0 180762 800
rect 181902 0 181958 800
rect 183098 0 183154 800
rect 184294 0 184350 800
rect 185490 0 185546 800
rect 186686 0 186742 800
rect 187882 0 187938 800
rect 189078 0 189134 800
rect 190274 0 190330 800
rect 191470 0 191526 800
rect 192666 0 192722 800
rect 193862 0 193918 800
rect 195058 0 195114 800
<< obsm2 >>
rect 938 199144 4838 199322
rect 5006 199144 6034 199322
rect 6202 199144 7230 199322
rect 7398 199144 8426 199322
rect 8594 199144 9622 199322
rect 9790 199144 10818 199322
rect 10986 199144 12014 199322
rect 12182 199144 13210 199322
rect 13378 199144 14406 199322
rect 14574 199144 15602 199322
rect 15770 199144 16798 199322
rect 16966 199144 17994 199322
rect 18162 199144 19190 199322
rect 19358 199144 20386 199322
rect 20554 199144 21582 199322
rect 21750 199144 22778 199322
rect 22946 199144 23974 199322
rect 24142 199144 25170 199322
rect 25338 199144 26366 199322
rect 26534 199144 27562 199322
rect 27730 199144 28758 199322
rect 28926 199144 29954 199322
rect 30122 199144 31150 199322
rect 31318 199144 32346 199322
rect 32514 199144 33542 199322
rect 33710 199144 34738 199322
rect 34906 199144 35934 199322
rect 36102 199144 37130 199322
rect 37298 199144 38326 199322
rect 38494 199144 39522 199322
rect 39690 199144 40718 199322
rect 40886 199144 41914 199322
rect 42082 199144 43110 199322
rect 43278 199144 44306 199322
rect 44474 199144 45502 199322
rect 45670 199144 46698 199322
rect 46866 199144 47894 199322
rect 48062 199144 49090 199322
rect 49258 199144 50286 199322
rect 50454 199144 51482 199322
rect 51650 199144 52678 199322
rect 52846 199144 53874 199322
rect 54042 199144 55070 199322
rect 55238 199144 56266 199322
rect 56434 199144 57462 199322
rect 57630 199144 58658 199322
rect 58826 199144 59854 199322
rect 60022 199144 61050 199322
rect 61218 199144 62246 199322
rect 62414 199144 63442 199322
rect 63610 199144 64638 199322
rect 64806 199144 65834 199322
rect 66002 199144 67030 199322
rect 67198 199144 68226 199322
rect 68394 199144 69422 199322
rect 69590 199144 70618 199322
rect 70786 199144 71814 199322
rect 71982 199144 73010 199322
rect 73178 199144 74206 199322
rect 74374 199144 75402 199322
rect 75570 199144 76598 199322
rect 76766 199144 77794 199322
rect 77962 199144 78990 199322
rect 79158 199144 80186 199322
rect 80354 199144 81382 199322
rect 81550 199144 82578 199322
rect 82746 199144 83774 199322
rect 83942 199144 84970 199322
rect 85138 199144 86166 199322
rect 86334 199144 87362 199322
rect 87530 199144 88558 199322
rect 88726 199144 89754 199322
rect 89922 199144 90950 199322
rect 91118 199144 92146 199322
rect 92314 199144 93342 199322
rect 93510 199144 94538 199322
rect 94706 199144 95734 199322
rect 95902 199144 96930 199322
rect 97098 199144 98126 199322
rect 98294 199144 99322 199322
rect 99490 199144 100518 199322
rect 100686 199144 101714 199322
rect 101882 199144 102910 199322
rect 103078 199144 104106 199322
rect 104274 199144 105302 199322
rect 105470 199144 106498 199322
rect 106666 199144 107694 199322
rect 107862 199144 108890 199322
rect 109058 199144 110086 199322
rect 110254 199144 111282 199322
rect 111450 199144 112478 199322
rect 112646 199144 113674 199322
rect 113842 199144 114870 199322
rect 115038 199144 116066 199322
rect 116234 199144 117262 199322
rect 117430 199144 118458 199322
rect 118626 199144 119654 199322
rect 119822 199144 120850 199322
rect 121018 199144 122046 199322
rect 122214 199144 123242 199322
rect 123410 199144 124438 199322
rect 124606 199144 125634 199322
rect 125802 199144 126830 199322
rect 126998 199144 128026 199322
rect 128194 199144 129222 199322
rect 129390 199144 130418 199322
rect 130586 199144 131614 199322
rect 131782 199144 132810 199322
rect 132978 199144 134006 199322
rect 134174 199144 135202 199322
rect 135370 199144 136398 199322
rect 136566 199144 137594 199322
rect 137762 199144 138790 199322
rect 138958 199144 139986 199322
rect 140154 199144 141182 199322
rect 141350 199144 142378 199322
rect 142546 199144 143574 199322
rect 143742 199144 144770 199322
rect 144938 199144 145966 199322
rect 146134 199144 147162 199322
rect 147330 199144 148358 199322
rect 148526 199144 149554 199322
rect 149722 199144 150750 199322
rect 150918 199144 151946 199322
rect 152114 199144 153142 199322
rect 153310 199144 154338 199322
rect 154506 199144 155534 199322
rect 155702 199144 156730 199322
rect 156898 199144 157926 199322
rect 158094 199144 159122 199322
rect 159290 199144 160318 199322
rect 160486 199144 161514 199322
rect 161682 199144 162710 199322
rect 162878 199144 163906 199322
rect 164074 199144 165102 199322
rect 165270 199144 166298 199322
rect 166466 199144 167494 199322
rect 167662 199144 168690 199322
rect 168858 199144 169886 199322
rect 170054 199144 171082 199322
rect 171250 199144 172278 199322
rect 172446 199144 173474 199322
rect 173642 199144 174670 199322
rect 174838 199144 175866 199322
rect 176034 199144 177062 199322
rect 177230 199144 178258 199322
rect 178426 199144 179454 199322
rect 179622 199144 180650 199322
rect 180818 199144 181846 199322
rect 182014 199144 183042 199322
rect 183210 199144 184238 199322
rect 184406 199144 185434 199322
rect 185602 199144 186630 199322
rect 186798 199144 187826 199322
rect 187994 199144 189022 199322
rect 189190 199144 190218 199322
rect 190386 199144 191414 199322
rect 191582 199144 192610 199322
rect 192778 199144 193806 199322
rect 193974 199144 195002 199322
rect 195170 199144 198978 199322
rect 938 856 198978 199144
rect 938 734 4838 856
rect 5006 734 6034 856
rect 6202 734 7230 856
rect 7398 734 8426 856
rect 8594 734 9622 856
rect 9790 734 10818 856
rect 10986 734 12014 856
rect 12182 734 13210 856
rect 13378 734 14406 856
rect 14574 734 15602 856
rect 15770 734 16798 856
rect 16966 734 17994 856
rect 18162 734 19190 856
rect 19358 734 20386 856
rect 20554 734 21582 856
rect 21750 734 22778 856
rect 22946 734 23974 856
rect 24142 734 25170 856
rect 25338 734 26366 856
rect 26534 734 27562 856
rect 27730 734 28758 856
rect 28926 734 29954 856
rect 30122 734 31150 856
rect 31318 734 32346 856
rect 32514 734 33542 856
rect 33710 734 34738 856
rect 34906 734 35934 856
rect 36102 734 37130 856
rect 37298 734 38326 856
rect 38494 734 39522 856
rect 39690 734 40718 856
rect 40886 734 41914 856
rect 42082 734 43110 856
rect 43278 734 44306 856
rect 44474 734 45502 856
rect 45670 734 46698 856
rect 46866 734 47894 856
rect 48062 734 49090 856
rect 49258 734 50286 856
rect 50454 734 51482 856
rect 51650 734 52678 856
rect 52846 734 53874 856
rect 54042 734 55070 856
rect 55238 734 56266 856
rect 56434 734 57462 856
rect 57630 734 58658 856
rect 58826 734 59854 856
rect 60022 734 61050 856
rect 61218 734 62246 856
rect 62414 734 63442 856
rect 63610 734 64638 856
rect 64806 734 65834 856
rect 66002 734 67030 856
rect 67198 734 68226 856
rect 68394 734 69422 856
rect 69590 734 70618 856
rect 70786 734 71814 856
rect 71982 734 73010 856
rect 73178 734 74206 856
rect 74374 734 75402 856
rect 75570 734 76598 856
rect 76766 734 77794 856
rect 77962 734 78990 856
rect 79158 734 80186 856
rect 80354 734 81382 856
rect 81550 734 82578 856
rect 82746 734 83774 856
rect 83942 734 84970 856
rect 85138 734 86166 856
rect 86334 734 87362 856
rect 87530 734 88558 856
rect 88726 734 89754 856
rect 89922 734 90950 856
rect 91118 734 92146 856
rect 92314 734 93342 856
rect 93510 734 94538 856
rect 94706 734 95734 856
rect 95902 734 96930 856
rect 97098 734 98126 856
rect 98294 734 99322 856
rect 99490 734 100518 856
rect 100686 734 101714 856
rect 101882 734 102910 856
rect 103078 734 104106 856
rect 104274 734 105302 856
rect 105470 734 106498 856
rect 106666 734 107694 856
rect 107862 734 108890 856
rect 109058 734 110086 856
rect 110254 734 111282 856
rect 111450 734 112478 856
rect 112646 734 113674 856
rect 113842 734 114870 856
rect 115038 734 116066 856
rect 116234 734 117262 856
rect 117430 734 118458 856
rect 118626 734 119654 856
rect 119822 734 120850 856
rect 121018 734 122046 856
rect 122214 734 123242 856
rect 123410 734 124438 856
rect 124606 734 125634 856
rect 125802 734 126830 856
rect 126998 734 128026 856
rect 128194 734 129222 856
rect 129390 734 130418 856
rect 130586 734 131614 856
rect 131782 734 132810 856
rect 132978 734 134006 856
rect 134174 734 135202 856
rect 135370 734 136398 856
rect 136566 734 137594 856
rect 137762 734 138790 856
rect 138958 734 139986 856
rect 140154 734 141182 856
rect 141350 734 142378 856
rect 142546 734 143574 856
rect 143742 734 144770 856
rect 144938 734 145966 856
rect 146134 734 147162 856
rect 147330 734 148358 856
rect 148526 734 149554 856
rect 149722 734 150750 856
rect 150918 734 151946 856
rect 152114 734 153142 856
rect 153310 734 154338 856
rect 154506 734 155534 856
rect 155702 734 156730 856
rect 156898 734 157926 856
rect 158094 734 159122 856
rect 159290 734 160318 856
rect 160486 734 161514 856
rect 161682 734 162710 856
rect 162878 734 163906 856
rect 164074 734 165102 856
rect 165270 734 166298 856
rect 166466 734 167494 856
rect 167662 734 168690 856
rect 168858 734 169886 856
rect 170054 734 171082 856
rect 171250 734 172278 856
rect 172446 734 173474 856
rect 173642 734 174670 856
rect 174838 734 175866 856
rect 176034 734 177062 856
rect 177230 734 178258 856
rect 178426 734 179454 856
rect 179622 734 180650 856
rect 180818 734 181846 856
rect 182014 734 183042 856
rect 183210 734 184238 856
rect 184406 734 185434 856
rect 185602 734 186630 856
rect 186798 734 187826 856
rect 187994 734 189022 856
rect 189190 734 190218 856
rect 190386 734 191414 856
rect 191582 734 192610 856
rect 192778 734 193806 856
rect 193974 734 195002 856
rect 195170 734 198978 856
<< metal3 >>
rect 0 190136 800 190256
rect 0 188232 800 188352
rect 0 186328 800 186448
rect 199200 186328 200000 186448
rect 199200 185240 200000 185360
rect 0 184424 800 184544
rect 199200 184152 200000 184272
rect 199200 183064 200000 183184
rect 0 182520 800 182640
rect 199200 181976 200000 182096
rect 199200 180888 200000 181008
rect 0 180616 800 180736
rect 199200 179800 200000 179920
rect 0 178712 800 178832
rect 199200 178712 200000 178832
rect 199200 177624 200000 177744
rect 0 176808 800 176928
rect 199200 176536 200000 176656
rect 199200 175448 200000 175568
rect 0 174904 800 175024
rect 199200 174360 200000 174480
rect 199200 173272 200000 173392
rect 0 173000 800 173120
rect 199200 172184 200000 172304
rect 0 171096 800 171216
rect 199200 171096 200000 171216
rect 199200 170008 200000 170128
rect 0 169192 800 169312
rect 199200 168920 200000 169040
rect 199200 167832 200000 167952
rect 0 167288 800 167408
rect 199200 166744 200000 166864
rect 199200 165656 200000 165776
rect 0 165384 800 165504
rect 199200 164568 200000 164688
rect 0 163480 800 163600
rect 199200 163480 200000 163600
rect 199200 162392 200000 162512
rect 0 161576 800 161696
rect 199200 161304 200000 161424
rect 199200 160216 200000 160336
rect 0 159672 800 159792
rect 199200 159128 200000 159248
rect 199200 158040 200000 158160
rect 0 157768 800 157888
rect 199200 156952 200000 157072
rect 0 155864 800 155984
rect 199200 155864 200000 155984
rect 199200 154776 200000 154896
rect 0 153960 800 154080
rect 199200 153688 200000 153808
rect 199200 152600 200000 152720
rect 0 152056 800 152176
rect 199200 151512 200000 151632
rect 199200 150424 200000 150544
rect 0 150152 800 150272
rect 199200 149336 200000 149456
rect 0 148248 800 148368
rect 199200 148248 200000 148368
rect 199200 147160 200000 147280
rect 0 146344 800 146464
rect 199200 146072 200000 146192
rect 199200 144984 200000 145104
rect 0 144440 800 144560
rect 199200 143896 200000 144016
rect 199200 142808 200000 142928
rect 0 142536 800 142656
rect 199200 141720 200000 141840
rect 0 140632 800 140752
rect 199200 140632 200000 140752
rect 199200 139544 200000 139664
rect 0 138728 800 138848
rect 199200 138456 200000 138576
rect 199200 137368 200000 137488
rect 0 136824 800 136944
rect 199200 136280 200000 136400
rect 199200 135192 200000 135312
rect 0 134920 800 135040
rect 199200 134104 200000 134224
rect 0 133016 800 133136
rect 199200 133016 200000 133136
rect 199200 131928 200000 132048
rect 0 131112 800 131232
rect 199200 130840 200000 130960
rect 199200 129752 200000 129872
rect 0 129208 800 129328
rect 199200 128664 200000 128784
rect 199200 127576 200000 127696
rect 0 127304 800 127424
rect 199200 126488 200000 126608
rect 0 125400 800 125520
rect 199200 125400 200000 125520
rect 199200 124312 200000 124432
rect 0 123496 800 123616
rect 199200 123224 200000 123344
rect 199200 122136 200000 122256
rect 0 121592 800 121712
rect 199200 121048 200000 121168
rect 199200 119960 200000 120080
rect 0 119688 800 119808
rect 199200 118872 200000 118992
rect 0 117784 800 117904
rect 199200 117784 200000 117904
rect 199200 116696 200000 116816
rect 0 115880 800 116000
rect 199200 115608 200000 115728
rect 199200 114520 200000 114640
rect 0 113976 800 114096
rect 199200 113432 200000 113552
rect 199200 112344 200000 112464
rect 0 112072 800 112192
rect 199200 111256 200000 111376
rect 0 110168 800 110288
rect 199200 110168 200000 110288
rect 199200 109080 200000 109200
rect 0 108264 800 108384
rect 199200 107992 200000 108112
rect 199200 106904 200000 107024
rect 0 106360 800 106480
rect 199200 105816 200000 105936
rect 199200 104728 200000 104848
rect 0 104456 800 104576
rect 199200 103640 200000 103760
rect 0 102552 800 102672
rect 199200 102552 200000 102672
rect 199200 101464 200000 101584
rect 0 100648 800 100768
rect 199200 100376 200000 100496
rect 199200 99288 200000 99408
rect 0 98744 800 98864
rect 199200 98200 200000 98320
rect 199200 97112 200000 97232
rect 0 96840 800 96960
rect 199200 96024 200000 96144
rect 0 94936 800 95056
rect 199200 94936 200000 95056
rect 199200 93848 200000 93968
rect 0 93032 800 93152
rect 199200 92760 200000 92880
rect 199200 91672 200000 91792
rect 0 91128 800 91248
rect 199200 90584 200000 90704
rect 199200 89496 200000 89616
rect 0 89224 800 89344
rect 199200 88408 200000 88528
rect 0 87320 800 87440
rect 199200 87320 200000 87440
rect 199200 86232 200000 86352
rect 0 85416 800 85536
rect 199200 85144 200000 85264
rect 199200 84056 200000 84176
rect 0 83512 800 83632
rect 199200 82968 200000 83088
rect 199200 81880 200000 82000
rect 0 81608 800 81728
rect 199200 80792 200000 80912
rect 0 79704 800 79824
rect 199200 79704 200000 79824
rect 199200 78616 200000 78736
rect 0 77800 800 77920
rect 199200 77528 200000 77648
rect 199200 76440 200000 76560
rect 0 75896 800 76016
rect 199200 75352 200000 75472
rect 199200 74264 200000 74384
rect 0 73992 800 74112
rect 199200 73176 200000 73296
rect 0 72088 800 72208
rect 199200 72088 200000 72208
rect 199200 71000 200000 71120
rect 0 70184 800 70304
rect 199200 69912 200000 70032
rect 199200 68824 200000 68944
rect 0 68280 800 68400
rect 199200 67736 200000 67856
rect 199200 66648 200000 66768
rect 0 66376 800 66496
rect 199200 65560 200000 65680
rect 0 64472 800 64592
rect 199200 64472 200000 64592
rect 199200 63384 200000 63504
rect 0 62568 800 62688
rect 199200 62296 200000 62416
rect 199200 61208 200000 61328
rect 0 60664 800 60784
rect 199200 60120 200000 60240
rect 199200 59032 200000 59152
rect 0 58760 800 58880
rect 199200 57944 200000 58064
rect 0 56856 800 56976
rect 199200 56856 200000 56976
rect 199200 55768 200000 55888
rect 0 54952 800 55072
rect 199200 54680 200000 54800
rect 199200 53592 200000 53712
rect 0 53048 800 53168
rect 199200 52504 200000 52624
rect 199200 51416 200000 51536
rect 0 51144 800 51264
rect 199200 50328 200000 50448
rect 0 49240 800 49360
rect 199200 49240 200000 49360
rect 199200 48152 200000 48272
rect 0 47336 800 47456
rect 199200 47064 200000 47184
rect 199200 45976 200000 46096
rect 0 45432 800 45552
rect 199200 44888 200000 45008
rect 199200 43800 200000 43920
rect 0 43528 800 43648
rect 199200 42712 200000 42832
rect 0 41624 800 41744
rect 199200 41624 200000 41744
rect 199200 40536 200000 40656
rect 0 39720 800 39840
rect 199200 39448 200000 39568
rect 199200 38360 200000 38480
rect 0 37816 800 37936
rect 199200 37272 200000 37392
rect 199200 36184 200000 36304
rect 0 35912 800 36032
rect 199200 35096 200000 35216
rect 0 34008 800 34128
rect 199200 34008 200000 34128
rect 199200 32920 200000 33040
rect 0 32104 800 32224
rect 199200 31832 200000 31952
rect 199200 30744 200000 30864
rect 0 30200 800 30320
rect 199200 29656 200000 29776
rect 199200 28568 200000 28688
rect 0 28296 800 28416
rect 199200 27480 200000 27600
rect 0 26392 800 26512
rect 199200 26392 200000 26512
rect 199200 25304 200000 25424
rect 0 24488 800 24608
rect 199200 24216 200000 24336
rect 199200 23128 200000 23248
rect 0 22584 800 22704
rect 199200 22040 200000 22160
rect 199200 20952 200000 21072
rect 0 20680 800 20800
rect 199200 19864 200000 19984
rect 0 18776 800 18896
rect 199200 18776 200000 18896
rect 199200 17688 200000 17808
rect 0 16872 800 16992
rect 199200 16600 200000 16720
rect 199200 15512 200000 15632
rect 0 14968 800 15088
rect 199200 14424 200000 14544
rect 199200 13336 200000 13456
rect 0 13064 800 13184
rect 0 11160 800 11280
rect 0 9256 800 9376
<< obsm3 >>
rect 798 190336 199200 197505
rect 880 190056 199200 190336
rect 798 188432 199200 190056
rect 880 188152 199200 188432
rect 798 186528 199200 188152
rect 880 186248 199120 186528
rect 798 185440 199200 186248
rect 798 185160 199120 185440
rect 798 184624 199200 185160
rect 880 184352 199200 184624
rect 880 184344 199120 184352
rect 798 184072 199120 184344
rect 798 183264 199200 184072
rect 798 182984 199120 183264
rect 798 182720 199200 182984
rect 880 182440 199200 182720
rect 798 182176 199200 182440
rect 798 181896 199120 182176
rect 798 181088 199200 181896
rect 798 180816 199120 181088
rect 880 180808 199120 180816
rect 880 180536 199200 180808
rect 798 180000 199200 180536
rect 798 179720 199120 180000
rect 798 178912 199200 179720
rect 880 178632 199120 178912
rect 798 177824 199200 178632
rect 798 177544 199120 177824
rect 798 177008 199200 177544
rect 880 176736 199200 177008
rect 880 176728 199120 176736
rect 798 176456 199120 176728
rect 798 175648 199200 176456
rect 798 175368 199120 175648
rect 798 175104 199200 175368
rect 880 174824 199200 175104
rect 798 174560 199200 174824
rect 798 174280 199120 174560
rect 798 173472 199200 174280
rect 798 173200 199120 173472
rect 880 173192 199120 173200
rect 880 172920 199200 173192
rect 798 172384 199200 172920
rect 798 172104 199120 172384
rect 798 171296 199200 172104
rect 880 171016 199120 171296
rect 798 170208 199200 171016
rect 798 169928 199120 170208
rect 798 169392 199200 169928
rect 880 169120 199200 169392
rect 880 169112 199120 169120
rect 798 168840 199120 169112
rect 798 168032 199200 168840
rect 798 167752 199120 168032
rect 798 167488 199200 167752
rect 880 167208 199200 167488
rect 798 166944 199200 167208
rect 798 166664 199120 166944
rect 798 165856 199200 166664
rect 798 165584 199120 165856
rect 880 165576 199120 165584
rect 880 165304 199200 165576
rect 798 164768 199200 165304
rect 798 164488 199120 164768
rect 798 163680 199200 164488
rect 880 163400 199120 163680
rect 798 162592 199200 163400
rect 798 162312 199120 162592
rect 798 161776 199200 162312
rect 880 161504 199200 161776
rect 880 161496 199120 161504
rect 798 161224 199120 161496
rect 798 160416 199200 161224
rect 798 160136 199120 160416
rect 798 159872 199200 160136
rect 880 159592 199200 159872
rect 798 159328 199200 159592
rect 798 159048 199120 159328
rect 798 158240 199200 159048
rect 798 157968 199120 158240
rect 880 157960 199120 157968
rect 880 157688 199200 157960
rect 798 157152 199200 157688
rect 798 156872 199120 157152
rect 798 156064 199200 156872
rect 880 155784 199120 156064
rect 798 154976 199200 155784
rect 798 154696 199120 154976
rect 798 154160 199200 154696
rect 880 153888 199200 154160
rect 880 153880 199120 153888
rect 798 153608 199120 153880
rect 798 152800 199200 153608
rect 798 152520 199120 152800
rect 798 152256 199200 152520
rect 880 151976 199200 152256
rect 798 151712 199200 151976
rect 798 151432 199120 151712
rect 798 150624 199200 151432
rect 798 150352 199120 150624
rect 880 150344 199120 150352
rect 880 150072 199200 150344
rect 798 149536 199200 150072
rect 798 149256 199120 149536
rect 798 148448 199200 149256
rect 880 148168 199120 148448
rect 798 147360 199200 148168
rect 798 147080 199120 147360
rect 798 146544 199200 147080
rect 880 146272 199200 146544
rect 880 146264 199120 146272
rect 798 145992 199120 146264
rect 798 145184 199200 145992
rect 798 144904 199120 145184
rect 798 144640 199200 144904
rect 880 144360 199200 144640
rect 798 144096 199200 144360
rect 798 143816 199120 144096
rect 798 143008 199200 143816
rect 798 142736 199120 143008
rect 880 142728 199120 142736
rect 880 142456 199200 142728
rect 798 141920 199200 142456
rect 798 141640 199120 141920
rect 798 140832 199200 141640
rect 880 140552 199120 140832
rect 798 139744 199200 140552
rect 798 139464 199120 139744
rect 798 138928 199200 139464
rect 880 138656 199200 138928
rect 880 138648 199120 138656
rect 798 138376 199120 138648
rect 798 137568 199200 138376
rect 798 137288 199120 137568
rect 798 137024 199200 137288
rect 880 136744 199200 137024
rect 798 136480 199200 136744
rect 798 136200 199120 136480
rect 798 135392 199200 136200
rect 798 135120 199120 135392
rect 880 135112 199120 135120
rect 880 134840 199200 135112
rect 798 134304 199200 134840
rect 798 134024 199120 134304
rect 798 133216 199200 134024
rect 880 132936 199120 133216
rect 798 132128 199200 132936
rect 798 131848 199120 132128
rect 798 131312 199200 131848
rect 880 131040 199200 131312
rect 880 131032 199120 131040
rect 798 130760 199120 131032
rect 798 129952 199200 130760
rect 798 129672 199120 129952
rect 798 129408 199200 129672
rect 880 129128 199200 129408
rect 798 128864 199200 129128
rect 798 128584 199120 128864
rect 798 127776 199200 128584
rect 798 127504 199120 127776
rect 880 127496 199120 127504
rect 880 127224 199200 127496
rect 798 126688 199200 127224
rect 798 126408 199120 126688
rect 798 125600 199200 126408
rect 880 125320 199120 125600
rect 798 124512 199200 125320
rect 798 124232 199120 124512
rect 798 123696 199200 124232
rect 880 123424 199200 123696
rect 880 123416 199120 123424
rect 798 123144 199120 123416
rect 798 122336 199200 123144
rect 798 122056 199120 122336
rect 798 121792 199200 122056
rect 880 121512 199200 121792
rect 798 121248 199200 121512
rect 798 120968 199120 121248
rect 798 120160 199200 120968
rect 798 119888 199120 120160
rect 880 119880 199120 119888
rect 880 119608 199200 119880
rect 798 119072 199200 119608
rect 798 118792 199120 119072
rect 798 117984 199200 118792
rect 880 117704 199120 117984
rect 798 116896 199200 117704
rect 798 116616 199120 116896
rect 798 116080 199200 116616
rect 880 115808 199200 116080
rect 880 115800 199120 115808
rect 798 115528 199120 115800
rect 798 114720 199200 115528
rect 798 114440 199120 114720
rect 798 114176 199200 114440
rect 880 113896 199200 114176
rect 798 113632 199200 113896
rect 798 113352 199120 113632
rect 798 112544 199200 113352
rect 798 112272 199120 112544
rect 880 112264 199120 112272
rect 880 111992 199200 112264
rect 798 111456 199200 111992
rect 798 111176 199120 111456
rect 798 110368 199200 111176
rect 880 110088 199120 110368
rect 798 109280 199200 110088
rect 798 109000 199120 109280
rect 798 108464 199200 109000
rect 880 108192 199200 108464
rect 880 108184 199120 108192
rect 798 107912 199120 108184
rect 798 107104 199200 107912
rect 798 106824 199120 107104
rect 798 106560 199200 106824
rect 880 106280 199200 106560
rect 798 106016 199200 106280
rect 798 105736 199120 106016
rect 798 104928 199200 105736
rect 798 104656 199120 104928
rect 880 104648 199120 104656
rect 880 104376 199200 104648
rect 798 103840 199200 104376
rect 798 103560 199120 103840
rect 798 102752 199200 103560
rect 880 102472 199120 102752
rect 798 101664 199200 102472
rect 798 101384 199120 101664
rect 798 100848 199200 101384
rect 880 100576 199200 100848
rect 880 100568 199120 100576
rect 798 100296 199120 100568
rect 798 99488 199200 100296
rect 798 99208 199120 99488
rect 798 98944 199200 99208
rect 880 98664 199200 98944
rect 798 98400 199200 98664
rect 798 98120 199120 98400
rect 798 97312 199200 98120
rect 798 97040 199120 97312
rect 880 97032 199120 97040
rect 880 96760 199200 97032
rect 798 96224 199200 96760
rect 798 95944 199120 96224
rect 798 95136 199200 95944
rect 880 94856 199120 95136
rect 798 94048 199200 94856
rect 798 93768 199120 94048
rect 798 93232 199200 93768
rect 880 92960 199200 93232
rect 880 92952 199120 92960
rect 798 92680 199120 92952
rect 798 91872 199200 92680
rect 798 91592 199120 91872
rect 798 91328 199200 91592
rect 880 91048 199200 91328
rect 798 90784 199200 91048
rect 798 90504 199120 90784
rect 798 89696 199200 90504
rect 798 89424 199120 89696
rect 880 89416 199120 89424
rect 880 89144 199200 89416
rect 798 88608 199200 89144
rect 798 88328 199120 88608
rect 798 87520 199200 88328
rect 880 87240 199120 87520
rect 798 86432 199200 87240
rect 798 86152 199120 86432
rect 798 85616 199200 86152
rect 880 85344 199200 85616
rect 880 85336 199120 85344
rect 798 85064 199120 85336
rect 798 84256 199200 85064
rect 798 83976 199120 84256
rect 798 83712 199200 83976
rect 880 83432 199200 83712
rect 798 83168 199200 83432
rect 798 82888 199120 83168
rect 798 82080 199200 82888
rect 798 81808 199120 82080
rect 880 81800 199120 81808
rect 880 81528 199200 81800
rect 798 80992 199200 81528
rect 798 80712 199120 80992
rect 798 79904 199200 80712
rect 880 79624 199120 79904
rect 798 78816 199200 79624
rect 798 78536 199120 78816
rect 798 78000 199200 78536
rect 880 77728 199200 78000
rect 880 77720 199120 77728
rect 798 77448 199120 77720
rect 798 76640 199200 77448
rect 798 76360 199120 76640
rect 798 76096 199200 76360
rect 880 75816 199200 76096
rect 798 75552 199200 75816
rect 798 75272 199120 75552
rect 798 74464 199200 75272
rect 798 74192 199120 74464
rect 880 74184 199120 74192
rect 880 73912 199200 74184
rect 798 73376 199200 73912
rect 798 73096 199120 73376
rect 798 72288 199200 73096
rect 880 72008 199120 72288
rect 798 71200 199200 72008
rect 798 70920 199120 71200
rect 798 70384 199200 70920
rect 880 70112 199200 70384
rect 880 70104 199120 70112
rect 798 69832 199120 70104
rect 798 69024 199200 69832
rect 798 68744 199120 69024
rect 798 68480 199200 68744
rect 880 68200 199200 68480
rect 798 67936 199200 68200
rect 798 67656 199120 67936
rect 798 66848 199200 67656
rect 798 66576 199120 66848
rect 880 66568 199120 66576
rect 880 66296 199200 66568
rect 798 65760 199200 66296
rect 798 65480 199120 65760
rect 798 64672 199200 65480
rect 880 64392 199120 64672
rect 798 63584 199200 64392
rect 798 63304 199120 63584
rect 798 62768 199200 63304
rect 880 62496 199200 62768
rect 880 62488 199120 62496
rect 798 62216 199120 62488
rect 798 61408 199200 62216
rect 798 61128 199120 61408
rect 798 60864 199200 61128
rect 880 60584 199200 60864
rect 798 60320 199200 60584
rect 798 60040 199120 60320
rect 798 59232 199200 60040
rect 798 58960 199120 59232
rect 880 58952 199120 58960
rect 880 58680 199200 58952
rect 798 58144 199200 58680
rect 798 57864 199120 58144
rect 798 57056 199200 57864
rect 880 56776 199120 57056
rect 798 55968 199200 56776
rect 798 55688 199120 55968
rect 798 55152 199200 55688
rect 880 54880 199200 55152
rect 880 54872 199120 54880
rect 798 54600 199120 54872
rect 798 53792 199200 54600
rect 798 53512 199120 53792
rect 798 53248 199200 53512
rect 880 52968 199200 53248
rect 798 52704 199200 52968
rect 798 52424 199120 52704
rect 798 51616 199200 52424
rect 798 51344 199120 51616
rect 880 51336 199120 51344
rect 880 51064 199200 51336
rect 798 50528 199200 51064
rect 798 50248 199120 50528
rect 798 49440 199200 50248
rect 880 49160 199120 49440
rect 798 48352 199200 49160
rect 798 48072 199120 48352
rect 798 47536 199200 48072
rect 880 47264 199200 47536
rect 880 47256 199120 47264
rect 798 46984 199120 47256
rect 798 46176 199200 46984
rect 798 45896 199120 46176
rect 798 45632 199200 45896
rect 880 45352 199200 45632
rect 798 45088 199200 45352
rect 798 44808 199120 45088
rect 798 44000 199200 44808
rect 798 43728 199120 44000
rect 880 43720 199120 43728
rect 880 43448 199200 43720
rect 798 42912 199200 43448
rect 798 42632 199120 42912
rect 798 41824 199200 42632
rect 880 41544 199120 41824
rect 798 40736 199200 41544
rect 798 40456 199120 40736
rect 798 39920 199200 40456
rect 880 39648 199200 39920
rect 880 39640 199120 39648
rect 798 39368 199120 39640
rect 798 38560 199200 39368
rect 798 38280 199120 38560
rect 798 38016 199200 38280
rect 880 37736 199200 38016
rect 798 37472 199200 37736
rect 798 37192 199120 37472
rect 798 36384 199200 37192
rect 798 36112 199120 36384
rect 880 36104 199120 36112
rect 880 35832 199200 36104
rect 798 35296 199200 35832
rect 798 35016 199120 35296
rect 798 34208 199200 35016
rect 880 33928 199120 34208
rect 798 33120 199200 33928
rect 798 32840 199120 33120
rect 798 32304 199200 32840
rect 880 32032 199200 32304
rect 880 32024 199120 32032
rect 798 31752 199120 32024
rect 798 30944 199200 31752
rect 798 30664 199120 30944
rect 798 30400 199200 30664
rect 880 30120 199200 30400
rect 798 29856 199200 30120
rect 798 29576 199120 29856
rect 798 28768 199200 29576
rect 798 28496 199120 28768
rect 880 28488 199120 28496
rect 880 28216 199200 28488
rect 798 27680 199200 28216
rect 798 27400 199120 27680
rect 798 26592 199200 27400
rect 880 26312 199120 26592
rect 798 25504 199200 26312
rect 798 25224 199120 25504
rect 798 24688 199200 25224
rect 880 24416 199200 24688
rect 880 24408 199120 24416
rect 798 24136 199120 24408
rect 798 23328 199200 24136
rect 798 23048 199120 23328
rect 798 22784 199200 23048
rect 880 22504 199200 22784
rect 798 22240 199200 22504
rect 798 21960 199120 22240
rect 798 21152 199200 21960
rect 798 20880 199120 21152
rect 880 20872 199120 20880
rect 880 20600 199200 20872
rect 798 20064 199200 20600
rect 798 19784 199120 20064
rect 798 18976 199200 19784
rect 880 18696 199120 18976
rect 798 17888 199200 18696
rect 798 17608 199120 17888
rect 798 17072 199200 17608
rect 880 16800 199200 17072
rect 880 16792 199120 16800
rect 798 16520 199120 16792
rect 798 15712 199200 16520
rect 798 15432 199120 15712
rect 798 15168 199200 15432
rect 880 14888 199200 15168
rect 798 14624 199200 14888
rect 798 14344 199120 14624
rect 798 13536 199200 14344
rect 798 13264 199120 13536
rect 880 13256 199120 13264
rect 880 12984 199200 13256
rect 798 11360 199200 12984
rect 880 11080 199200 11360
rect 798 9456 199200 11080
rect 880 9176 199200 9456
rect 798 2143 199200 9176
<< metal4 >>
rect 4208 2128 4528 197520
rect 19568 2128 19888 197520
rect 34928 2128 35248 197520
rect 50288 2128 50608 197520
rect 65648 2128 65968 197520
rect 81008 2128 81328 197520
rect 96368 2128 96688 197520
rect 111728 2128 112048 197520
rect 127088 2128 127408 197520
rect 142448 2128 142768 197520
rect 157808 2128 158128 197520
rect 173168 2128 173488 197520
rect 188528 2128 188848 197520
<< obsm4 >>
rect 2819 2347 4128 197165
rect 4608 2347 19488 197165
rect 19968 2347 34848 197165
rect 35328 2347 50208 197165
rect 50688 2347 65568 197165
rect 66048 2347 80928 197165
rect 81408 2347 96288 197165
rect 96768 2347 111648 197165
rect 112128 2347 127008 197165
rect 127488 2347 142368 197165
rect 142848 2347 146957 197165
<< labels >>
rlabel metal3 s 0 188232 800 188352 6 busy_o
port 1 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 clk_i
port 2 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 mport_i[0]
port 3 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 mport_i[10]
port 4 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 mport_i[11]
port 5 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 mport_i[12]
port 6 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 mport_i[13]
port 7 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 mport_i[14]
port 8 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 mport_i[15]
port 9 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 mport_i[16]
port 10 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 mport_i[17]
port 11 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 mport_i[18]
port 12 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 mport_i[19]
port 13 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 mport_i[1]
port 14 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 mport_i[20]
port 15 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 mport_i[21]
port 16 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 mport_i[22]
port 17 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 mport_i[23]
port 18 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 mport_i[24]
port 19 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 mport_i[25]
port 20 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 mport_i[26]
port 21 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 mport_i[27]
port 22 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 mport_i[28]
port 23 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 mport_i[29]
port 24 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 mport_i[2]
port 25 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 mport_i[30]
port 26 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 mport_i[31]
port 27 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 mport_i[32]
port 28 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 mport_i[33]
port 29 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 mport_i[3]
port 30 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 mport_i[4]
port 31 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 mport_i[5]
port 32 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 mport_i[6]
port 33 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 mport_i[7]
port 34 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 mport_i[8]
port 35 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 mport_i[9]
port 36 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 mport_o[0]
port 37 nsew signal output
rlabel metal3 s 0 96840 800 96960 6 mport_o[10]
port 38 nsew signal output
rlabel metal3 s 0 98744 800 98864 6 mport_o[11]
port 39 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 mport_o[12]
port 40 nsew signal output
rlabel metal3 s 0 102552 800 102672 6 mport_o[13]
port 41 nsew signal output
rlabel metal3 s 0 104456 800 104576 6 mport_o[14]
port 42 nsew signal output
rlabel metal3 s 0 106360 800 106480 6 mport_o[15]
port 43 nsew signal output
rlabel metal3 s 0 108264 800 108384 6 mport_o[16]
port 44 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 mport_o[17]
port 45 nsew signal output
rlabel metal3 s 0 112072 800 112192 6 mport_o[18]
port 46 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 mport_o[19]
port 47 nsew signal output
rlabel metal3 s 0 79704 800 79824 6 mport_o[1]
port 48 nsew signal output
rlabel metal3 s 0 115880 800 116000 6 mport_o[20]
port 49 nsew signal output
rlabel metal3 s 0 117784 800 117904 6 mport_o[21]
port 50 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 mport_o[22]
port 51 nsew signal output
rlabel metal3 s 0 121592 800 121712 6 mport_o[23]
port 52 nsew signal output
rlabel metal3 s 0 123496 800 123616 6 mport_o[24]
port 53 nsew signal output
rlabel metal3 s 0 125400 800 125520 6 mport_o[25]
port 54 nsew signal output
rlabel metal3 s 0 127304 800 127424 6 mport_o[26]
port 55 nsew signal output
rlabel metal3 s 0 129208 800 129328 6 mport_o[27]
port 56 nsew signal output
rlabel metal3 s 0 131112 800 131232 6 mport_o[28]
port 57 nsew signal output
rlabel metal3 s 0 133016 800 133136 6 mport_o[29]
port 58 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 mport_o[2]
port 59 nsew signal output
rlabel metal3 s 0 134920 800 135040 6 mport_o[30]
port 60 nsew signal output
rlabel metal3 s 0 136824 800 136944 6 mport_o[31]
port 61 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 mport_o[32]
port 62 nsew signal output
rlabel metal3 s 0 140632 800 140752 6 mport_o[33]
port 63 nsew signal output
rlabel metal3 s 0 142536 800 142656 6 mport_o[34]
port 64 nsew signal output
rlabel metal3 s 0 144440 800 144560 6 mport_o[35]
port 65 nsew signal output
rlabel metal3 s 0 146344 800 146464 6 mport_o[36]
port 66 nsew signal output
rlabel metal3 s 0 148248 800 148368 6 mport_o[37]
port 67 nsew signal output
rlabel metal3 s 0 150152 800 150272 6 mport_o[38]
port 68 nsew signal output
rlabel metal3 s 0 152056 800 152176 6 mport_o[39]
port 69 nsew signal output
rlabel metal3 s 0 83512 800 83632 6 mport_o[3]
port 70 nsew signal output
rlabel metal3 s 0 153960 800 154080 6 mport_o[40]
port 71 nsew signal output
rlabel metal3 s 0 155864 800 155984 6 mport_o[41]
port 72 nsew signal output
rlabel metal3 s 0 157768 800 157888 6 mport_o[42]
port 73 nsew signal output
rlabel metal3 s 0 159672 800 159792 6 mport_o[43]
port 74 nsew signal output
rlabel metal3 s 0 161576 800 161696 6 mport_o[44]
port 75 nsew signal output
rlabel metal3 s 0 163480 800 163600 6 mport_o[45]
port 76 nsew signal output
rlabel metal3 s 0 165384 800 165504 6 mport_o[46]
port 77 nsew signal output
rlabel metal3 s 0 167288 800 167408 6 mport_o[47]
port 78 nsew signal output
rlabel metal3 s 0 169192 800 169312 6 mport_o[48]
port 79 nsew signal output
rlabel metal3 s 0 171096 800 171216 6 mport_o[49]
port 80 nsew signal output
rlabel metal3 s 0 85416 800 85536 6 mport_o[4]
port 81 nsew signal output
rlabel metal3 s 0 173000 800 173120 6 mport_o[50]
port 82 nsew signal output
rlabel metal3 s 0 174904 800 175024 6 mport_o[51]
port 83 nsew signal output
rlabel metal3 s 0 176808 800 176928 6 mport_o[52]
port 84 nsew signal output
rlabel metal3 s 0 178712 800 178832 6 mport_o[53]
port 85 nsew signal output
rlabel metal3 s 0 180616 800 180736 6 mport_o[54]
port 86 nsew signal output
rlabel metal3 s 0 182520 800 182640 6 mport_o[55]
port 87 nsew signal output
rlabel metal3 s 0 184424 800 184544 6 mport_o[56]
port 88 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 mport_o[5]
port 89 nsew signal output
rlabel metal3 s 0 89224 800 89344 6 mport_o[6]
port 90 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 mport_o[7]
port 91 nsew signal output
rlabel metal3 s 0 93032 800 93152 6 mport_o[8]
port 92 nsew signal output
rlabel metal3 s 0 94936 800 95056 6 mport_o[9]
port 93 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 nrst_i
port 94 nsew signal input
rlabel metal3 s 0 190136 800 190256 6 output_ready_o
port 95 nsew signal output
rlabel metal3 s 0 186328 800 186448 6 run_i
port 96 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 t0x[0]
port 97 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 t0x[10]
port 98 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 t0x[11]
port 99 nsew signal input
rlabel metal2 s 148414 0 148470 800 6 t0x[12]
port 100 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 t0x[13]
port 101 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 t0x[14]
port 102 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 t0x[15]
port 103 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 t0x[16]
port 104 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 t0x[17]
port 105 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 t0x[18]
port 106 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 t0x[19]
port 107 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 t0x[1]
port 108 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 t0x[20]
port 109 nsew signal input
rlabel metal2 s 169942 0 169998 800 6 t0x[21]
port 110 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 t0x[22]
port 111 nsew signal input
rlabel metal2 s 174726 0 174782 800 6 t0x[23]
port 112 nsew signal input
rlabel metal2 s 177118 0 177174 800 6 t0x[24]
port 113 nsew signal input
rlabel metal2 s 179510 0 179566 800 6 t0x[25]
port 114 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 t0x[26]
port 115 nsew signal input
rlabel metal2 s 184294 0 184350 800 6 t0x[27]
port 116 nsew signal input
rlabel metal2 s 186686 0 186742 800 6 t0x[28]
port 117 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 t0x[29]
port 118 nsew signal input
rlabel metal2 s 124494 0 124550 800 6 t0x[2]
port 119 nsew signal input
rlabel metal2 s 191470 0 191526 800 6 t0x[30]
port 120 nsew signal input
rlabel metal2 s 193862 0 193918 800 6 t0x[31]
port 121 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 t0x[3]
port 122 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 t0x[4]
port 123 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 t0x[5]
port 124 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 t0x[6]
port 125 nsew signal input
rlabel metal2 s 136454 0 136510 800 6 t0x[7]
port 126 nsew signal input
rlabel metal2 s 138846 0 138902 800 6 t0x[8]
port 127 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 t0x[9]
port 128 nsew signal input
rlabel metal2 s 120906 0 120962 800 6 t0y[0]
port 129 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 t0y[10]
port 130 nsew signal input
rlabel metal2 s 147218 0 147274 800 6 t0y[11]
port 131 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 t0y[12]
port 132 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 t0y[13]
port 133 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 t0y[14]
port 134 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 t0y[15]
port 135 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 t0y[16]
port 136 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 t0y[17]
port 137 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 t0y[18]
port 138 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 t0y[19]
port 139 nsew signal input
rlabel metal2 s 123298 0 123354 800 6 t0y[1]
port 140 nsew signal input
rlabel metal2 s 168746 0 168802 800 6 t0y[20]
port 141 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 t0y[21]
port 142 nsew signal input
rlabel metal2 s 173530 0 173586 800 6 t0y[22]
port 143 nsew signal input
rlabel metal2 s 175922 0 175978 800 6 t0y[23]
port 144 nsew signal input
rlabel metal2 s 178314 0 178370 800 6 t0y[24]
port 145 nsew signal input
rlabel metal2 s 180706 0 180762 800 6 t0y[25]
port 146 nsew signal input
rlabel metal2 s 183098 0 183154 800 6 t0y[26]
port 147 nsew signal input
rlabel metal2 s 185490 0 185546 800 6 t0y[27]
port 148 nsew signal input
rlabel metal2 s 187882 0 187938 800 6 t0y[28]
port 149 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 t0y[29]
port 150 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 t0y[2]
port 151 nsew signal input
rlabel metal2 s 192666 0 192722 800 6 t0y[30]
port 152 nsew signal input
rlabel metal2 s 195058 0 195114 800 6 t0y[31]
port 153 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 t0y[3]
port 154 nsew signal input
rlabel metal2 s 130474 0 130530 800 6 t0y[4]
port 155 nsew signal input
rlabel metal2 s 132866 0 132922 800 6 t0y[5]
port 156 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 t0y[6]
port 157 nsew signal input
rlabel metal2 s 137650 0 137706 800 6 t0y[7]
port 158 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 t0y[8]
port 159 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 t0y[9]
port 160 nsew signal input
rlabel metal2 s 119710 199200 119766 200000 6 t1x[0]
port 161 nsew signal input
rlabel metal2 s 143630 199200 143686 200000 6 t1x[10]
port 162 nsew signal input
rlabel metal2 s 146022 199200 146078 200000 6 t1x[11]
port 163 nsew signal input
rlabel metal2 s 148414 199200 148470 200000 6 t1x[12]
port 164 nsew signal input
rlabel metal2 s 150806 199200 150862 200000 6 t1x[13]
port 165 nsew signal input
rlabel metal2 s 153198 199200 153254 200000 6 t1x[14]
port 166 nsew signal input
rlabel metal2 s 155590 199200 155646 200000 6 t1x[15]
port 167 nsew signal input
rlabel metal2 s 157982 199200 158038 200000 6 t1x[16]
port 168 nsew signal input
rlabel metal2 s 160374 199200 160430 200000 6 t1x[17]
port 169 nsew signal input
rlabel metal2 s 162766 199200 162822 200000 6 t1x[18]
port 170 nsew signal input
rlabel metal2 s 165158 199200 165214 200000 6 t1x[19]
port 171 nsew signal input
rlabel metal2 s 122102 199200 122158 200000 6 t1x[1]
port 172 nsew signal input
rlabel metal2 s 167550 199200 167606 200000 6 t1x[20]
port 173 nsew signal input
rlabel metal2 s 169942 199200 169998 200000 6 t1x[21]
port 174 nsew signal input
rlabel metal2 s 172334 199200 172390 200000 6 t1x[22]
port 175 nsew signal input
rlabel metal2 s 174726 199200 174782 200000 6 t1x[23]
port 176 nsew signal input
rlabel metal2 s 177118 199200 177174 200000 6 t1x[24]
port 177 nsew signal input
rlabel metal2 s 179510 199200 179566 200000 6 t1x[25]
port 178 nsew signal input
rlabel metal2 s 181902 199200 181958 200000 6 t1x[26]
port 179 nsew signal input
rlabel metal2 s 184294 199200 184350 200000 6 t1x[27]
port 180 nsew signal input
rlabel metal2 s 186686 199200 186742 200000 6 t1x[28]
port 181 nsew signal input
rlabel metal2 s 189078 199200 189134 200000 6 t1x[29]
port 182 nsew signal input
rlabel metal2 s 124494 199200 124550 200000 6 t1x[2]
port 183 nsew signal input
rlabel metal2 s 191470 199200 191526 200000 6 t1x[30]
port 184 nsew signal input
rlabel metal2 s 193862 199200 193918 200000 6 t1x[31]
port 185 nsew signal input
rlabel metal2 s 126886 199200 126942 200000 6 t1x[3]
port 186 nsew signal input
rlabel metal2 s 129278 199200 129334 200000 6 t1x[4]
port 187 nsew signal input
rlabel metal2 s 131670 199200 131726 200000 6 t1x[5]
port 188 nsew signal input
rlabel metal2 s 134062 199200 134118 200000 6 t1x[6]
port 189 nsew signal input
rlabel metal2 s 136454 199200 136510 200000 6 t1x[7]
port 190 nsew signal input
rlabel metal2 s 138846 199200 138902 200000 6 t1x[8]
port 191 nsew signal input
rlabel metal2 s 141238 199200 141294 200000 6 t1x[9]
port 192 nsew signal input
rlabel metal2 s 120906 199200 120962 200000 6 t1y[0]
port 193 nsew signal input
rlabel metal2 s 144826 199200 144882 200000 6 t1y[10]
port 194 nsew signal input
rlabel metal2 s 147218 199200 147274 200000 6 t1y[11]
port 195 nsew signal input
rlabel metal2 s 149610 199200 149666 200000 6 t1y[12]
port 196 nsew signal input
rlabel metal2 s 152002 199200 152058 200000 6 t1y[13]
port 197 nsew signal input
rlabel metal2 s 154394 199200 154450 200000 6 t1y[14]
port 198 nsew signal input
rlabel metal2 s 156786 199200 156842 200000 6 t1y[15]
port 199 nsew signal input
rlabel metal2 s 159178 199200 159234 200000 6 t1y[16]
port 200 nsew signal input
rlabel metal2 s 161570 199200 161626 200000 6 t1y[17]
port 201 nsew signal input
rlabel metal2 s 163962 199200 164018 200000 6 t1y[18]
port 202 nsew signal input
rlabel metal2 s 166354 199200 166410 200000 6 t1y[19]
port 203 nsew signal input
rlabel metal2 s 123298 199200 123354 200000 6 t1y[1]
port 204 nsew signal input
rlabel metal2 s 168746 199200 168802 200000 6 t1y[20]
port 205 nsew signal input
rlabel metal2 s 171138 199200 171194 200000 6 t1y[21]
port 206 nsew signal input
rlabel metal2 s 173530 199200 173586 200000 6 t1y[22]
port 207 nsew signal input
rlabel metal2 s 175922 199200 175978 200000 6 t1y[23]
port 208 nsew signal input
rlabel metal2 s 178314 199200 178370 200000 6 t1y[24]
port 209 nsew signal input
rlabel metal2 s 180706 199200 180762 200000 6 t1y[25]
port 210 nsew signal input
rlabel metal2 s 183098 199200 183154 200000 6 t1y[26]
port 211 nsew signal input
rlabel metal2 s 185490 199200 185546 200000 6 t1y[27]
port 212 nsew signal input
rlabel metal2 s 187882 199200 187938 200000 6 t1y[28]
port 213 nsew signal input
rlabel metal2 s 190274 199200 190330 200000 6 t1y[29]
port 214 nsew signal input
rlabel metal2 s 125690 199200 125746 200000 6 t1y[2]
port 215 nsew signal input
rlabel metal2 s 192666 199200 192722 200000 6 t1y[30]
port 216 nsew signal input
rlabel metal2 s 195058 199200 195114 200000 6 t1y[31]
port 217 nsew signal input
rlabel metal2 s 128082 199200 128138 200000 6 t1y[3]
port 218 nsew signal input
rlabel metal2 s 130474 199200 130530 200000 6 t1y[4]
port 219 nsew signal input
rlabel metal2 s 132866 199200 132922 200000 6 t1y[5]
port 220 nsew signal input
rlabel metal2 s 135258 199200 135314 200000 6 t1y[6]
port 221 nsew signal input
rlabel metal2 s 137650 199200 137706 200000 6 t1y[7]
port 222 nsew signal input
rlabel metal2 s 140042 199200 140098 200000 6 t1y[8]
port 223 nsew signal input
rlabel metal2 s 142434 199200 142490 200000 6 t1y[9]
port 224 nsew signal input
rlabel metal3 s 199200 117784 200000 117904 6 t2x[0]
port 225 nsew signal input
rlabel metal3 s 199200 139544 200000 139664 6 t2x[10]
port 226 nsew signal input
rlabel metal3 s 199200 141720 200000 141840 6 t2x[11]
port 227 nsew signal input
rlabel metal3 s 199200 143896 200000 144016 6 t2x[12]
port 228 nsew signal input
rlabel metal3 s 199200 146072 200000 146192 6 t2x[13]
port 229 nsew signal input
rlabel metal3 s 199200 148248 200000 148368 6 t2x[14]
port 230 nsew signal input
rlabel metal3 s 199200 150424 200000 150544 6 t2x[15]
port 231 nsew signal input
rlabel metal3 s 199200 152600 200000 152720 6 t2x[16]
port 232 nsew signal input
rlabel metal3 s 199200 154776 200000 154896 6 t2x[17]
port 233 nsew signal input
rlabel metal3 s 199200 156952 200000 157072 6 t2x[18]
port 234 nsew signal input
rlabel metal3 s 199200 159128 200000 159248 6 t2x[19]
port 235 nsew signal input
rlabel metal3 s 199200 119960 200000 120080 6 t2x[1]
port 236 nsew signal input
rlabel metal3 s 199200 161304 200000 161424 6 t2x[20]
port 237 nsew signal input
rlabel metal3 s 199200 163480 200000 163600 6 t2x[21]
port 238 nsew signal input
rlabel metal3 s 199200 165656 200000 165776 6 t2x[22]
port 239 nsew signal input
rlabel metal3 s 199200 167832 200000 167952 6 t2x[23]
port 240 nsew signal input
rlabel metal3 s 199200 170008 200000 170128 6 t2x[24]
port 241 nsew signal input
rlabel metal3 s 199200 172184 200000 172304 6 t2x[25]
port 242 nsew signal input
rlabel metal3 s 199200 174360 200000 174480 6 t2x[26]
port 243 nsew signal input
rlabel metal3 s 199200 176536 200000 176656 6 t2x[27]
port 244 nsew signal input
rlabel metal3 s 199200 178712 200000 178832 6 t2x[28]
port 245 nsew signal input
rlabel metal3 s 199200 180888 200000 181008 6 t2x[29]
port 246 nsew signal input
rlabel metal3 s 199200 122136 200000 122256 6 t2x[2]
port 247 nsew signal input
rlabel metal3 s 199200 183064 200000 183184 6 t2x[30]
port 248 nsew signal input
rlabel metal3 s 199200 185240 200000 185360 6 t2x[31]
port 249 nsew signal input
rlabel metal3 s 199200 124312 200000 124432 6 t2x[3]
port 250 nsew signal input
rlabel metal3 s 199200 126488 200000 126608 6 t2x[4]
port 251 nsew signal input
rlabel metal3 s 199200 128664 200000 128784 6 t2x[5]
port 252 nsew signal input
rlabel metal3 s 199200 130840 200000 130960 6 t2x[6]
port 253 nsew signal input
rlabel metal3 s 199200 133016 200000 133136 6 t2x[7]
port 254 nsew signal input
rlabel metal3 s 199200 135192 200000 135312 6 t2x[8]
port 255 nsew signal input
rlabel metal3 s 199200 137368 200000 137488 6 t2x[9]
port 256 nsew signal input
rlabel metal3 s 199200 118872 200000 118992 6 t2y[0]
port 257 nsew signal input
rlabel metal3 s 199200 140632 200000 140752 6 t2y[10]
port 258 nsew signal input
rlabel metal3 s 199200 142808 200000 142928 6 t2y[11]
port 259 nsew signal input
rlabel metal3 s 199200 144984 200000 145104 6 t2y[12]
port 260 nsew signal input
rlabel metal3 s 199200 147160 200000 147280 6 t2y[13]
port 261 nsew signal input
rlabel metal3 s 199200 149336 200000 149456 6 t2y[14]
port 262 nsew signal input
rlabel metal3 s 199200 151512 200000 151632 6 t2y[15]
port 263 nsew signal input
rlabel metal3 s 199200 153688 200000 153808 6 t2y[16]
port 264 nsew signal input
rlabel metal3 s 199200 155864 200000 155984 6 t2y[17]
port 265 nsew signal input
rlabel metal3 s 199200 158040 200000 158160 6 t2y[18]
port 266 nsew signal input
rlabel metal3 s 199200 160216 200000 160336 6 t2y[19]
port 267 nsew signal input
rlabel metal3 s 199200 121048 200000 121168 6 t2y[1]
port 268 nsew signal input
rlabel metal3 s 199200 162392 200000 162512 6 t2y[20]
port 269 nsew signal input
rlabel metal3 s 199200 164568 200000 164688 6 t2y[21]
port 270 nsew signal input
rlabel metal3 s 199200 166744 200000 166864 6 t2y[22]
port 271 nsew signal input
rlabel metal3 s 199200 168920 200000 169040 6 t2y[23]
port 272 nsew signal input
rlabel metal3 s 199200 171096 200000 171216 6 t2y[24]
port 273 nsew signal input
rlabel metal3 s 199200 173272 200000 173392 6 t2y[25]
port 274 nsew signal input
rlabel metal3 s 199200 175448 200000 175568 6 t2y[26]
port 275 nsew signal input
rlabel metal3 s 199200 177624 200000 177744 6 t2y[27]
port 276 nsew signal input
rlabel metal3 s 199200 179800 200000 179920 6 t2y[28]
port 277 nsew signal input
rlabel metal3 s 199200 181976 200000 182096 6 t2y[29]
port 278 nsew signal input
rlabel metal3 s 199200 123224 200000 123344 6 t2y[2]
port 279 nsew signal input
rlabel metal3 s 199200 184152 200000 184272 6 t2y[30]
port 280 nsew signal input
rlabel metal3 s 199200 186328 200000 186448 6 t2y[31]
port 281 nsew signal input
rlabel metal3 s 199200 125400 200000 125520 6 t2y[3]
port 282 nsew signal input
rlabel metal3 s 199200 127576 200000 127696 6 t2y[4]
port 283 nsew signal input
rlabel metal3 s 199200 129752 200000 129872 6 t2y[5]
port 284 nsew signal input
rlabel metal3 s 199200 131928 200000 132048 6 t2y[6]
port 285 nsew signal input
rlabel metal3 s 199200 134104 200000 134224 6 t2y[7]
port 286 nsew signal input
rlabel metal3 s 199200 136280 200000 136400 6 t2y[8]
port 287 nsew signal input
rlabel metal3 s 199200 138456 200000 138576 6 t2y[9]
port 288 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 v0x[0]
port 289 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 v0x[10]
port 290 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 v0x[11]
port 291 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 v0x[12]
port 292 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 v0x[13]
port 293 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 v0x[14]
port 294 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 v0x[15]
port 295 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 v0x[16]
port 296 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 v0x[17]
port 297 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 v0x[18]
port 298 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 v0x[19]
port 299 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 v0x[1]
port 300 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 v0x[20]
port 301 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 v0x[21]
port 302 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 v0x[22]
port 303 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 v0x[23]
port 304 nsew signal input
rlabel metal2 s 91006 0 91062 800 6 v0x[24]
port 305 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 v0x[25]
port 306 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 v0x[26]
port 307 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 v0x[27]
port 308 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 v0x[28]
port 309 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 v0x[29]
port 310 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 v0x[2]
port 311 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 v0x[30]
port 312 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 v0x[31]
port 313 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 v0x[3]
port 314 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 v0x[4]
port 315 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 v0x[5]
port 316 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 v0x[6]
port 317 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 v0x[7]
port 318 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 v0x[8]
port 319 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 v0x[9]
port 320 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 v0y[0]
port 321 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 v0y[10]
port 322 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 v0y[11]
port 323 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 v0y[12]
port 324 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 v0y[13]
port 325 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 v0y[14]
port 326 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 v0y[15]
port 327 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 v0y[16]
port 328 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 v0y[17]
port 329 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 v0y[18]
port 330 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 v0y[19]
port 331 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 v0y[1]
port 332 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 v0y[20]
port 333 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 v0y[21]
port 334 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 v0y[22]
port 335 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 v0y[23]
port 336 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 v0y[24]
port 337 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 v0y[25]
port 338 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 v0y[26]
port 339 nsew signal input
rlabel metal2 s 102966 0 103022 800 6 v0y[27]
port 340 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 v0y[28]
port 341 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 v0y[29]
port 342 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 v0y[2]
port 343 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 v0y[30]
port 344 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 v0y[31]
port 345 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 v0y[3]
port 346 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 v0y[4]
port 347 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 v0y[5]
port 348 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 v0y[6]
port 349 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 v0y[7]
port 350 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 v0y[8]
port 351 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 v0y[9]
port 352 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 v0z[0]
port 353 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 v0z[10]
port 354 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 v0z[11]
port 355 nsew signal input
rlabel metal2 s 50342 0 50398 800 6 v0z[12]
port 356 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 v0z[13]
port 357 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 v0z[14]
port 358 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 v0z[15]
port 359 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 v0z[16]
port 360 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 v0z[17]
port 361 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 v0z[18]
port 362 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 v0z[19]
port 363 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 v0z[1]
port 364 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 v0z[20]
port 365 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 v0z[21]
port 366 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 v0z[22]
port 367 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 v0z[23]
port 368 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 v0z[24]
port 369 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 v0z[25]
port 370 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 v0z[26]
port 371 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 v0z[27]
port 372 nsew signal input
rlabel metal2 s 107750 0 107806 800 6 v0z[28]
port 373 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 v0z[29]
port 374 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 v0z[2]
port 375 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 v0z[30]
port 376 nsew signal input
rlabel metal2 s 118514 0 118570 800 6 v0z[31]
port 377 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 v0z[3]
port 378 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 v0z[4]
port 379 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 v0z[5]
port 380 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 v0z[6]
port 381 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 v0z[7]
port 382 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 v0z[8]
port 383 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 v0z[9]
port 384 nsew signal input
rlabel metal2 s 4894 199200 4950 200000 6 v1x[0]
port 385 nsew signal input
rlabel metal2 s 40774 199200 40830 200000 6 v1x[10]
port 386 nsew signal input
rlabel metal2 s 44362 199200 44418 200000 6 v1x[11]
port 387 nsew signal input
rlabel metal2 s 47950 199200 48006 200000 6 v1x[12]
port 388 nsew signal input
rlabel metal2 s 51538 199200 51594 200000 6 v1x[13]
port 389 nsew signal input
rlabel metal2 s 55126 199200 55182 200000 6 v1x[14]
port 390 nsew signal input
rlabel metal2 s 58714 199200 58770 200000 6 v1x[15]
port 391 nsew signal input
rlabel metal2 s 62302 199200 62358 200000 6 v1x[16]
port 392 nsew signal input
rlabel metal2 s 65890 199200 65946 200000 6 v1x[17]
port 393 nsew signal input
rlabel metal2 s 69478 199200 69534 200000 6 v1x[18]
port 394 nsew signal input
rlabel metal2 s 73066 199200 73122 200000 6 v1x[19]
port 395 nsew signal input
rlabel metal2 s 8482 199200 8538 200000 6 v1x[1]
port 396 nsew signal input
rlabel metal2 s 76654 199200 76710 200000 6 v1x[20]
port 397 nsew signal input
rlabel metal2 s 80242 199200 80298 200000 6 v1x[21]
port 398 nsew signal input
rlabel metal2 s 83830 199200 83886 200000 6 v1x[22]
port 399 nsew signal input
rlabel metal2 s 87418 199200 87474 200000 6 v1x[23]
port 400 nsew signal input
rlabel metal2 s 91006 199200 91062 200000 6 v1x[24]
port 401 nsew signal input
rlabel metal2 s 94594 199200 94650 200000 6 v1x[25]
port 402 nsew signal input
rlabel metal2 s 98182 199200 98238 200000 6 v1x[26]
port 403 nsew signal input
rlabel metal2 s 101770 199200 101826 200000 6 v1x[27]
port 404 nsew signal input
rlabel metal2 s 105358 199200 105414 200000 6 v1x[28]
port 405 nsew signal input
rlabel metal2 s 108946 199200 109002 200000 6 v1x[29]
port 406 nsew signal input
rlabel metal2 s 12070 199200 12126 200000 6 v1x[2]
port 407 nsew signal input
rlabel metal2 s 112534 199200 112590 200000 6 v1x[30]
port 408 nsew signal input
rlabel metal2 s 116122 199200 116178 200000 6 v1x[31]
port 409 nsew signal input
rlabel metal2 s 15658 199200 15714 200000 6 v1x[3]
port 410 nsew signal input
rlabel metal2 s 19246 199200 19302 200000 6 v1x[4]
port 411 nsew signal input
rlabel metal2 s 22834 199200 22890 200000 6 v1x[5]
port 412 nsew signal input
rlabel metal2 s 26422 199200 26478 200000 6 v1x[6]
port 413 nsew signal input
rlabel metal2 s 30010 199200 30066 200000 6 v1x[7]
port 414 nsew signal input
rlabel metal2 s 33598 199200 33654 200000 6 v1x[8]
port 415 nsew signal input
rlabel metal2 s 37186 199200 37242 200000 6 v1x[9]
port 416 nsew signal input
rlabel metal2 s 6090 199200 6146 200000 6 v1y[0]
port 417 nsew signal input
rlabel metal2 s 41970 199200 42026 200000 6 v1y[10]
port 418 nsew signal input
rlabel metal2 s 45558 199200 45614 200000 6 v1y[11]
port 419 nsew signal input
rlabel metal2 s 49146 199200 49202 200000 6 v1y[12]
port 420 nsew signal input
rlabel metal2 s 52734 199200 52790 200000 6 v1y[13]
port 421 nsew signal input
rlabel metal2 s 56322 199200 56378 200000 6 v1y[14]
port 422 nsew signal input
rlabel metal2 s 59910 199200 59966 200000 6 v1y[15]
port 423 nsew signal input
rlabel metal2 s 63498 199200 63554 200000 6 v1y[16]
port 424 nsew signal input
rlabel metal2 s 67086 199200 67142 200000 6 v1y[17]
port 425 nsew signal input
rlabel metal2 s 70674 199200 70730 200000 6 v1y[18]
port 426 nsew signal input
rlabel metal2 s 74262 199200 74318 200000 6 v1y[19]
port 427 nsew signal input
rlabel metal2 s 9678 199200 9734 200000 6 v1y[1]
port 428 nsew signal input
rlabel metal2 s 77850 199200 77906 200000 6 v1y[20]
port 429 nsew signal input
rlabel metal2 s 81438 199200 81494 200000 6 v1y[21]
port 430 nsew signal input
rlabel metal2 s 85026 199200 85082 200000 6 v1y[22]
port 431 nsew signal input
rlabel metal2 s 88614 199200 88670 200000 6 v1y[23]
port 432 nsew signal input
rlabel metal2 s 92202 199200 92258 200000 6 v1y[24]
port 433 nsew signal input
rlabel metal2 s 95790 199200 95846 200000 6 v1y[25]
port 434 nsew signal input
rlabel metal2 s 99378 199200 99434 200000 6 v1y[26]
port 435 nsew signal input
rlabel metal2 s 102966 199200 103022 200000 6 v1y[27]
port 436 nsew signal input
rlabel metal2 s 106554 199200 106610 200000 6 v1y[28]
port 437 nsew signal input
rlabel metal2 s 110142 199200 110198 200000 6 v1y[29]
port 438 nsew signal input
rlabel metal2 s 13266 199200 13322 200000 6 v1y[2]
port 439 nsew signal input
rlabel metal2 s 113730 199200 113786 200000 6 v1y[30]
port 440 nsew signal input
rlabel metal2 s 117318 199200 117374 200000 6 v1y[31]
port 441 nsew signal input
rlabel metal2 s 16854 199200 16910 200000 6 v1y[3]
port 442 nsew signal input
rlabel metal2 s 20442 199200 20498 200000 6 v1y[4]
port 443 nsew signal input
rlabel metal2 s 24030 199200 24086 200000 6 v1y[5]
port 444 nsew signal input
rlabel metal2 s 27618 199200 27674 200000 6 v1y[6]
port 445 nsew signal input
rlabel metal2 s 31206 199200 31262 200000 6 v1y[7]
port 446 nsew signal input
rlabel metal2 s 34794 199200 34850 200000 6 v1y[8]
port 447 nsew signal input
rlabel metal2 s 38382 199200 38438 200000 6 v1y[9]
port 448 nsew signal input
rlabel metal2 s 7286 199200 7342 200000 6 v1z[0]
port 449 nsew signal input
rlabel metal2 s 43166 199200 43222 200000 6 v1z[10]
port 450 nsew signal input
rlabel metal2 s 46754 199200 46810 200000 6 v1z[11]
port 451 nsew signal input
rlabel metal2 s 50342 199200 50398 200000 6 v1z[12]
port 452 nsew signal input
rlabel metal2 s 53930 199200 53986 200000 6 v1z[13]
port 453 nsew signal input
rlabel metal2 s 57518 199200 57574 200000 6 v1z[14]
port 454 nsew signal input
rlabel metal2 s 61106 199200 61162 200000 6 v1z[15]
port 455 nsew signal input
rlabel metal2 s 64694 199200 64750 200000 6 v1z[16]
port 456 nsew signal input
rlabel metal2 s 68282 199200 68338 200000 6 v1z[17]
port 457 nsew signal input
rlabel metal2 s 71870 199200 71926 200000 6 v1z[18]
port 458 nsew signal input
rlabel metal2 s 75458 199200 75514 200000 6 v1z[19]
port 459 nsew signal input
rlabel metal2 s 10874 199200 10930 200000 6 v1z[1]
port 460 nsew signal input
rlabel metal2 s 79046 199200 79102 200000 6 v1z[20]
port 461 nsew signal input
rlabel metal2 s 82634 199200 82690 200000 6 v1z[21]
port 462 nsew signal input
rlabel metal2 s 86222 199200 86278 200000 6 v1z[22]
port 463 nsew signal input
rlabel metal2 s 89810 199200 89866 200000 6 v1z[23]
port 464 nsew signal input
rlabel metal2 s 93398 199200 93454 200000 6 v1z[24]
port 465 nsew signal input
rlabel metal2 s 96986 199200 97042 200000 6 v1z[25]
port 466 nsew signal input
rlabel metal2 s 100574 199200 100630 200000 6 v1z[26]
port 467 nsew signal input
rlabel metal2 s 104162 199200 104218 200000 6 v1z[27]
port 468 nsew signal input
rlabel metal2 s 107750 199200 107806 200000 6 v1z[28]
port 469 nsew signal input
rlabel metal2 s 111338 199200 111394 200000 6 v1z[29]
port 470 nsew signal input
rlabel metal2 s 14462 199200 14518 200000 6 v1z[2]
port 471 nsew signal input
rlabel metal2 s 114926 199200 114982 200000 6 v1z[30]
port 472 nsew signal input
rlabel metal2 s 118514 199200 118570 200000 6 v1z[31]
port 473 nsew signal input
rlabel metal2 s 18050 199200 18106 200000 6 v1z[3]
port 474 nsew signal input
rlabel metal2 s 21638 199200 21694 200000 6 v1z[4]
port 475 nsew signal input
rlabel metal2 s 25226 199200 25282 200000 6 v1z[5]
port 476 nsew signal input
rlabel metal2 s 28814 199200 28870 200000 6 v1z[6]
port 477 nsew signal input
rlabel metal2 s 32402 199200 32458 200000 6 v1z[7]
port 478 nsew signal input
rlabel metal2 s 35990 199200 36046 200000 6 v1z[8]
port 479 nsew signal input
rlabel metal2 s 39578 199200 39634 200000 6 v1z[9]
port 480 nsew signal input
rlabel metal3 s 199200 13336 200000 13456 6 v2x[0]
port 481 nsew signal input
rlabel metal3 s 199200 45976 200000 46096 6 v2x[10]
port 482 nsew signal input
rlabel metal3 s 199200 49240 200000 49360 6 v2x[11]
port 483 nsew signal input
rlabel metal3 s 199200 52504 200000 52624 6 v2x[12]
port 484 nsew signal input
rlabel metal3 s 199200 55768 200000 55888 6 v2x[13]
port 485 nsew signal input
rlabel metal3 s 199200 59032 200000 59152 6 v2x[14]
port 486 nsew signal input
rlabel metal3 s 199200 62296 200000 62416 6 v2x[15]
port 487 nsew signal input
rlabel metal3 s 199200 65560 200000 65680 6 v2x[16]
port 488 nsew signal input
rlabel metal3 s 199200 68824 200000 68944 6 v2x[17]
port 489 nsew signal input
rlabel metal3 s 199200 72088 200000 72208 6 v2x[18]
port 490 nsew signal input
rlabel metal3 s 199200 75352 200000 75472 6 v2x[19]
port 491 nsew signal input
rlabel metal3 s 199200 16600 200000 16720 6 v2x[1]
port 492 nsew signal input
rlabel metal3 s 199200 78616 200000 78736 6 v2x[20]
port 493 nsew signal input
rlabel metal3 s 199200 81880 200000 82000 6 v2x[21]
port 494 nsew signal input
rlabel metal3 s 199200 85144 200000 85264 6 v2x[22]
port 495 nsew signal input
rlabel metal3 s 199200 88408 200000 88528 6 v2x[23]
port 496 nsew signal input
rlabel metal3 s 199200 91672 200000 91792 6 v2x[24]
port 497 nsew signal input
rlabel metal3 s 199200 94936 200000 95056 6 v2x[25]
port 498 nsew signal input
rlabel metal3 s 199200 98200 200000 98320 6 v2x[26]
port 499 nsew signal input
rlabel metal3 s 199200 101464 200000 101584 6 v2x[27]
port 500 nsew signal input
rlabel metal3 s 199200 104728 200000 104848 6 v2x[28]
port 501 nsew signal input
rlabel metal3 s 199200 107992 200000 108112 6 v2x[29]
port 502 nsew signal input
rlabel metal3 s 199200 19864 200000 19984 6 v2x[2]
port 503 nsew signal input
rlabel metal3 s 199200 111256 200000 111376 6 v2x[30]
port 504 nsew signal input
rlabel metal3 s 199200 114520 200000 114640 6 v2x[31]
port 505 nsew signal input
rlabel metal3 s 199200 23128 200000 23248 6 v2x[3]
port 506 nsew signal input
rlabel metal3 s 199200 26392 200000 26512 6 v2x[4]
port 507 nsew signal input
rlabel metal3 s 199200 29656 200000 29776 6 v2x[5]
port 508 nsew signal input
rlabel metal3 s 199200 32920 200000 33040 6 v2x[6]
port 509 nsew signal input
rlabel metal3 s 199200 36184 200000 36304 6 v2x[7]
port 510 nsew signal input
rlabel metal3 s 199200 39448 200000 39568 6 v2x[8]
port 511 nsew signal input
rlabel metal3 s 199200 42712 200000 42832 6 v2x[9]
port 512 nsew signal input
rlabel metal3 s 199200 14424 200000 14544 6 v2y[0]
port 513 nsew signal input
rlabel metal3 s 199200 47064 200000 47184 6 v2y[10]
port 514 nsew signal input
rlabel metal3 s 199200 50328 200000 50448 6 v2y[11]
port 515 nsew signal input
rlabel metal3 s 199200 53592 200000 53712 6 v2y[12]
port 516 nsew signal input
rlabel metal3 s 199200 56856 200000 56976 6 v2y[13]
port 517 nsew signal input
rlabel metal3 s 199200 60120 200000 60240 6 v2y[14]
port 518 nsew signal input
rlabel metal3 s 199200 63384 200000 63504 6 v2y[15]
port 519 nsew signal input
rlabel metal3 s 199200 66648 200000 66768 6 v2y[16]
port 520 nsew signal input
rlabel metal3 s 199200 69912 200000 70032 6 v2y[17]
port 521 nsew signal input
rlabel metal3 s 199200 73176 200000 73296 6 v2y[18]
port 522 nsew signal input
rlabel metal3 s 199200 76440 200000 76560 6 v2y[19]
port 523 nsew signal input
rlabel metal3 s 199200 17688 200000 17808 6 v2y[1]
port 524 nsew signal input
rlabel metal3 s 199200 79704 200000 79824 6 v2y[20]
port 525 nsew signal input
rlabel metal3 s 199200 82968 200000 83088 6 v2y[21]
port 526 nsew signal input
rlabel metal3 s 199200 86232 200000 86352 6 v2y[22]
port 527 nsew signal input
rlabel metal3 s 199200 89496 200000 89616 6 v2y[23]
port 528 nsew signal input
rlabel metal3 s 199200 92760 200000 92880 6 v2y[24]
port 529 nsew signal input
rlabel metal3 s 199200 96024 200000 96144 6 v2y[25]
port 530 nsew signal input
rlabel metal3 s 199200 99288 200000 99408 6 v2y[26]
port 531 nsew signal input
rlabel metal3 s 199200 102552 200000 102672 6 v2y[27]
port 532 nsew signal input
rlabel metal3 s 199200 105816 200000 105936 6 v2y[28]
port 533 nsew signal input
rlabel metal3 s 199200 109080 200000 109200 6 v2y[29]
port 534 nsew signal input
rlabel metal3 s 199200 20952 200000 21072 6 v2y[2]
port 535 nsew signal input
rlabel metal3 s 199200 112344 200000 112464 6 v2y[30]
port 536 nsew signal input
rlabel metal3 s 199200 115608 200000 115728 6 v2y[31]
port 537 nsew signal input
rlabel metal3 s 199200 24216 200000 24336 6 v2y[3]
port 538 nsew signal input
rlabel metal3 s 199200 27480 200000 27600 6 v2y[4]
port 539 nsew signal input
rlabel metal3 s 199200 30744 200000 30864 6 v2y[5]
port 540 nsew signal input
rlabel metal3 s 199200 34008 200000 34128 6 v2y[6]
port 541 nsew signal input
rlabel metal3 s 199200 37272 200000 37392 6 v2y[7]
port 542 nsew signal input
rlabel metal3 s 199200 40536 200000 40656 6 v2y[8]
port 543 nsew signal input
rlabel metal3 s 199200 43800 200000 43920 6 v2y[9]
port 544 nsew signal input
rlabel metal3 s 199200 15512 200000 15632 6 v2z[0]
port 545 nsew signal input
rlabel metal3 s 199200 48152 200000 48272 6 v2z[10]
port 546 nsew signal input
rlabel metal3 s 199200 51416 200000 51536 6 v2z[11]
port 547 nsew signal input
rlabel metal3 s 199200 54680 200000 54800 6 v2z[12]
port 548 nsew signal input
rlabel metal3 s 199200 57944 200000 58064 6 v2z[13]
port 549 nsew signal input
rlabel metal3 s 199200 61208 200000 61328 6 v2z[14]
port 550 nsew signal input
rlabel metal3 s 199200 64472 200000 64592 6 v2z[15]
port 551 nsew signal input
rlabel metal3 s 199200 67736 200000 67856 6 v2z[16]
port 552 nsew signal input
rlabel metal3 s 199200 71000 200000 71120 6 v2z[17]
port 553 nsew signal input
rlabel metal3 s 199200 74264 200000 74384 6 v2z[18]
port 554 nsew signal input
rlabel metal3 s 199200 77528 200000 77648 6 v2z[19]
port 555 nsew signal input
rlabel metal3 s 199200 18776 200000 18896 6 v2z[1]
port 556 nsew signal input
rlabel metal3 s 199200 80792 200000 80912 6 v2z[20]
port 557 nsew signal input
rlabel metal3 s 199200 84056 200000 84176 6 v2z[21]
port 558 nsew signal input
rlabel metal3 s 199200 87320 200000 87440 6 v2z[22]
port 559 nsew signal input
rlabel metal3 s 199200 90584 200000 90704 6 v2z[23]
port 560 nsew signal input
rlabel metal3 s 199200 93848 200000 93968 6 v2z[24]
port 561 nsew signal input
rlabel metal3 s 199200 97112 200000 97232 6 v2z[25]
port 562 nsew signal input
rlabel metal3 s 199200 100376 200000 100496 6 v2z[26]
port 563 nsew signal input
rlabel metal3 s 199200 103640 200000 103760 6 v2z[27]
port 564 nsew signal input
rlabel metal3 s 199200 106904 200000 107024 6 v2z[28]
port 565 nsew signal input
rlabel metal3 s 199200 110168 200000 110288 6 v2z[29]
port 566 nsew signal input
rlabel metal3 s 199200 22040 200000 22160 6 v2z[2]
port 567 nsew signal input
rlabel metal3 s 199200 113432 200000 113552 6 v2z[30]
port 568 nsew signal input
rlabel metal3 s 199200 116696 200000 116816 6 v2z[31]
port 569 nsew signal input
rlabel metal3 s 199200 25304 200000 25424 6 v2z[3]
port 570 nsew signal input
rlabel metal3 s 199200 28568 200000 28688 6 v2z[4]
port 571 nsew signal input
rlabel metal3 s 199200 31832 200000 31952 6 v2z[5]
port 572 nsew signal input
rlabel metal3 s 199200 35096 200000 35216 6 v2z[6]
port 573 nsew signal input
rlabel metal3 s 199200 38360 200000 38480 6 v2z[7]
port 574 nsew signal input
rlabel metal3 s 199200 41624 200000 41744 6 v2z[8]
port 575 nsew signal input
rlabel metal3 s 199200 44888 200000 45008 6 v2z[9]
port 576 nsew signal input
rlabel metal4 s 4208 2128 4528 197520 6 vccd1
port 577 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 197520 6 vccd1
port 577 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 197520 6 vccd1
port 577 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 197520 6 vccd1
port 577 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 197520 6 vccd1
port 577 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 197520 6 vccd1
port 577 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 197520 6 vccd1
port 577 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 197520 6 vssd1
port 578 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 197520 6 vssd1
port 578 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 197520 6 vssd1
port 578 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 197520 6 vssd1
port 578 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 197520 6 vssd1
port 578 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 197520 6 vssd1
port 578 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 200000 200000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 61558854
string GDS_FILE /local/colinm22/sdmay26-24/openlane/rasterizer/runs/25_10_06_09_59/results/signoff/rasterizer_m.magic.gds
string GDS_START 997486
<< end >>

