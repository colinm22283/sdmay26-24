module vga_tb();

endmodule
