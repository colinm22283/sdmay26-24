VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rasterizer_m
  CLASS BLOCK ;
  FOREIGN rasterizer_m ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN busy_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 941.160 4.000 941.760 ;
    END
  END busy_o
  PIN clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END clk_i
  PIN mport_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END mport_i[0]
  PIN mport_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END mport_i[10]
  PIN mport_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END mport_i[11]
  PIN mport_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END mport_i[12]
  PIN mport_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END mport_i[13]
  PIN mport_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END mport_i[14]
  PIN mport_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END mport_i[15]
  PIN mport_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END mport_i[16]
  PIN mport_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END mport_i[17]
  PIN mport_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END mport_i[18]
  PIN mport_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.200 4.000 246.800 ;
    END
  END mport_i[19]
  PIN mport_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END mport_i[1]
  PIN mport_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END mport_i[20]
  PIN mport_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END mport_i[21]
  PIN mport_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END mport_i[22]
  PIN mport_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END mport_i[23]
  PIN mport_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.800 4.000 294.400 ;
    END
  END mport_i[24]
  PIN mport_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END mport_i[25]
  PIN mport_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END mport_i[26]
  PIN mport_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END mport_i[27]
  PIN mport_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END mport_i[28]
  PIN mport_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END mport_i[29]
  PIN mport_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END mport_i[2]
  PIN mport_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END mport_i[30]
  PIN mport_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END mport_i[31]
  PIN mport_i[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END mport_i[32]
  PIN mport_i[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END mport_i[33]
  PIN mport_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END mport_i[3]
  PIN mport_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END mport_i[4]
  PIN mport_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END mport_i[5]
  PIN mport_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END mport_i[6]
  PIN mport_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.960 4.000 132.560 ;
    END
  END mport_i[7]
  PIN mport_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 141.480 4.000 142.080 ;
    END
  END mport_i[8]
  PIN mport_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END mport_i[9]
  PIN mport_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END mport_o[0]
  PIN mport_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END mport_o[10]
  PIN mport_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END mport_o[11]
  PIN mport_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END mport_o[12]
  PIN mport_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END mport_o[13]
  PIN mport_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END mport_o[14]
  PIN mport_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 531.800 4.000 532.400 ;
    END
  END mport_o[15]
  PIN mport_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END mport_o[16]
  PIN mport_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END mport_o[17]
  PIN mport_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 560.360 4.000 560.960 ;
    END
  END mport_o[18]
  PIN mport_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.880 4.000 570.480 ;
    END
  END mport_o[19]
  PIN mport_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END mport_o[1]
  PIN mport_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END mport_o[20]
  PIN mport_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.920 4.000 589.520 ;
    END
  END mport_o[21]
  PIN mport_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END mport_o[22]
  PIN mport_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END mport_o[23]
  PIN mport_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END mport_o[24]
  PIN mport_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END mport_o[25]
  PIN mport_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END mport_o[26]
  PIN mport_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END mport_o[27]
  PIN mport_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END mport_o[28]
  PIN mport_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.080 4.000 665.680 ;
    END
  END mport_o[29]
  PIN mport_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END mport_o[2]
  PIN mport_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 674.600 4.000 675.200 ;
    END
  END mport_o[30]
  PIN mport_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END mport_o[31]
  PIN mport_o[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 693.640 4.000 694.240 ;
    END
  END mport_o[32]
  PIN mport_o[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.160 4.000 703.760 ;
    END
  END mport_o[33]
  PIN mport_o[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 4.000 713.280 ;
    END
  END mport_o[34]
  PIN mport_o[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END mport_o[35]
  PIN mport_o[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.720 4.000 732.320 ;
    END
  END mport_o[36]
  PIN mport_o[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END mport_o[37]
  PIN mport_o[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.760 4.000 751.360 ;
    END
  END mport_o[38]
  PIN mport_o[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 760.280 4.000 760.880 ;
    END
  END mport_o[39]
  PIN mport_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END mport_o[3]
  PIN mport_o[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END mport_o[40]
  PIN mport_o[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 779.320 4.000 779.920 ;
    END
  END mport_o[41]
  PIN mport_o[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END mport_o[42]
  PIN mport_o[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 798.360 4.000 798.960 ;
    END
  END mport_o[43]
  PIN mport_o[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 807.880 4.000 808.480 ;
    END
  END mport_o[44]
  PIN mport_o[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 817.400 4.000 818.000 ;
    END
  END mport_o[45]
  PIN mport_o[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.920 4.000 827.520 ;
    END
  END mport_o[46]
  PIN mport_o[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 836.440 4.000 837.040 ;
    END
  END mport_o[47]
  PIN mport_o[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 845.960 4.000 846.560 ;
    END
  END mport_o[48]
  PIN mport_o[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 855.480 4.000 856.080 ;
    END
  END mport_o[49]
  PIN mport_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END mport_o[4]
  PIN mport_o[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 865.000 4.000 865.600 ;
    END
  END mport_o[50]
  PIN mport_o[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 874.520 4.000 875.120 ;
    END
  END mport_o[51]
  PIN mport_o[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 884.040 4.000 884.640 ;
    END
  END mport_o[52]
  PIN mport_o[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 893.560 4.000 894.160 ;
    END
  END mport_o[53]
  PIN mport_o[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 903.080 4.000 903.680 ;
    END
  END mport_o[54]
  PIN mport_o[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 912.600 4.000 913.200 ;
    END
  END mport_o[55]
  PIN mport_o[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 922.120 4.000 922.720 ;
    END
  END mport_o[56]
  PIN mport_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END mport_o[5]
  PIN mport_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END mport_o[6]
  PIN mport_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END mport_o[7]
  PIN mport_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.160 4.000 465.760 ;
    END
  END mport_o[8]
  PIN mport_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END mport_o[9]
  PIN nrst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END nrst_i
  PIN output_ready_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 950.680 4.000 951.280 ;
    END
  END output_ready_o
  PIN run_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 931.640 4.000 932.240 ;
    END
  END run_i
  PIN t0x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 0.000 598.830 4.000 ;
    END
  END t0x[0]
  PIN t0x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 0.000 718.430 4.000 ;
    END
  END t0x[10]
  PIN t0x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END t0x[11]
  PIN t0x[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 0.000 742.350 4.000 ;
    END
  END t0x[12]
  PIN t0x[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 4.000 ;
    END
  END t0x[13]
  PIN t0x[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END t0x[14]
  PIN t0x[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END t0x[15]
  PIN t0x[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 0.000 790.190 4.000 ;
    END
  END t0x[16]
  PIN t0x[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END t0x[17]
  PIN t0x[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 0.000 814.110 4.000 ;
    END
  END t0x[18]
  PIN t0x[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 0.000 826.070 4.000 ;
    END
  END t0x[19]
  PIN t0x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END t0x[1]
  PIN t0x[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 0.000 838.030 4.000 ;
    END
  END t0x[20]
  PIN t0x[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 0.000 849.990 4.000 ;
    END
  END t0x[21]
  PIN t0x[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 0.000 861.950 4.000 ;
    END
  END t0x[22]
  PIN t0x[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 0.000 873.910 4.000 ;
    END
  END t0x[23]
  PIN t0x[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 0.000 885.870 4.000 ;
    END
  END t0x[24]
  PIN t0x[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 0.000 897.830 4.000 ;
    END
  END t0x[25]
  PIN t0x[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 0.000 909.790 4.000 ;
    END
  END t0x[26]
  PIN t0x[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 0.000 921.750 4.000 ;
    END
  END t0x[27]
  PIN t0x[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 0.000 933.710 4.000 ;
    END
  END t0x[28]
  PIN t0x[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.390 0.000 945.670 4.000 ;
    END
  END t0x[29]
  PIN t0x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END t0x[2]
  PIN t0x[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 0.000 957.630 4.000 ;
    END
  END t0x[30]
  PIN t0x[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 0.000 969.590 4.000 ;
    END
  END t0x[31]
  PIN t0x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END t0x[3]
  PIN t0x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END t0x[4]
  PIN t0x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 0.000 658.630 4.000 ;
    END
  END t0x[5]
  PIN t0x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END t0x[6]
  PIN t0x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 0.000 682.550 4.000 ;
    END
  END t0x[7]
  PIN t0x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END t0x[8]
  PIN t0x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END t0x[9]
  PIN t0y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END t0y[0]
  PIN t0y[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 0.000 724.410 4.000 ;
    END
  END t0y[10]
  PIN t0y[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 0.000 736.370 4.000 ;
    END
  END t0y[11]
  PIN t0y[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 4.000 ;
    END
  END t0y[12]
  PIN t0y[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END t0y[13]
  PIN t0y[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 0.000 772.250 4.000 ;
    END
  END t0y[14]
  PIN t0y[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 0.000 784.210 4.000 ;
    END
  END t0y[15]
  PIN t0y[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END t0y[16]
  PIN t0y[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 0.000 808.130 4.000 ;
    END
  END t0y[17]
  PIN t0y[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END t0y[18]
  PIN t0y[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.770 0.000 832.050 4.000 ;
    END
  END t0y[19]
  PIN t0y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END t0y[1]
  PIN t0y[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 0.000 844.010 4.000 ;
    END
  END t0y[20]
  PIN t0y[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 0.000 855.970 4.000 ;
    END
  END t0y[21]
  PIN t0y[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.650 0.000 867.930 4.000 ;
    END
  END t0y[22]
  PIN t0y[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 0.000 879.890 4.000 ;
    END
  END t0y[23]
  PIN t0y[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 0.000 891.850 4.000 ;
    END
  END t0y[24]
  PIN t0y[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.530 0.000 903.810 4.000 ;
    END
  END t0y[25]
  PIN t0y[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.490 0.000 915.770 4.000 ;
    END
  END t0y[26]
  PIN t0y[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 0.000 927.730 4.000 ;
    END
  END t0y[27]
  PIN t0y[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.410 0.000 939.690 4.000 ;
    END
  END t0y[28]
  PIN t0y[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 0.000 951.650 4.000 ;
    END
  END t0y[29]
  PIN t0y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 0.000 628.730 4.000 ;
    END
  END t0y[2]
  PIN t0y[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.330 0.000 963.610 4.000 ;
    END
  END t0y[30]
  PIN t0y[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 0.000 975.570 4.000 ;
    END
  END t0y[31]
  PIN t0y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END t0y[3]
  PIN t0y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 0.000 652.650 4.000 ;
    END
  END t0y[4]
  PIN t0y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 0.000 664.610 4.000 ;
    END
  END t0y[5]
  PIN t0y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END t0y[6]
  PIN t0y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 0.000 688.530 4.000 ;
    END
  END t0y[7]
  PIN t0y[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END t0y[8]
  PIN t0y[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 0.000 712.450 4.000 ;
    END
  END t0y[9]
  PIN t1x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 996.000 598.830 1000.000 ;
    END
  END t1x[0]
  PIN t1x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 996.000 718.430 1000.000 ;
    END
  END t1x[10]
  PIN t1x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 996.000 730.390 1000.000 ;
    END
  END t1x[11]
  PIN t1x[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 996.000 742.350 1000.000 ;
    END
  END t1x[12]
  PIN t1x[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 996.000 754.310 1000.000 ;
    END
  END t1x[13]
  PIN t1x[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 996.000 766.270 1000.000 ;
    END
  END t1x[14]
  PIN t1x[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 996.000 778.230 1000.000 ;
    END
  END t1x[15]
  PIN t1x[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 996.000 790.190 1000.000 ;
    END
  END t1x[16]
  PIN t1x[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 996.000 802.150 1000.000 ;
    END
  END t1x[17]
  PIN t1x[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 996.000 814.110 1000.000 ;
    END
  END t1x[18]
  PIN t1x[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.790 996.000 826.070 1000.000 ;
    END
  END t1x[19]
  PIN t1x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 996.000 610.790 1000.000 ;
    END
  END t1x[1]
  PIN t1x[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 996.000 838.030 1000.000 ;
    END
  END t1x[20]
  PIN t1x[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.710 996.000 849.990 1000.000 ;
    END
  END t1x[21]
  PIN t1x[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 996.000 861.950 1000.000 ;
    END
  END t1x[22]
  PIN t1x[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.630 996.000 873.910 1000.000 ;
    END
  END t1x[23]
  PIN t1x[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 996.000 885.870 1000.000 ;
    END
  END t1x[24]
  PIN t1x[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.550 996.000 897.830 1000.000 ;
    END
  END t1x[25]
  PIN t1x[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.510 996.000 909.790 1000.000 ;
    END
  END t1x[26]
  PIN t1x[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 996.000 921.750 1000.000 ;
    END
  END t1x[27]
  PIN t1x[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 996.000 933.710 1000.000 ;
    END
  END t1x[28]
  PIN t1x[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.390 996.000 945.670 1000.000 ;
    END
  END t1x[29]
  PIN t1x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 996.000 622.750 1000.000 ;
    END
  END t1x[2]
  PIN t1x[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 996.000 957.630 1000.000 ;
    END
  END t1x[30]
  PIN t1x[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 969.310 996.000 969.590 1000.000 ;
    END
  END t1x[31]
  PIN t1x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 996.000 634.710 1000.000 ;
    END
  END t1x[3]
  PIN t1x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 996.000 646.670 1000.000 ;
    END
  END t1x[4]
  PIN t1x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 996.000 658.630 1000.000 ;
    END
  END t1x[5]
  PIN t1x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 996.000 670.590 1000.000 ;
    END
  END t1x[6]
  PIN t1x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.270 996.000 682.550 1000.000 ;
    END
  END t1x[7]
  PIN t1x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 996.000 694.510 1000.000 ;
    END
  END t1x[8]
  PIN t1x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 996.000 706.470 1000.000 ;
    END
  END t1x[9]
  PIN t1y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.530 996.000 604.810 1000.000 ;
    END
  END t1y[0]
  PIN t1y[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 996.000 724.410 1000.000 ;
    END
  END t1y[10]
  PIN t1y[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 996.000 736.370 1000.000 ;
    END
  END t1y[11]
  PIN t1y[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 996.000 748.330 1000.000 ;
    END
  END t1y[12]
  PIN t1y[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 996.000 760.290 1000.000 ;
    END
  END t1y[13]
  PIN t1y[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 996.000 772.250 1000.000 ;
    END
  END t1y[14]
  PIN t1y[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 996.000 784.210 1000.000 ;
    END
  END t1y[15]
  PIN t1y[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 996.000 796.170 1000.000 ;
    END
  END t1y[16]
  PIN t1y[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 996.000 808.130 1000.000 ;
    END
  END t1y[17]
  PIN t1y[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 996.000 820.090 1000.000 ;
    END
  END t1y[18]
  PIN t1y[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.770 996.000 832.050 1000.000 ;
    END
  END t1y[19]
  PIN t1y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.490 996.000 616.770 1000.000 ;
    END
  END t1y[1]
  PIN t1y[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 996.000 844.010 1000.000 ;
    END
  END t1y[20]
  PIN t1y[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.690 996.000 855.970 1000.000 ;
    END
  END t1y[21]
  PIN t1y[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.650 996.000 867.930 1000.000 ;
    END
  END t1y[22]
  PIN t1y[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.610 996.000 879.890 1000.000 ;
    END
  END t1y[23]
  PIN t1y[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 996.000 891.850 1000.000 ;
    END
  END t1y[24]
  PIN t1y[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.530 996.000 903.810 1000.000 ;
    END
  END t1y[25]
  PIN t1y[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.490 996.000 915.770 1000.000 ;
    END
  END t1y[26]
  PIN t1y[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.450 996.000 927.730 1000.000 ;
    END
  END t1y[27]
  PIN t1y[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.410 996.000 939.690 1000.000 ;
    END
  END t1y[28]
  PIN t1y[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 996.000 951.650 1000.000 ;
    END
  END t1y[29]
  PIN t1y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 996.000 628.730 1000.000 ;
    END
  END t1y[2]
  PIN t1y[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.330 996.000 963.610 1000.000 ;
    END
  END t1y[30]
  PIN t1y[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 975.290 996.000 975.570 1000.000 ;
    END
  END t1y[31]
  PIN t1y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 996.000 640.690 1000.000 ;
    END
  END t1y[3]
  PIN t1y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.370 996.000 652.650 1000.000 ;
    END
  END t1y[4]
  PIN t1y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 996.000 664.610 1000.000 ;
    END
  END t1y[5]
  PIN t1y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 996.000 676.570 1000.000 ;
    END
  END t1y[6]
  PIN t1y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 996.000 688.530 1000.000 ;
    END
  END t1y[7]
  PIN t1y[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 996.000 700.490 1000.000 ;
    END
  END t1y[8]
  PIN t1y[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 996.000 712.450 1000.000 ;
    END
  END t1y[9]
  PIN t2x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 588.920 1000.000 589.520 ;
    END
  END t2x[0]
  PIN t2x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 697.720 1000.000 698.320 ;
    END
  END t2x[10]
  PIN t2x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 708.600 1000.000 709.200 ;
    END
  END t2x[11]
  PIN t2x[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 719.480 1000.000 720.080 ;
    END
  END t2x[12]
  PIN t2x[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 730.360 1000.000 730.960 ;
    END
  END t2x[13]
  PIN t2x[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 741.240 1000.000 741.840 ;
    END
  END t2x[14]
  PIN t2x[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 752.120 1000.000 752.720 ;
    END
  END t2x[15]
  PIN t2x[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 763.000 1000.000 763.600 ;
    END
  END t2x[16]
  PIN t2x[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 773.880 1000.000 774.480 ;
    END
  END t2x[17]
  PIN t2x[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 784.760 1000.000 785.360 ;
    END
  END t2x[18]
  PIN t2x[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 795.640 1000.000 796.240 ;
    END
  END t2x[19]
  PIN t2x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 599.800 1000.000 600.400 ;
    END
  END t2x[1]
  PIN t2x[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 806.520 1000.000 807.120 ;
    END
  END t2x[20]
  PIN t2x[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 817.400 1000.000 818.000 ;
    END
  END t2x[21]
  PIN t2x[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 828.280 1000.000 828.880 ;
    END
  END t2x[22]
  PIN t2x[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 839.160 1000.000 839.760 ;
    END
  END t2x[23]
  PIN t2x[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 850.040 1000.000 850.640 ;
    END
  END t2x[24]
  PIN t2x[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 860.920 1000.000 861.520 ;
    END
  END t2x[25]
  PIN t2x[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 871.800 1000.000 872.400 ;
    END
  END t2x[26]
  PIN t2x[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 882.680 1000.000 883.280 ;
    END
  END t2x[27]
  PIN t2x[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 893.560 1000.000 894.160 ;
    END
  END t2x[28]
  PIN t2x[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 904.440 1000.000 905.040 ;
    END
  END t2x[29]
  PIN t2x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 610.680 1000.000 611.280 ;
    END
  END t2x[2]
  PIN t2x[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 915.320 1000.000 915.920 ;
    END
  END t2x[30]
  PIN t2x[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 926.200 1000.000 926.800 ;
    END
  END t2x[31]
  PIN t2x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 621.560 1000.000 622.160 ;
    END
  END t2x[3]
  PIN t2x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 632.440 1000.000 633.040 ;
    END
  END t2x[4]
  PIN t2x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 643.320 1000.000 643.920 ;
    END
  END t2x[5]
  PIN t2x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 654.200 1000.000 654.800 ;
    END
  END t2x[6]
  PIN t2x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 665.080 1000.000 665.680 ;
    END
  END t2x[7]
  PIN t2x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 675.960 1000.000 676.560 ;
    END
  END t2x[8]
  PIN t2x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 686.840 1000.000 687.440 ;
    END
  END t2x[9]
  PIN t2y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 594.360 1000.000 594.960 ;
    END
  END t2y[0]
  PIN t2y[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 703.160 1000.000 703.760 ;
    END
  END t2y[10]
  PIN t2y[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 714.040 1000.000 714.640 ;
    END
  END t2y[11]
  PIN t2y[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 724.920 1000.000 725.520 ;
    END
  END t2y[12]
  PIN t2y[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 735.800 1000.000 736.400 ;
    END
  END t2y[13]
  PIN t2y[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 746.680 1000.000 747.280 ;
    END
  END t2y[14]
  PIN t2y[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 757.560 1000.000 758.160 ;
    END
  END t2y[15]
  PIN t2y[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 768.440 1000.000 769.040 ;
    END
  END t2y[16]
  PIN t2y[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 779.320 1000.000 779.920 ;
    END
  END t2y[17]
  PIN t2y[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 790.200 1000.000 790.800 ;
    END
  END t2y[18]
  PIN t2y[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 801.080 1000.000 801.680 ;
    END
  END t2y[19]
  PIN t2y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 605.240 1000.000 605.840 ;
    END
  END t2y[1]
  PIN t2y[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 811.960 1000.000 812.560 ;
    END
  END t2y[20]
  PIN t2y[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 822.840 1000.000 823.440 ;
    END
  END t2y[21]
  PIN t2y[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 833.720 1000.000 834.320 ;
    END
  END t2y[22]
  PIN t2y[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 844.600 1000.000 845.200 ;
    END
  END t2y[23]
  PIN t2y[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 855.480 1000.000 856.080 ;
    END
  END t2y[24]
  PIN t2y[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 866.360 1000.000 866.960 ;
    END
  END t2y[25]
  PIN t2y[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 877.240 1000.000 877.840 ;
    END
  END t2y[26]
  PIN t2y[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 888.120 1000.000 888.720 ;
    END
  END t2y[27]
  PIN t2y[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 899.000 1000.000 899.600 ;
    END
  END t2y[28]
  PIN t2y[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 909.880 1000.000 910.480 ;
    END
  END t2y[29]
  PIN t2y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 616.120 1000.000 616.720 ;
    END
  END t2y[2]
  PIN t2y[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 920.760 1000.000 921.360 ;
    END
  END t2y[30]
  PIN t2y[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 931.640 1000.000 932.240 ;
    END
  END t2y[31]
  PIN t2y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 627.000 1000.000 627.600 ;
    END
  END t2y[3]
  PIN t2y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 637.880 1000.000 638.480 ;
    END
  END t2y[4]
  PIN t2y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 648.760 1000.000 649.360 ;
    END
  END t2y[5]
  PIN t2y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 659.640 1000.000 660.240 ;
    END
  END t2y[6]
  PIN t2y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 670.520 1000.000 671.120 ;
    END
  END t2y[7]
  PIN t2y[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 681.400 1000.000 682.000 ;
    END
  END t2y[8]
  PIN t2y[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 692.280 1000.000 692.880 ;
    END
  END t2y[9]
  PIN v0x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END v0x[0]
  PIN v0x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END v0x[10]
  PIN v0x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END v0x[11]
  PIN v0x[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END v0x[12]
  PIN v0x[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END v0x[13]
  PIN v0x[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END v0x[14]
  PIN v0x[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END v0x[15]
  PIN v0x[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 311.510 0.000 311.790 4.000 ;
    END
  END v0x[16]
  PIN v0x[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END v0x[17]
  PIN v0x[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END v0x[18]
  PIN v0x[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END v0x[19]
  PIN v0x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END v0x[1]
  PIN v0x[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END v0x[20]
  PIN v0x[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END v0x[21]
  PIN v0x[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END v0x[22]
  PIN v0x[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END v0x[23]
  PIN v0x[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 455.030 0.000 455.310 4.000 ;
    END
  END v0x[24]
  PIN v0x[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 4.000 ;
    END
  END v0x[25]
  PIN v0x[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END v0x[26]
  PIN v0x[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 508.850 0.000 509.130 4.000 ;
    END
  END v0x[27]
  PIN v0x[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 4.000 ;
    END
  END v0x[28]
  PIN v0x[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END v0x[29]
  PIN v0x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END v0x[2]
  PIN v0x[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END v0x[30]
  PIN v0x[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END v0x[31]
  PIN v0x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END v0x[3]
  PIN v0x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END v0x[4]
  PIN v0x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END v0x[5]
  PIN v0x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END v0x[6]
  PIN v0x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END v0x[7]
  PIN v0x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END v0x[8]
  PIN v0x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END v0x[9]
  PIN v0y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END v0y[0]
  PIN v0y[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END v0y[10]
  PIN v0y[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END v0y[11]
  PIN v0y[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 245.730 0.000 246.010 4.000 ;
    END
  END v0y[12]
  PIN v0y[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 263.670 0.000 263.950 4.000 ;
    END
  END v0y[13]
  PIN v0y[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END v0y[14]
  PIN v0y[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END v0y[15]
  PIN v0y[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END v0y[16]
  PIN v0y[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END v0y[17]
  PIN v0y[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END v0y[18]
  PIN v0y[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 371.310 0.000 371.590 4.000 ;
    END
  END v0y[19]
  PIN v0y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END v0y[1]
  PIN v0y[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 389.250 0.000 389.530 4.000 ;
    END
  END v0y[20]
  PIN v0y[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END v0y[21]
  PIN v0y[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END v0y[22]
  PIN v0y[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END v0y[23]
  PIN v0y[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END v0y[24]
  PIN v0y[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END v0y[25]
  PIN v0y[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 496.890 0.000 497.170 4.000 ;
    END
  END v0y[26]
  PIN v0y[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END v0y[27]
  PIN v0y[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 4.000 ;
    END
  END v0y[28]
  PIN v0y[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END v0y[29]
  PIN v0y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END v0y[2]
  PIN v0y[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 568.650 0.000 568.930 4.000 ;
    END
  END v0y[30]
  PIN v0y[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END v0y[31]
  PIN v0y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END v0y[3]
  PIN v0y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END v0y[4]
  PIN v0y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END v0y[5]
  PIN v0y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END v0y[6]
  PIN v0y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END v0y[7]
  PIN v0y[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END v0y[8]
  PIN v0y[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END v0y[9]
  PIN v0z[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END v0z[0]
  PIN v0z[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END v0z[10]
  PIN v0z[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END v0z[11]
  PIN v0z[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 4.000 ;
    END
  END v0z[12]
  PIN v0z[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END v0z[13]
  PIN v0z[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END v0z[14]
  PIN v0z[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END v0z[15]
  PIN v0z[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 0.000 323.750 4.000 ;
    END
  END v0z[16]
  PIN v0z[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END v0z[17]
  PIN v0z[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END v0z[18]
  PIN v0z[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 0.000 377.570 4.000 ;
    END
  END v0z[19]
  PIN v0z[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END v0z[1]
  PIN v0z[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 0.000 395.510 4.000 ;
    END
  END v0z[20]
  PIN v0z[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END v0z[21]
  PIN v0z[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 0.000 431.390 4.000 ;
    END
  END v0z[22]
  PIN v0z[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END v0z[23]
  PIN v0z[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END v0z[24]
  PIN v0z[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END v0z[25]
  PIN v0z[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 0.000 503.150 4.000 ;
    END
  END v0z[26]
  PIN v0z[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END v0z[27]
  PIN v0z[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 4.000 ;
    END
  END v0z[28]
  PIN v0z[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END v0z[29]
  PIN v0z[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END v0z[2]
  PIN v0z[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END v0z[30]
  PIN v0z[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 0.000 592.850 4.000 ;
    END
  END v0z[31]
  PIN v0z[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END v0z[3]
  PIN v0z[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END v0z[4]
  PIN v0z[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END v0z[5]
  PIN v0z[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END v0z[6]
  PIN v0z[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END v0z[7]
  PIN v0z[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END v0z[8]
  PIN v0z[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END v0z[9]
  PIN v1x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 24.470 996.000 24.750 1000.000 ;
    END
  END v1x[0]
  PIN v1x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 203.870 996.000 204.150 1000.000 ;
    END
  END v1x[10]
  PIN v1x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 221.810 996.000 222.090 1000.000 ;
    END
  END v1x[11]
  PIN v1x[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 239.750 996.000 240.030 1000.000 ;
    END
  END v1x[12]
  PIN v1x[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 257.690 996.000 257.970 1000.000 ;
    END
  END v1x[13]
  PIN v1x[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 275.630 996.000 275.910 1000.000 ;
    END
  END v1x[14]
  PIN v1x[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 293.570 996.000 293.850 1000.000 ;
    END
  END v1x[15]
  PIN v1x[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 311.510 996.000 311.790 1000.000 ;
    END
  END v1x[16]
  PIN v1x[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 329.450 996.000 329.730 1000.000 ;
    END
  END v1x[17]
  PIN v1x[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 347.390 996.000 347.670 1000.000 ;
    END
  END v1x[18]
  PIN v1x[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 365.330 996.000 365.610 1000.000 ;
    END
  END v1x[19]
  PIN v1x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 42.410 996.000 42.690 1000.000 ;
    END
  END v1x[1]
  PIN v1x[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 383.270 996.000 383.550 1000.000 ;
    END
  END v1x[20]
  PIN v1x[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 401.210 996.000 401.490 1000.000 ;
    END
  END v1x[21]
  PIN v1x[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 419.150 996.000 419.430 1000.000 ;
    END
  END v1x[22]
  PIN v1x[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 437.090 996.000 437.370 1000.000 ;
    END
  END v1x[23]
  PIN v1x[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 455.030 996.000 455.310 1000.000 ;
    END
  END v1x[24]
  PIN v1x[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 472.970 996.000 473.250 1000.000 ;
    END
  END v1x[25]
  PIN v1x[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 490.910 996.000 491.190 1000.000 ;
    END
  END v1x[26]
  PIN v1x[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 508.850 996.000 509.130 1000.000 ;
    END
  END v1x[27]
  PIN v1x[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 526.790 996.000 527.070 1000.000 ;
    END
  END v1x[28]
  PIN v1x[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 544.730 996.000 545.010 1000.000 ;
    END
  END v1x[29]
  PIN v1x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 60.350 996.000 60.630 1000.000 ;
    END
  END v1x[2]
  PIN v1x[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 562.670 996.000 562.950 1000.000 ;
    END
  END v1x[30]
  PIN v1x[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 580.610 996.000 580.890 1000.000 ;
    END
  END v1x[31]
  PIN v1x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 78.290 996.000 78.570 1000.000 ;
    END
  END v1x[3]
  PIN v1x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 96.230 996.000 96.510 1000.000 ;
    END
  END v1x[4]
  PIN v1x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 114.170 996.000 114.450 1000.000 ;
    END
  END v1x[5]
  PIN v1x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 132.110 996.000 132.390 1000.000 ;
    END
  END v1x[6]
  PIN v1x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 150.050 996.000 150.330 1000.000 ;
    END
  END v1x[7]
  PIN v1x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 167.990 996.000 168.270 1000.000 ;
    END
  END v1x[8]
  PIN v1x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 185.930 996.000 186.210 1000.000 ;
    END
  END v1x[9]
  PIN v1y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 30.450 996.000 30.730 1000.000 ;
    END
  END v1y[0]
  PIN v1y[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 209.850 996.000 210.130 1000.000 ;
    END
  END v1y[10]
  PIN v1y[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 227.790 996.000 228.070 1000.000 ;
    END
  END v1y[11]
  PIN v1y[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 245.730 996.000 246.010 1000.000 ;
    END
  END v1y[12]
  PIN v1y[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 263.670 996.000 263.950 1000.000 ;
    END
  END v1y[13]
  PIN v1y[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 281.610 996.000 281.890 1000.000 ;
    END
  END v1y[14]
  PIN v1y[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 299.550 996.000 299.830 1000.000 ;
    END
  END v1y[15]
  PIN v1y[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 317.490 996.000 317.770 1000.000 ;
    END
  END v1y[16]
  PIN v1y[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 335.430 996.000 335.710 1000.000 ;
    END
  END v1y[17]
  PIN v1y[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 353.370 996.000 353.650 1000.000 ;
    END
  END v1y[18]
  PIN v1y[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 371.310 996.000 371.590 1000.000 ;
    END
  END v1y[19]
  PIN v1y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 996.000 48.670 1000.000 ;
    END
  END v1y[1]
  PIN v1y[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 389.250 996.000 389.530 1000.000 ;
    END
  END v1y[20]
  PIN v1y[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 407.190 996.000 407.470 1000.000 ;
    END
  END v1y[21]
  PIN v1y[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 425.130 996.000 425.410 1000.000 ;
    END
  END v1y[22]
  PIN v1y[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 443.070 996.000 443.350 1000.000 ;
    END
  END v1y[23]
  PIN v1y[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 461.010 996.000 461.290 1000.000 ;
    END
  END v1y[24]
  PIN v1y[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 478.950 996.000 479.230 1000.000 ;
    END
  END v1y[25]
  PIN v1y[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 496.890 996.000 497.170 1000.000 ;
    END
  END v1y[26]
  PIN v1y[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 514.830 996.000 515.110 1000.000 ;
    END
  END v1y[27]
  PIN v1y[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met2 ;
        RECT 532.770 996.000 533.050 1000.000 ;
    END
  END v1y[28]
  PIN v1y[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 550.710 996.000 550.990 1000.000 ;
    END
  END v1y[29]
  PIN v1y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 66.330 996.000 66.610 1000.000 ;
    END
  END v1y[2]
  PIN v1y[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met2 ;
        RECT 568.650 996.000 568.930 1000.000 ;
    END
  END v1y[30]
  PIN v1y[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 586.590 996.000 586.870 1000.000 ;
    END
  END v1y[31]
  PIN v1y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    PORT
      LAYER met2 ;
        RECT 84.270 996.000 84.550 1000.000 ;
    END
  END v1y[3]
  PIN v1y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 102.210 996.000 102.490 1000.000 ;
    END
  END v1y[4]
  PIN v1y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 120.150 996.000 120.430 1000.000 ;
    END
  END v1y[5]
  PIN v1y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 138.090 996.000 138.370 1000.000 ;
    END
  END v1y[6]
  PIN v1y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 156.030 996.000 156.310 1000.000 ;
    END
  END v1y[7]
  PIN v1y[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 173.970 996.000 174.250 1000.000 ;
    END
  END v1y[8]
  PIN v1y[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met2 ;
        RECT 191.910 996.000 192.190 1000.000 ;
    END
  END v1y[9]
  PIN v1z[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 996.000 36.710 1000.000 ;
    END
  END v1z[0]
  PIN v1z[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 996.000 216.110 1000.000 ;
    END
  END v1z[10]
  PIN v1z[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 996.000 234.050 1000.000 ;
    END
  END v1z[11]
  PIN v1z[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 996.000 251.990 1000.000 ;
    END
  END v1z[12]
  PIN v1z[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 996.000 269.930 1000.000 ;
    END
  END v1z[13]
  PIN v1z[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 996.000 287.870 1000.000 ;
    END
  END v1z[14]
  PIN v1z[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 996.000 305.810 1000.000 ;
    END
  END v1z[15]
  PIN v1z[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 996.000 323.750 1000.000 ;
    END
  END v1z[16]
  PIN v1z[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 996.000 341.690 1000.000 ;
    END
  END v1z[17]
  PIN v1z[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 996.000 359.630 1000.000 ;
    END
  END v1z[18]
  PIN v1z[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 996.000 377.570 1000.000 ;
    END
  END v1z[19]
  PIN v1z[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 996.000 54.650 1000.000 ;
    END
  END v1z[1]
  PIN v1z[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.230 996.000 395.510 1000.000 ;
    END
  END v1z[20]
  PIN v1z[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 996.000 413.450 1000.000 ;
    END
  END v1z[21]
  PIN v1z[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.110 996.000 431.390 1000.000 ;
    END
  END v1z[22]
  PIN v1z[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 996.000 449.330 1000.000 ;
    END
  END v1z[23]
  PIN v1z[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 996.000 467.270 1000.000 ;
    END
  END v1z[24]
  PIN v1z[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.930 996.000 485.210 1000.000 ;
    END
  END v1z[25]
  PIN v1z[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 996.000 503.150 1000.000 ;
    END
  END v1z[26]
  PIN v1z[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 996.000 521.090 1000.000 ;
    END
  END v1z[27]
  PIN v1z[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.750 996.000 539.030 1000.000 ;
    END
  END v1z[28]
  PIN v1z[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 996.000 556.970 1000.000 ;
    END
  END v1z[29]
  PIN v1z[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 996.000 72.590 1000.000 ;
    END
  END v1z[2]
  PIN v1z[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 996.000 574.910 1000.000 ;
    END
  END v1z[30]
  PIN v1z[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.570 996.000 592.850 1000.000 ;
    END
  END v1z[31]
  PIN v1z[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 996.000 90.530 1000.000 ;
    END
  END v1z[3]
  PIN v1z[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 996.000 108.470 1000.000 ;
    END
  END v1z[4]
  PIN v1z[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 996.000 126.410 1000.000 ;
    END
  END v1z[5]
  PIN v1z[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 996.000 144.350 1000.000 ;
    END
  END v1z[6]
  PIN v1z[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 996.000 162.290 1000.000 ;
    END
  END v1z[7]
  PIN v1z[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 996.000 180.230 1000.000 ;
    END
  END v1z[8]
  PIN v1z[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 996.000 198.170 1000.000 ;
    END
  END v1z[9]
  PIN v2x[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 66.680 1000.000 67.280 ;
    END
  END v2x[0]
  PIN v2x[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 229.880 1000.000 230.480 ;
    END
  END v2x[10]
  PIN v2x[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 246.200 1000.000 246.800 ;
    END
  END v2x[11]
  PIN v2x[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 262.520 1000.000 263.120 ;
    END
  END v2x[12]
  PIN v2x[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 278.840 1000.000 279.440 ;
    END
  END v2x[13]
  PIN v2x[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 295.160 1000.000 295.760 ;
    END
  END v2x[14]
  PIN v2x[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 311.480 1000.000 312.080 ;
    END
  END v2x[15]
  PIN v2x[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 327.800 1000.000 328.400 ;
    END
  END v2x[16]
  PIN v2x[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 344.120 1000.000 344.720 ;
    END
  END v2x[17]
  PIN v2x[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 360.440 1000.000 361.040 ;
    END
  END v2x[18]
  PIN v2x[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 376.760 1000.000 377.360 ;
    END
  END v2x[19]
  PIN v2x[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 83.000 1000.000 83.600 ;
    END
  END v2x[1]
  PIN v2x[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 393.080 1000.000 393.680 ;
    END
  END v2x[20]
  PIN v2x[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 409.400 1000.000 410.000 ;
    END
  END v2x[21]
  PIN v2x[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 425.720 1000.000 426.320 ;
    END
  END v2x[22]
  PIN v2x[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 442.040 1000.000 442.640 ;
    END
  END v2x[23]
  PIN v2x[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 458.360 1000.000 458.960 ;
    END
  END v2x[24]
  PIN v2x[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 474.680 1000.000 475.280 ;
    END
  END v2x[25]
  PIN v2x[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 491.000 1000.000 491.600 ;
    END
  END v2x[26]
  PIN v2x[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 507.320 1000.000 507.920 ;
    END
  END v2x[27]
  PIN v2x[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 523.640 1000.000 524.240 ;
    END
  END v2x[28]
  PIN v2x[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 539.960 1000.000 540.560 ;
    END
  END v2x[29]
  PIN v2x[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 99.320 1000.000 99.920 ;
    END
  END v2x[2]
  PIN v2x[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 556.280 1000.000 556.880 ;
    END
  END v2x[30]
  PIN v2x[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 572.600 1000.000 573.200 ;
    END
  END v2x[31]
  PIN v2x[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 115.640 1000.000 116.240 ;
    END
  END v2x[3]
  PIN v2x[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 131.960 1000.000 132.560 ;
    END
  END v2x[4]
  PIN v2x[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 148.280 1000.000 148.880 ;
    END
  END v2x[5]
  PIN v2x[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 164.600 1000.000 165.200 ;
    END
  END v2x[6]
  PIN v2x[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 180.920 1000.000 181.520 ;
    END
  END v2x[7]
  PIN v2x[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 197.240 1000.000 197.840 ;
    END
  END v2x[8]
  PIN v2x[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 213.560 1000.000 214.160 ;
    END
  END v2x[9]
  PIN v2y[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 72.120 1000.000 72.720 ;
    END
  END v2y[0]
  PIN v2y[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 235.320 1000.000 235.920 ;
    END
  END v2y[10]
  PIN v2y[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 251.640 1000.000 252.240 ;
    END
  END v2y[11]
  PIN v2y[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 267.960 1000.000 268.560 ;
    END
  END v2y[12]
  PIN v2y[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 284.280 1000.000 284.880 ;
    END
  END v2y[13]
  PIN v2y[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 300.600 1000.000 301.200 ;
    END
  END v2y[14]
  PIN v2y[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 316.920 1000.000 317.520 ;
    END
  END v2y[15]
  PIN v2y[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 333.240 1000.000 333.840 ;
    END
  END v2y[16]
  PIN v2y[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 349.560 1000.000 350.160 ;
    END
  END v2y[17]
  PIN v2y[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 365.880 1000.000 366.480 ;
    END
  END v2y[18]
  PIN v2y[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 382.200 1000.000 382.800 ;
    END
  END v2y[19]
  PIN v2y[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 88.440 1000.000 89.040 ;
    END
  END v2y[1]
  PIN v2y[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 398.520 1000.000 399.120 ;
    END
  END v2y[20]
  PIN v2y[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 414.840 1000.000 415.440 ;
    END
  END v2y[21]
  PIN v2y[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 431.160 1000.000 431.760 ;
    END
  END v2y[22]
  PIN v2y[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 447.480 1000.000 448.080 ;
    END
  END v2y[23]
  PIN v2y[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 463.800 1000.000 464.400 ;
    END
  END v2y[24]
  PIN v2y[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 480.120 1000.000 480.720 ;
    END
  END v2y[25]
  PIN v2y[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 496.440 1000.000 497.040 ;
    END
  END v2y[26]
  PIN v2y[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 512.760 1000.000 513.360 ;
    END
  END v2y[27]
  PIN v2y[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 529.080 1000.000 529.680 ;
    END
  END v2y[28]
  PIN v2y[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 545.400 1000.000 546.000 ;
    END
  END v2y[29]
  PIN v2y[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 104.760 1000.000 105.360 ;
    END
  END v2y[2]
  PIN v2y[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 561.720 1000.000 562.320 ;
    END
  END v2y[30]
  PIN v2y[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 578.040 1000.000 578.640 ;
    END
  END v2y[31]
  PIN v2y[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 121.080 1000.000 121.680 ;
    END
  END v2y[3]
  PIN v2y[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 137.400 1000.000 138.000 ;
    END
  END v2y[4]
  PIN v2y[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 153.720 1000.000 154.320 ;
    END
  END v2y[5]
  PIN v2y[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 170.040 1000.000 170.640 ;
    END
  END v2y[6]
  PIN v2y[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 186.360 1000.000 186.960 ;
    END
  END v2y[7]
  PIN v2y[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.742500 ;
    PORT
      LAYER met3 ;
        RECT 996.000 202.680 1000.000 203.280 ;
    END
  END v2y[8]
  PIN v2y[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.495000 ;
    PORT
      LAYER met3 ;
        RECT 996.000 219.000 1000.000 219.600 ;
    END
  END v2y[9]
  PIN v2z[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 77.560 1000.000 78.160 ;
    END
  END v2z[0]
  PIN v2z[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 240.760 1000.000 241.360 ;
    END
  END v2z[10]
  PIN v2z[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 257.080 1000.000 257.680 ;
    END
  END v2z[11]
  PIN v2z[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 273.400 1000.000 274.000 ;
    END
  END v2z[12]
  PIN v2z[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 289.720 1000.000 290.320 ;
    END
  END v2z[13]
  PIN v2z[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 306.040 1000.000 306.640 ;
    END
  END v2z[14]
  PIN v2z[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 322.360 1000.000 322.960 ;
    END
  END v2z[15]
  PIN v2z[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 338.680 1000.000 339.280 ;
    END
  END v2z[16]
  PIN v2z[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 355.000 1000.000 355.600 ;
    END
  END v2z[17]
  PIN v2z[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 371.320 1000.000 371.920 ;
    END
  END v2z[18]
  PIN v2z[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 387.640 1000.000 388.240 ;
    END
  END v2z[19]
  PIN v2z[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 93.880 1000.000 94.480 ;
    END
  END v2z[1]
  PIN v2z[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 403.960 1000.000 404.560 ;
    END
  END v2z[20]
  PIN v2z[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 420.280 1000.000 420.880 ;
    END
  END v2z[21]
  PIN v2z[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 436.600 1000.000 437.200 ;
    END
  END v2z[22]
  PIN v2z[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 452.920 1000.000 453.520 ;
    END
  END v2z[23]
  PIN v2z[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 469.240 1000.000 469.840 ;
    END
  END v2z[24]
  PIN v2z[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 485.560 1000.000 486.160 ;
    END
  END v2z[25]
  PIN v2z[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 501.880 1000.000 502.480 ;
    END
  END v2z[26]
  PIN v2z[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 518.200 1000.000 518.800 ;
    END
  END v2z[27]
  PIN v2z[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 534.520 1000.000 535.120 ;
    END
  END v2z[28]
  PIN v2z[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 550.840 1000.000 551.440 ;
    END
  END v2z[29]
  PIN v2z[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 110.200 1000.000 110.800 ;
    END
  END v2z[2]
  PIN v2z[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 567.160 1000.000 567.760 ;
    END
  END v2z[30]
  PIN v2z[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 583.480 1000.000 584.080 ;
    END
  END v2z[31]
  PIN v2z[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 126.520 1000.000 127.120 ;
    END
  END v2z[3]
  PIN v2z[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 142.840 1000.000 143.440 ;
    END
  END v2z[4]
  PIN v2z[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 159.160 1000.000 159.760 ;
    END
  END v2z[5]
  PIN v2z[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 175.480 1000.000 176.080 ;
    END
  END v2z[6]
  PIN v2z[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 191.800 1000.000 192.400 ;
    END
  END v2z[7]
  PIN v2z[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 208.120 1000.000 208.720 ;
    END
  END v2z[8]
  PIN v2z[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 996.000 224.440 1000.000 225.040 ;
    END
  END v2z[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 987.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 987.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 987.600 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 994.060 987.445 ;
      LAYER met1 ;
        RECT 4.670 6.160 994.910 987.600 ;
      LAYER met2 ;
        RECT 4.690 995.720 24.190 996.610 ;
        RECT 25.030 995.720 30.170 996.610 ;
        RECT 31.010 995.720 36.150 996.610 ;
        RECT 36.990 995.720 42.130 996.610 ;
        RECT 42.970 995.720 48.110 996.610 ;
        RECT 48.950 995.720 54.090 996.610 ;
        RECT 54.930 995.720 60.070 996.610 ;
        RECT 60.910 995.720 66.050 996.610 ;
        RECT 66.890 995.720 72.030 996.610 ;
        RECT 72.870 995.720 78.010 996.610 ;
        RECT 78.850 995.720 83.990 996.610 ;
        RECT 84.830 995.720 89.970 996.610 ;
        RECT 90.810 995.720 95.950 996.610 ;
        RECT 96.790 995.720 101.930 996.610 ;
        RECT 102.770 995.720 107.910 996.610 ;
        RECT 108.750 995.720 113.890 996.610 ;
        RECT 114.730 995.720 119.870 996.610 ;
        RECT 120.710 995.720 125.850 996.610 ;
        RECT 126.690 995.720 131.830 996.610 ;
        RECT 132.670 995.720 137.810 996.610 ;
        RECT 138.650 995.720 143.790 996.610 ;
        RECT 144.630 995.720 149.770 996.610 ;
        RECT 150.610 995.720 155.750 996.610 ;
        RECT 156.590 995.720 161.730 996.610 ;
        RECT 162.570 995.720 167.710 996.610 ;
        RECT 168.550 995.720 173.690 996.610 ;
        RECT 174.530 995.720 179.670 996.610 ;
        RECT 180.510 995.720 185.650 996.610 ;
        RECT 186.490 995.720 191.630 996.610 ;
        RECT 192.470 995.720 197.610 996.610 ;
        RECT 198.450 995.720 203.590 996.610 ;
        RECT 204.430 995.720 209.570 996.610 ;
        RECT 210.410 995.720 215.550 996.610 ;
        RECT 216.390 995.720 221.530 996.610 ;
        RECT 222.370 995.720 227.510 996.610 ;
        RECT 228.350 995.720 233.490 996.610 ;
        RECT 234.330 995.720 239.470 996.610 ;
        RECT 240.310 995.720 245.450 996.610 ;
        RECT 246.290 995.720 251.430 996.610 ;
        RECT 252.270 995.720 257.410 996.610 ;
        RECT 258.250 995.720 263.390 996.610 ;
        RECT 264.230 995.720 269.370 996.610 ;
        RECT 270.210 995.720 275.350 996.610 ;
        RECT 276.190 995.720 281.330 996.610 ;
        RECT 282.170 995.720 287.310 996.610 ;
        RECT 288.150 995.720 293.290 996.610 ;
        RECT 294.130 995.720 299.270 996.610 ;
        RECT 300.110 995.720 305.250 996.610 ;
        RECT 306.090 995.720 311.230 996.610 ;
        RECT 312.070 995.720 317.210 996.610 ;
        RECT 318.050 995.720 323.190 996.610 ;
        RECT 324.030 995.720 329.170 996.610 ;
        RECT 330.010 995.720 335.150 996.610 ;
        RECT 335.990 995.720 341.130 996.610 ;
        RECT 341.970 995.720 347.110 996.610 ;
        RECT 347.950 995.720 353.090 996.610 ;
        RECT 353.930 995.720 359.070 996.610 ;
        RECT 359.910 995.720 365.050 996.610 ;
        RECT 365.890 995.720 371.030 996.610 ;
        RECT 371.870 995.720 377.010 996.610 ;
        RECT 377.850 995.720 382.990 996.610 ;
        RECT 383.830 995.720 388.970 996.610 ;
        RECT 389.810 995.720 394.950 996.610 ;
        RECT 395.790 995.720 400.930 996.610 ;
        RECT 401.770 995.720 406.910 996.610 ;
        RECT 407.750 995.720 412.890 996.610 ;
        RECT 413.730 995.720 418.870 996.610 ;
        RECT 419.710 995.720 424.850 996.610 ;
        RECT 425.690 995.720 430.830 996.610 ;
        RECT 431.670 995.720 436.810 996.610 ;
        RECT 437.650 995.720 442.790 996.610 ;
        RECT 443.630 995.720 448.770 996.610 ;
        RECT 449.610 995.720 454.750 996.610 ;
        RECT 455.590 995.720 460.730 996.610 ;
        RECT 461.570 995.720 466.710 996.610 ;
        RECT 467.550 995.720 472.690 996.610 ;
        RECT 473.530 995.720 478.670 996.610 ;
        RECT 479.510 995.720 484.650 996.610 ;
        RECT 485.490 995.720 490.630 996.610 ;
        RECT 491.470 995.720 496.610 996.610 ;
        RECT 497.450 995.720 502.590 996.610 ;
        RECT 503.430 995.720 508.570 996.610 ;
        RECT 509.410 995.720 514.550 996.610 ;
        RECT 515.390 995.720 520.530 996.610 ;
        RECT 521.370 995.720 526.510 996.610 ;
        RECT 527.350 995.720 532.490 996.610 ;
        RECT 533.330 995.720 538.470 996.610 ;
        RECT 539.310 995.720 544.450 996.610 ;
        RECT 545.290 995.720 550.430 996.610 ;
        RECT 551.270 995.720 556.410 996.610 ;
        RECT 557.250 995.720 562.390 996.610 ;
        RECT 563.230 995.720 568.370 996.610 ;
        RECT 569.210 995.720 574.350 996.610 ;
        RECT 575.190 995.720 580.330 996.610 ;
        RECT 581.170 995.720 586.310 996.610 ;
        RECT 587.150 995.720 592.290 996.610 ;
        RECT 593.130 995.720 598.270 996.610 ;
        RECT 599.110 995.720 604.250 996.610 ;
        RECT 605.090 995.720 610.230 996.610 ;
        RECT 611.070 995.720 616.210 996.610 ;
        RECT 617.050 995.720 622.190 996.610 ;
        RECT 623.030 995.720 628.170 996.610 ;
        RECT 629.010 995.720 634.150 996.610 ;
        RECT 634.990 995.720 640.130 996.610 ;
        RECT 640.970 995.720 646.110 996.610 ;
        RECT 646.950 995.720 652.090 996.610 ;
        RECT 652.930 995.720 658.070 996.610 ;
        RECT 658.910 995.720 664.050 996.610 ;
        RECT 664.890 995.720 670.030 996.610 ;
        RECT 670.870 995.720 676.010 996.610 ;
        RECT 676.850 995.720 681.990 996.610 ;
        RECT 682.830 995.720 687.970 996.610 ;
        RECT 688.810 995.720 693.950 996.610 ;
        RECT 694.790 995.720 699.930 996.610 ;
        RECT 700.770 995.720 705.910 996.610 ;
        RECT 706.750 995.720 711.890 996.610 ;
        RECT 712.730 995.720 717.870 996.610 ;
        RECT 718.710 995.720 723.850 996.610 ;
        RECT 724.690 995.720 729.830 996.610 ;
        RECT 730.670 995.720 735.810 996.610 ;
        RECT 736.650 995.720 741.790 996.610 ;
        RECT 742.630 995.720 747.770 996.610 ;
        RECT 748.610 995.720 753.750 996.610 ;
        RECT 754.590 995.720 759.730 996.610 ;
        RECT 760.570 995.720 765.710 996.610 ;
        RECT 766.550 995.720 771.690 996.610 ;
        RECT 772.530 995.720 777.670 996.610 ;
        RECT 778.510 995.720 783.650 996.610 ;
        RECT 784.490 995.720 789.630 996.610 ;
        RECT 790.470 995.720 795.610 996.610 ;
        RECT 796.450 995.720 801.590 996.610 ;
        RECT 802.430 995.720 807.570 996.610 ;
        RECT 808.410 995.720 813.550 996.610 ;
        RECT 814.390 995.720 819.530 996.610 ;
        RECT 820.370 995.720 825.510 996.610 ;
        RECT 826.350 995.720 831.490 996.610 ;
        RECT 832.330 995.720 837.470 996.610 ;
        RECT 838.310 995.720 843.450 996.610 ;
        RECT 844.290 995.720 849.430 996.610 ;
        RECT 850.270 995.720 855.410 996.610 ;
        RECT 856.250 995.720 861.390 996.610 ;
        RECT 862.230 995.720 867.370 996.610 ;
        RECT 868.210 995.720 873.350 996.610 ;
        RECT 874.190 995.720 879.330 996.610 ;
        RECT 880.170 995.720 885.310 996.610 ;
        RECT 886.150 995.720 891.290 996.610 ;
        RECT 892.130 995.720 897.270 996.610 ;
        RECT 898.110 995.720 903.250 996.610 ;
        RECT 904.090 995.720 909.230 996.610 ;
        RECT 910.070 995.720 915.210 996.610 ;
        RECT 916.050 995.720 921.190 996.610 ;
        RECT 922.030 995.720 927.170 996.610 ;
        RECT 928.010 995.720 933.150 996.610 ;
        RECT 933.990 995.720 939.130 996.610 ;
        RECT 939.970 995.720 945.110 996.610 ;
        RECT 945.950 995.720 951.090 996.610 ;
        RECT 951.930 995.720 957.070 996.610 ;
        RECT 957.910 995.720 963.050 996.610 ;
        RECT 963.890 995.720 969.030 996.610 ;
        RECT 969.870 995.720 975.010 996.610 ;
        RECT 975.850 995.720 994.890 996.610 ;
        RECT 4.690 4.280 994.890 995.720 ;
        RECT 4.690 3.670 24.190 4.280 ;
        RECT 25.030 3.670 30.170 4.280 ;
        RECT 31.010 3.670 36.150 4.280 ;
        RECT 36.990 3.670 42.130 4.280 ;
        RECT 42.970 3.670 48.110 4.280 ;
        RECT 48.950 3.670 54.090 4.280 ;
        RECT 54.930 3.670 60.070 4.280 ;
        RECT 60.910 3.670 66.050 4.280 ;
        RECT 66.890 3.670 72.030 4.280 ;
        RECT 72.870 3.670 78.010 4.280 ;
        RECT 78.850 3.670 83.990 4.280 ;
        RECT 84.830 3.670 89.970 4.280 ;
        RECT 90.810 3.670 95.950 4.280 ;
        RECT 96.790 3.670 101.930 4.280 ;
        RECT 102.770 3.670 107.910 4.280 ;
        RECT 108.750 3.670 113.890 4.280 ;
        RECT 114.730 3.670 119.870 4.280 ;
        RECT 120.710 3.670 125.850 4.280 ;
        RECT 126.690 3.670 131.830 4.280 ;
        RECT 132.670 3.670 137.810 4.280 ;
        RECT 138.650 3.670 143.790 4.280 ;
        RECT 144.630 3.670 149.770 4.280 ;
        RECT 150.610 3.670 155.750 4.280 ;
        RECT 156.590 3.670 161.730 4.280 ;
        RECT 162.570 3.670 167.710 4.280 ;
        RECT 168.550 3.670 173.690 4.280 ;
        RECT 174.530 3.670 179.670 4.280 ;
        RECT 180.510 3.670 185.650 4.280 ;
        RECT 186.490 3.670 191.630 4.280 ;
        RECT 192.470 3.670 197.610 4.280 ;
        RECT 198.450 3.670 203.590 4.280 ;
        RECT 204.430 3.670 209.570 4.280 ;
        RECT 210.410 3.670 215.550 4.280 ;
        RECT 216.390 3.670 221.530 4.280 ;
        RECT 222.370 3.670 227.510 4.280 ;
        RECT 228.350 3.670 233.490 4.280 ;
        RECT 234.330 3.670 239.470 4.280 ;
        RECT 240.310 3.670 245.450 4.280 ;
        RECT 246.290 3.670 251.430 4.280 ;
        RECT 252.270 3.670 257.410 4.280 ;
        RECT 258.250 3.670 263.390 4.280 ;
        RECT 264.230 3.670 269.370 4.280 ;
        RECT 270.210 3.670 275.350 4.280 ;
        RECT 276.190 3.670 281.330 4.280 ;
        RECT 282.170 3.670 287.310 4.280 ;
        RECT 288.150 3.670 293.290 4.280 ;
        RECT 294.130 3.670 299.270 4.280 ;
        RECT 300.110 3.670 305.250 4.280 ;
        RECT 306.090 3.670 311.230 4.280 ;
        RECT 312.070 3.670 317.210 4.280 ;
        RECT 318.050 3.670 323.190 4.280 ;
        RECT 324.030 3.670 329.170 4.280 ;
        RECT 330.010 3.670 335.150 4.280 ;
        RECT 335.990 3.670 341.130 4.280 ;
        RECT 341.970 3.670 347.110 4.280 ;
        RECT 347.950 3.670 353.090 4.280 ;
        RECT 353.930 3.670 359.070 4.280 ;
        RECT 359.910 3.670 365.050 4.280 ;
        RECT 365.890 3.670 371.030 4.280 ;
        RECT 371.870 3.670 377.010 4.280 ;
        RECT 377.850 3.670 382.990 4.280 ;
        RECT 383.830 3.670 388.970 4.280 ;
        RECT 389.810 3.670 394.950 4.280 ;
        RECT 395.790 3.670 400.930 4.280 ;
        RECT 401.770 3.670 406.910 4.280 ;
        RECT 407.750 3.670 412.890 4.280 ;
        RECT 413.730 3.670 418.870 4.280 ;
        RECT 419.710 3.670 424.850 4.280 ;
        RECT 425.690 3.670 430.830 4.280 ;
        RECT 431.670 3.670 436.810 4.280 ;
        RECT 437.650 3.670 442.790 4.280 ;
        RECT 443.630 3.670 448.770 4.280 ;
        RECT 449.610 3.670 454.750 4.280 ;
        RECT 455.590 3.670 460.730 4.280 ;
        RECT 461.570 3.670 466.710 4.280 ;
        RECT 467.550 3.670 472.690 4.280 ;
        RECT 473.530 3.670 478.670 4.280 ;
        RECT 479.510 3.670 484.650 4.280 ;
        RECT 485.490 3.670 490.630 4.280 ;
        RECT 491.470 3.670 496.610 4.280 ;
        RECT 497.450 3.670 502.590 4.280 ;
        RECT 503.430 3.670 508.570 4.280 ;
        RECT 509.410 3.670 514.550 4.280 ;
        RECT 515.390 3.670 520.530 4.280 ;
        RECT 521.370 3.670 526.510 4.280 ;
        RECT 527.350 3.670 532.490 4.280 ;
        RECT 533.330 3.670 538.470 4.280 ;
        RECT 539.310 3.670 544.450 4.280 ;
        RECT 545.290 3.670 550.430 4.280 ;
        RECT 551.270 3.670 556.410 4.280 ;
        RECT 557.250 3.670 562.390 4.280 ;
        RECT 563.230 3.670 568.370 4.280 ;
        RECT 569.210 3.670 574.350 4.280 ;
        RECT 575.190 3.670 580.330 4.280 ;
        RECT 581.170 3.670 586.310 4.280 ;
        RECT 587.150 3.670 592.290 4.280 ;
        RECT 593.130 3.670 598.270 4.280 ;
        RECT 599.110 3.670 604.250 4.280 ;
        RECT 605.090 3.670 610.230 4.280 ;
        RECT 611.070 3.670 616.210 4.280 ;
        RECT 617.050 3.670 622.190 4.280 ;
        RECT 623.030 3.670 628.170 4.280 ;
        RECT 629.010 3.670 634.150 4.280 ;
        RECT 634.990 3.670 640.130 4.280 ;
        RECT 640.970 3.670 646.110 4.280 ;
        RECT 646.950 3.670 652.090 4.280 ;
        RECT 652.930 3.670 658.070 4.280 ;
        RECT 658.910 3.670 664.050 4.280 ;
        RECT 664.890 3.670 670.030 4.280 ;
        RECT 670.870 3.670 676.010 4.280 ;
        RECT 676.850 3.670 681.990 4.280 ;
        RECT 682.830 3.670 687.970 4.280 ;
        RECT 688.810 3.670 693.950 4.280 ;
        RECT 694.790 3.670 699.930 4.280 ;
        RECT 700.770 3.670 705.910 4.280 ;
        RECT 706.750 3.670 711.890 4.280 ;
        RECT 712.730 3.670 717.870 4.280 ;
        RECT 718.710 3.670 723.850 4.280 ;
        RECT 724.690 3.670 729.830 4.280 ;
        RECT 730.670 3.670 735.810 4.280 ;
        RECT 736.650 3.670 741.790 4.280 ;
        RECT 742.630 3.670 747.770 4.280 ;
        RECT 748.610 3.670 753.750 4.280 ;
        RECT 754.590 3.670 759.730 4.280 ;
        RECT 760.570 3.670 765.710 4.280 ;
        RECT 766.550 3.670 771.690 4.280 ;
        RECT 772.530 3.670 777.670 4.280 ;
        RECT 778.510 3.670 783.650 4.280 ;
        RECT 784.490 3.670 789.630 4.280 ;
        RECT 790.470 3.670 795.610 4.280 ;
        RECT 796.450 3.670 801.590 4.280 ;
        RECT 802.430 3.670 807.570 4.280 ;
        RECT 808.410 3.670 813.550 4.280 ;
        RECT 814.390 3.670 819.530 4.280 ;
        RECT 820.370 3.670 825.510 4.280 ;
        RECT 826.350 3.670 831.490 4.280 ;
        RECT 832.330 3.670 837.470 4.280 ;
        RECT 838.310 3.670 843.450 4.280 ;
        RECT 844.290 3.670 849.430 4.280 ;
        RECT 850.270 3.670 855.410 4.280 ;
        RECT 856.250 3.670 861.390 4.280 ;
        RECT 862.230 3.670 867.370 4.280 ;
        RECT 868.210 3.670 873.350 4.280 ;
        RECT 874.190 3.670 879.330 4.280 ;
        RECT 880.170 3.670 885.310 4.280 ;
        RECT 886.150 3.670 891.290 4.280 ;
        RECT 892.130 3.670 897.270 4.280 ;
        RECT 898.110 3.670 903.250 4.280 ;
        RECT 904.090 3.670 909.230 4.280 ;
        RECT 910.070 3.670 915.210 4.280 ;
        RECT 916.050 3.670 921.190 4.280 ;
        RECT 922.030 3.670 927.170 4.280 ;
        RECT 928.010 3.670 933.150 4.280 ;
        RECT 933.990 3.670 939.130 4.280 ;
        RECT 939.970 3.670 945.110 4.280 ;
        RECT 945.950 3.670 951.090 4.280 ;
        RECT 951.930 3.670 957.070 4.280 ;
        RECT 957.910 3.670 963.050 4.280 ;
        RECT 963.890 3.670 969.030 4.280 ;
        RECT 969.870 3.670 975.010 4.280 ;
        RECT 975.850 3.670 994.890 4.280 ;
      LAYER met3 ;
        RECT 3.990 951.680 996.000 987.525 ;
        RECT 4.400 950.280 996.000 951.680 ;
        RECT 3.990 942.160 996.000 950.280 ;
        RECT 4.400 940.760 996.000 942.160 ;
        RECT 3.990 932.640 996.000 940.760 ;
        RECT 4.400 931.240 995.600 932.640 ;
        RECT 3.990 927.200 996.000 931.240 ;
        RECT 3.990 925.800 995.600 927.200 ;
        RECT 3.990 923.120 996.000 925.800 ;
        RECT 4.400 921.760 996.000 923.120 ;
        RECT 4.400 921.720 995.600 921.760 ;
        RECT 3.990 920.360 995.600 921.720 ;
        RECT 3.990 916.320 996.000 920.360 ;
        RECT 3.990 914.920 995.600 916.320 ;
        RECT 3.990 913.600 996.000 914.920 ;
        RECT 4.400 912.200 996.000 913.600 ;
        RECT 3.990 910.880 996.000 912.200 ;
        RECT 3.990 909.480 995.600 910.880 ;
        RECT 3.990 905.440 996.000 909.480 ;
        RECT 3.990 904.080 995.600 905.440 ;
        RECT 4.400 904.040 995.600 904.080 ;
        RECT 4.400 902.680 996.000 904.040 ;
        RECT 3.990 900.000 996.000 902.680 ;
        RECT 3.990 898.600 995.600 900.000 ;
        RECT 3.990 894.560 996.000 898.600 ;
        RECT 4.400 893.160 995.600 894.560 ;
        RECT 3.990 889.120 996.000 893.160 ;
        RECT 3.990 887.720 995.600 889.120 ;
        RECT 3.990 885.040 996.000 887.720 ;
        RECT 4.400 883.680 996.000 885.040 ;
        RECT 4.400 883.640 995.600 883.680 ;
        RECT 3.990 882.280 995.600 883.640 ;
        RECT 3.990 878.240 996.000 882.280 ;
        RECT 3.990 876.840 995.600 878.240 ;
        RECT 3.990 875.520 996.000 876.840 ;
        RECT 4.400 874.120 996.000 875.520 ;
        RECT 3.990 872.800 996.000 874.120 ;
        RECT 3.990 871.400 995.600 872.800 ;
        RECT 3.990 867.360 996.000 871.400 ;
        RECT 3.990 866.000 995.600 867.360 ;
        RECT 4.400 865.960 995.600 866.000 ;
        RECT 4.400 864.600 996.000 865.960 ;
        RECT 3.990 861.920 996.000 864.600 ;
        RECT 3.990 860.520 995.600 861.920 ;
        RECT 3.990 856.480 996.000 860.520 ;
        RECT 4.400 855.080 995.600 856.480 ;
        RECT 3.990 851.040 996.000 855.080 ;
        RECT 3.990 849.640 995.600 851.040 ;
        RECT 3.990 846.960 996.000 849.640 ;
        RECT 4.400 845.600 996.000 846.960 ;
        RECT 4.400 845.560 995.600 845.600 ;
        RECT 3.990 844.200 995.600 845.560 ;
        RECT 3.990 840.160 996.000 844.200 ;
        RECT 3.990 838.760 995.600 840.160 ;
        RECT 3.990 837.440 996.000 838.760 ;
        RECT 4.400 836.040 996.000 837.440 ;
        RECT 3.990 834.720 996.000 836.040 ;
        RECT 3.990 833.320 995.600 834.720 ;
        RECT 3.990 829.280 996.000 833.320 ;
        RECT 3.990 827.920 995.600 829.280 ;
        RECT 4.400 827.880 995.600 827.920 ;
        RECT 4.400 826.520 996.000 827.880 ;
        RECT 3.990 823.840 996.000 826.520 ;
        RECT 3.990 822.440 995.600 823.840 ;
        RECT 3.990 818.400 996.000 822.440 ;
        RECT 4.400 817.000 995.600 818.400 ;
        RECT 3.990 812.960 996.000 817.000 ;
        RECT 3.990 811.560 995.600 812.960 ;
        RECT 3.990 808.880 996.000 811.560 ;
        RECT 4.400 807.520 996.000 808.880 ;
        RECT 4.400 807.480 995.600 807.520 ;
        RECT 3.990 806.120 995.600 807.480 ;
        RECT 3.990 802.080 996.000 806.120 ;
        RECT 3.990 800.680 995.600 802.080 ;
        RECT 3.990 799.360 996.000 800.680 ;
        RECT 4.400 797.960 996.000 799.360 ;
        RECT 3.990 796.640 996.000 797.960 ;
        RECT 3.990 795.240 995.600 796.640 ;
        RECT 3.990 791.200 996.000 795.240 ;
        RECT 3.990 789.840 995.600 791.200 ;
        RECT 4.400 789.800 995.600 789.840 ;
        RECT 4.400 788.440 996.000 789.800 ;
        RECT 3.990 785.760 996.000 788.440 ;
        RECT 3.990 784.360 995.600 785.760 ;
        RECT 3.990 780.320 996.000 784.360 ;
        RECT 4.400 778.920 995.600 780.320 ;
        RECT 3.990 774.880 996.000 778.920 ;
        RECT 3.990 773.480 995.600 774.880 ;
        RECT 3.990 770.800 996.000 773.480 ;
        RECT 4.400 769.440 996.000 770.800 ;
        RECT 4.400 769.400 995.600 769.440 ;
        RECT 3.990 768.040 995.600 769.400 ;
        RECT 3.990 764.000 996.000 768.040 ;
        RECT 3.990 762.600 995.600 764.000 ;
        RECT 3.990 761.280 996.000 762.600 ;
        RECT 4.400 759.880 996.000 761.280 ;
        RECT 3.990 758.560 996.000 759.880 ;
        RECT 3.990 757.160 995.600 758.560 ;
        RECT 3.990 753.120 996.000 757.160 ;
        RECT 3.990 751.760 995.600 753.120 ;
        RECT 4.400 751.720 995.600 751.760 ;
        RECT 4.400 750.360 996.000 751.720 ;
        RECT 3.990 747.680 996.000 750.360 ;
        RECT 3.990 746.280 995.600 747.680 ;
        RECT 3.990 742.240 996.000 746.280 ;
        RECT 4.400 740.840 995.600 742.240 ;
        RECT 3.990 736.800 996.000 740.840 ;
        RECT 3.990 735.400 995.600 736.800 ;
        RECT 3.990 732.720 996.000 735.400 ;
        RECT 4.400 731.360 996.000 732.720 ;
        RECT 4.400 731.320 995.600 731.360 ;
        RECT 3.990 729.960 995.600 731.320 ;
        RECT 3.990 725.920 996.000 729.960 ;
        RECT 3.990 724.520 995.600 725.920 ;
        RECT 3.990 723.200 996.000 724.520 ;
        RECT 4.400 721.800 996.000 723.200 ;
        RECT 3.990 720.480 996.000 721.800 ;
        RECT 3.990 719.080 995.600 720.480 ;
        RECT 3.990 715.040 996.000 719.080 ;
        RECT 3.990 713.680 995.600 715.040 ;
        RECT 4.400 713.640 995.600 713.680 ;
        RECT 4.400 712.280 996.000 713.640 ;
        RECT 3.990 709.600 996.000 712.280 ;
        RECT 3.990 708.200 995.600 709.600 ;
        RECT 3.990 704.160 996.000 708.200 ;
        RECT 4.400 702.760 995.600 704.160 ;
        RECT 3.990 698.720 996.000 702.760 ;
        RECT 3.990 697.320 995.600 698.720 ;
        RECT 3.990 694.640 996.000 697.320 ;
        RECT 4.400 693.280 996.000 694.640 ;
        RECT 4.400 693.240 995.600 693.280 ;
        RECT 3.990 691.880 995.600 693.240 ;
        RECT 3.990 687.840 996.000 691.880 ;
        RECT 3.990 686.440 995.600 687.840 ;
        RECT 3.990 685.120 996.000 686.440 ;
        RECT 4.400 683.720 996.000 685.120 ;
        RECT 3.990 682.400 996.000 683.720 ;
        RECT 3.990 681.000 995.600 682.400 ;
        RECT 3.990 676.960 996.000 681.000 ;
        RECT 3.990 675.600 995.600 676.960 ;
        RECT 4.400 675.560 995.600 675.600 ;
        RECT 4.400 674.200 996.000 675.560 ;
        RECT 3.990 671.520 996.000 674.200 ;
        RECT 3.990 670.120 995.600 671.520 ;
        RECT 3.990 666.080 996.000 670.120 ;
        RECT 4.400 664.680 995.600 666.080 ;
        RECT 3.990 660.640 996.000 664.680 ;
        RECT 3.990 659.240 995.600 660.640 ;
        RECT 3.990 656.560 996.000 659.240 ;
        RECT 4.400 655.200 996.000 656.560 ;
        RECT 4.400 655.160 995.600 655.200 ;
        RECT 3.990 653.800 995.600 655.160 ;
        RECT 3.990 649.760 996.000 653.800 ;
        RECT 3.990 648.360 995.600 649.760 ;
        RECT 3.990 647.040 996.000 648.360 ;
        RECT 4.400 645.640 996.000 647.040 ;
        RECT 3.990 644.320 996.000 645.640 ;
        RECT 3.990 642.920 995.600 644.320 ;
        RECT 3.990 638.880 996.000 642.920 ;
        RECT 3.990 637.520 995.600 638.880 ;
        RECT 4.400 637.480 995.600 637.520 ;
        RECT 4.400 636.120 996.000 637.480 ;
        RECT 3.990 633.440 996.000 636.120 ;
        RECT 3.990 632.040 995.600 633.440 ;
        RECT 3.990 628.000 996.000 632.040 ;
        RECT 4.400 626.600 995.600 628.000 ;
        RECT 3.990 622.560 996.000 626.600 ;
        RECT 3.990 621.160 995.600 622.560 ;
        RECT 3.990 618.480 996.000 621.160 ;
        RECT 4.400 617.120 996.000 618.480 ;
        RECT 4.400 617.080 995.600 617.120 ;
        RECT 3.990 615.720 995.600 617.080 ;
        RECT 3.990 611.680 996.000 615.720 ;
        RECT 3.990 610.280 995.600 611.680 ;
        RECT 3.990 608.960 996.000 610.280 ;
        RECT 4.400 607.560 996.000 608.960 ;
        RECT 3.990 606.240 996.000 607.560 ;
        RECT 3.990 604.840 995.600 606.240 ;
        RECT 3.990 600.800 996.000 604.840 ;
        RECT 3.990 599.440 995.600 600.800 ;
        RECT 4.400 599.400 995.600 599.440 ;
        RECT 4.400 598.040 996.000 599.400 ;
        RECT 3.990 595.360 996.000 598.040 ;
        RECT 3.990 593.960 995.600 595.360 ;
        RECT 3.990 589.920 996.000 593.960 ;
        RECT 4.400 588.520 995.600 589.920 ;
        RECT 3.990 584.480 996.000 588.520 ;
        RECT 3.990 583.080 995.600 584.480 ;
        RECT 3.990 580.400 996.000 583.080 ;
        RECT 4.400 579.040 996.000 580.400 ;
        RECT 4.400 579.000 995.600 579.040 ;
        RECT 3.990 577.640 995.600 579.000 ;
        RECT 3.990 573.600 996.000 577.640 ;
        RECT 3.990 572.200 995.600 573.600 ;
        RECT 3.990 570.880 996.000 572.200 ;
        RECT 4.400 569.480 996.000 570.880 ;
        RECT 3.990 568.160 996.000 569.480 ;
        RECT 3.990 566.760 995.600 568.160 ;
        RECT 3.990 562.720 996.000 566.760 ;
        RECT 3.990 561.360 995.600 562.720 ;
        RECT 4.400 561.320 995.600 561.360 ;
        RECT 4.400 559.960 996.000 561.320 ;
        RECT 3.990 557.280 996.000 559.960 ;
        RECT 3.990 555.880 995.600 557.280 ;
        RECT 3.990 551.840 996.000 555.880 ;
        RECT 4.400 550.440 995.600 551.840 ;
        RECT 3.990 546.400 996.000 550.440 ;
        RECT 3.990 545.000 995.600 546.400 ;
        RECT 3.990 542.320 996.000 545.000 ;
        RECT 4.400 540.960 996.000 542.320 ;
        RECT 4.400 540.920 995.600 540.960 ;
        RECT 3.990 539.560 995.600 540.920 ;
        RECT 3.990 535.520 996.000 539.560 ;
        RECT 3.990 534.120 995.600 535.520 ;
        RECT 3.990 532.800 996.000 534.120 ;
        RECT 4.400 531.400 996.000 532.800 ;
        RECT 3.990 530.080 996.000 531.400 ;
        RECT 3.990 528.680 995.600 530.080 ;
        RECT 3.990 524.640 996.000 528.680 ;
        RECT 3.990 523.280 995.600 524.640 ;
        RECT 4.400 523.240 995.600 523.280 ;
        RECT 4.400 521.880 996.000 523.240 ;
        RECT 3.990 519.200 996.000 521.880 ;
        RECT 3.990 517.800 995.600 519.200 ;
        RECT 3.990 513.760 996.000 517.800 ;
        RECT 4.400 512.360 995.600 513.760 ;
        RECT 3.990 508.320 996.000 512.360 ;
        RECT 3.990 506.920 995.600 508.320 ;
        RECT 3.990 504.240 996.000 506.920 ;
        RECT 4.400 502.880 996.000 504.240 ;
        RECT 4.400 502.840 995.600 502.880 ;
        RECT 3.990 501.480 995.600 502.840 ;
        RECT 3.990 497.440 996.000 501.480 ;
        RECT 3.990 496.040 995.600 497.440 ;
        RECT 3.990 494.720 996.000 496.040 ;
        RECT 4.400 493.320 996.000 494.720 ;
        RECT 3.990 492.000 996.000 493.320 ;
        RECT 3.990 490.600 995.600 492.000 ;
        RECT 3.990 486.560 996.000 490.600 ;
        RECT 3.990 485.200 995.600 486.560 ;
        RECT 4.400 485.160 995.600 485.200 ;
        RECT 4.400 483.800 996.000 485.160 ;
        RECT 3.990 481.120 996.000 483.800 ;
        RECT 3.990 479.720 995.600 481.120 ;
        RECT 3.990 475.680 996.000 479.720 ;
        RECT 4.400 474.280 995.600 475.680 ;
        RECT 3.990 470.240 996.000 474.280 ;
        RECT 3.990 468.840 995.600 470.240 ;
        RECT 3.990 466.160 996.000 468.840 ;
        RECT 4.400 464.800 996.000 466.160 ;
        RECT 4.400 464.760 995.600 464.800 ;
        RECT 3.990 463.400 995.600 464.760 ;
        RECT 3.990 459.360 996.000 463.400 ;
        RECT 3.990 457.960 995.600 459.360 ;
        RECT 3.990 456.640 996.000 457.960 ;
        RECT 4.400 455.240 996.000 456.640 ;
        RECT 3.990 453.920 996.000 455.240 ;
        RECT 3.990 452.520 995.600 453.920 ;
        RECT 3.990 448.480 996.000 452.520 ;
        RECT 3.990 447.120 995.600 448.480 ;
        RECT 4.400 447.080 995.600 447.120 ;
        RECT 4.400 445.720 996.000 447.080 ;
        RECT 3.990 443.040 996.000 445.720 ;
        RECT 3.990 441.640 995.600 443.040 ;
        RECT 3.990 437.600 996.000 441.640 ;
        RECT 4.400 436.200 995.600 437.600 ;
        RECT 3.990 432.160 996.000 436.200 ;
        RECT 3.990 430.760 995.600 432.160 ;
        RECT 3.990 428.080 996.000 430.760 ;
        RECT 4.400 426.720 996.000 428.080 ;
        RECT 4.400 426.680 995.600 426.720 ;
        RECT 3.990 425.320 995.600 426.680 ;
        RECT 3.990 421.280 996.000 425.320 ;
        RECT 3.990 419.880 995.600 421.280 ;
        RECT 3.990 418.560 996.000 419.880 ;
        RECT 4.400 417.160 996.000 418.560 ;
        RECT 3.990 415.840 996.000 417.160 ;
        RECT 3.990 414.440 995.600 415.840 ;
        RECT 3.990 410.400 996.000 414.440 ;
        RECT 3.990 409.040 995.600 410.400 ;
        RECT 4.400 409.000 995.600 409.040 ;
        RECT 4.400 407.640 996.000 409.000 ;
        RECT 3.990 404.960 996.000 407.640 ;
        RECT 3.990 403.560 995.600 404.960 ;
        RECT 3.990 399.520 996.000 403.560 ;
        RECT 4.400 398.120 995.600 399.520 ;
        RECT 3.990 394.080 996.000 398.120 ;
        RECT 3.990 392.680 995.600 394.080 ;
        RECT 3.990 390.000 996.000 392.680 ;
        RECT 4.400 388.640 996.000 390.000 ;
        RECT 4.400 388.600 995.600 388.640 ;
        RECT 3.990 387.240 995.600 388.600 ;
        RECT 3.990 383.200 996.000 387.240 ;
        RECT 3.990 381.800 995.600 383.200 ;
        RECT 3.990 380.480 996.000 381.800 ;
        RECT 4.400 379.080 996.000 380.480 ;
        RECT 3.990 377.760 996.000 379.080 ;
        RECT 3.990 376.360 995.600 377.760 ;
        RECT 3.990 372.320 996.000 376.360 ;
        RECT 3.990 370.960 995.600 372.320 ;
        RECT 4.400 370.920 995.600 370.960 ;
        RECT 4.400 369.560 996.000 370.920 ;
        RECT 3.990 366.880 996.000 369.560 ;
        RECT 3.990 365.480 995.600 366.880 ;
        RECT 3.990 361.440 996.000 365.480 ;
        RECT 4.400 360.040 995.600 361.440 ;
        RECT 3.990 356.000 996.000 360.040 ;
        RECT 3.990 354.600 995.600 356.000 ;
        RECT 3.990 351.920 996.000 354.600 ;
        RECT 4.400 350.560 996.000 351.920 ;
        RECT 4.400 350.520 995.600 350.560 ;
        RECT 3.990 349.160 995.600 350.520 ;
        RECT 3.990 345.120 996.000 349.160 ;
        RECT 3.990 343.720 995.600 345.120 ;
        RECT 3.990 342.400 996.000 343.720 ;
        RECT 4.400 341.000 996.000 342.400 ;
        RECT 3.990 339.680 996.000 341.000 ;
        RECT 3.990 338.280 995.600 339.680 ;
        RECT 3.990 334.240 996.000 338.280 ;
        RECT 3.990 332.880 995.600 334.240 ;
        RECT 4.400 332.840 995.600 332.880 ;
        RECT 4.400 331.480 996.000 332.840 ;
        RECT 3.990 328.800 996.000 331.480 ;
        RECT 3.990 327.400 995.600 328.800 ;
        RECT 3.990 323.360 996.000 327.400 ;
        RECT 4.400 321.960 995.600 323.360 ;
        RECT 3.990 317.920 996.000 321.960 ;
        RECT 3.990 316.520 995.600 317.920 ;
        RECT 3.990 313.840 996.000 316.520 ;
        RECT 4.400 312.480 996.000 313.840 ;
        RECT 4.400 312.440 995.600 312.480 ;
        RECT 3.990 311.080 995.600 312.440 ;
        RECT 3.990 307.040 996.000 311.080 ;
        RECT 3.990 305.640 995.600 307.040 ;
        RECT 3.990 304.320 996.000 305.640 ;
        RECT 4.400 302.920 996.000 304.320 ;
        RECT 3.990 301.600 996.000 302.920 ;
        RECT 3.990 300.200 995.600 301.600 ;
        RECT 3.990 296.160 996.000 300.200 ;
        RECT 3.990 294.800 995.600 296.160 ;
        RECT 4.400 294.760 995.600 294.800 ;
        RECT 4.400 293.400 996.000 294.760 ;
        RECT 3.990 290.720 996.000 293.400 ;
        RECT 3.990 289.320 995.600 290.720 ;
        RECT 3.990 285.280 996.000 289.320 ;
        RECT 4.400 283.880 995.600 285.280 ;
        RECT 3.990 279.840 996.000 283.880 ;
        RECT 3.990 278.440 995.600 279.840 ;
        RECT 3.990 275.760 996.000 278.440 ;
        RECT 4.400 274.400 996.000 275.760 ;
        RECT 4.400 274.360 995.600 274.400 ;
        RECT 3.990 273.000 995.600 274.360 ;
        RECT 3.990 268.960 996.000 273.000 ;
        RECT 3.990 267.560 995.600 268.960 ;
        RECT 3.990 266.240 996.000 267.560 ;
        RECT 4.400 264.840 996.000 266.240 ;
        RECT 3.990 263.520 996.000 264.840 ;
        RECT 3.990 262.120 995.600 263.520 ;
        RECT 3.990 258.080 996.000 262.120 ;
        RECT 3.990 256.720 995.600 258.080 ;
        RECT 4.400 256.680 995.600 256.720 ;
        RECT 4.400 255.320 996.000 256.680 ;
        RECT 3.990 252.640 996.000 255.320 ;
        RECT 3.990 251.240 995.600 252.640 ;
        RECT 3.990 247.200 996.000 251.240 ;
        RECT 4.400 245.800 995.600 247.200 ;
        RECT 3.990 241.760 996.000 245.800 ;
        RECT 3.990 240.360 995.600 241.760 ;
        RECT 3.990 237.680 996.000 240.360 ;
        RECT 4.400 236.320 996.000 237.680 ;
        RECT 4.400 236.280 995.600 236.320 ;
        RECT 3.990 234.920 995.600 236.280 ;
        RECT 3.990 230.880 996.000 234.920 ;
        RECT 3.990 229.480 995.600 230.880 ;
        RECT 3.990 228.160 996.000 229.480 ;
        RECT 4.400 226.760 996.000 228.160 ;
        RECT 3.990 225.440 996.000 226.760 ;
        RECT 3.990 224.040 995.600 225.440 ;
        RECT 3.990 220.000 996.000 224.040 ;
        RECT 3.990 218.640 995.600 220.000 ;
        RECT 4.400 218.600 995.600 218.640 ;
        RECT 4.400 217.240 996.000 218.600 ;
        RECT 3.990 214.560 996.000 217.240 ;
        RECT 3.990 213.160 995.600 214.560 ;
        RECT 3.990 209.120 996.000 213.160 ;
        RECT 4.400 207.720 995.600 209.120 ;
        RECT 3.990 203.680 996.000 207.720 ;
        RECT 3.990 202.280 995.600 203.680 ;
        RECT 3.990 199.600 996.000 202.280 ;
        RECT 4.400 198.240 996.000 199.600 ;
        RECT 4.400 198.200 995.600 198.240 ;
        RECT 3.990 196.840 995.600 198.200 ;
        RECT 3.990 192.800 996.000 196.840 ;
        RECT 3.990 191.400 995.600 192.800 ;
        RECT 3.990 190.080 996.000 191.400 ;
        RECT 4.400 188.680 996.000 190.080 ;
        RECT 3.990 187.360 996.000 188.680 ;
        RECT 3.990 185.960 995.600 187.360 ;
        RECT 3.990 181.920 996.000 185.960 ;
        RECT 3.990 180.560 995.600 181.920 ;
        RECT 4.400 180.520 995.600 180.560 ;
        RECT 4.400 179.160 996.000 180.520 ;
        RECT 3.990 176.480 996.000 179.160 ;
        RECT 3.990 175.080 995.600 176.480 ;
        RECT 3.990 171.040 996.000 175.080 ;
        RECT 4.400 169.640 995.600 171.040 ;
        RECT 3.990 165.600 996.000 169.640 ;
        RECT 3.990 164.200 995.600 165.600 ;
        RECT 3.990 161.520 996.000 164.200 ;
        RECT 4.400 160.160 996.000 161.520 ;
        RECT 4.400 160.120 995.600 160.160 ;
        RECT 3.990 158.760 995.600 160.120 ;
        RECT 3.990 154.720 996.000 158.760 ;
        RECT 3.990 153.320 995.600 154.720 ;
        RECT 3.990 152.000 996.000 153.320 ;
        RECT 4.400 150.600 996.000 152.000 ;
        RECT 3.990 149.280 996.000 150.600 ;
        RECT 3.990 147.880 995.600 149.280 ;
        RECT 3.990 143.840 996.000 147.880 ;
        RECT 3.990 142.480 995.600 143.840 ;
        RECT 4.400 142.440 995.600 142.480 ;
        RECT 4.400 141.080 996.000 142.440 ;
        RECT 3.990 138.400 996.000 141.080 ;
        RECT 3.990 137.000 995.600 138.400 ;
        RECT 3.990 132.960 996.000 137.000 ;
        RECT 4.400 131.560 995.600 132.960 ;
        RECT 3.990 127.520 996.000 131.560 ;
        RECT 3.990 126.120 995.600 127.520 ;
        RECT 3.990 123.440 996.000 126.120 ;
        RECT 4.400 122.080 996.000 123.440 ;
        RECT 4.400 122.040 995.600 122.080 ;
        RECT 3.990 120.680 995.600 122.040 ;
        RECT 3.990 116.640 996.000 120.680 ;
        RECT 3.990 115.240 995.600 116.640 ;
        RECT 3.990 113.920 996.000 115.240 ;
        RECT 4.400 112.520 996.000 113.920 ;
        RECT 3.990 111.200 996.000 112.520 ;
        RECT 3.990 109.800 995.600 111.200 ;
        RECT 3.990 105.760 996.000 109.800 ;
        RECT 3.990 104.400 995.600 105.760 ;
        RECT 4.400 104.360 995.600 104.400 ;
        RECT 4.400 103.000 996.000 104.360 ;
        RECT 3.990 100.320 996.000 103.000 ;
        RECT 3.990 98.920 995.600 100.320 ;
        RECT 3.990 94.880 996.000 98.920 ;
        RECT 4.400 93.480 995.600 94.880 ;
        RECT 3.990 89.440 996.000 93.480 ;
        RECT 3.990 88.040 995.600 89.440 ;
        RECT 3.990 85.360 996.000 88.040 ;
        RECT 4.400 84.000 996.000 85.360 ;
        RECT 4.400 83.960 995.600 84.000 ;
        RECT 3.990 82.600 995.600 83.960 ;
        RECT 3.990 78.560 996.000 82.600 ;
        RECT 3.990 77.160 995.600 78.560 ;
        RECT 3.990 75.840 996.000 77.160 ;
        RECT 4.400 74.440 996.000 75.840 ;
        RECT 3.990 73.120 996.000 74.440 ;
        RECT 3.990 71.720 995.600 73.120 ;
        RECT 3.990 67.680 996.000 71.720 ;
        RECT 3.990 66.320 995.600 67.680 ;
        RECT 4.400 66.280 995.600 66.320 ;
        RECT 4.400 64.920 996.000 66.280 ;
        RECT 3.990 56.800 996.000 64.920 ;
        RECT 4.400 55.400 996.000 56.800 ;
        RECT 3.990 47.280 996.000 55.400 ;
        RECT 4.400 45.880 996.000 47.280 ;
        RECT 3.990 10.715 996.000 45.880 ;
      LAYER met4 ;
        RECT 14.095 11.735 20.640 985.825 ;
        RECT 23.040 11.735 97.440 985.825 ;
        RECT 99.840 11.735 174.240 985.825 ;
        RECT 176.640 11.735 251.040 985.825 ;
        RECT 253.440 11.735 327.840 985.825 ;
        RECT 330.240 11.735 404.640 985.825 ;
        RECT 407.040 11.735 481.440 985.825 ;
        RECT 483.840 11.735 558.240 985.825 ;
        RECT 560.640 11.735 635.040 985.825 ;
        RECT 637.440 11.735 711.840 985.825 ;
        RECT 714.240 11.735 734.785 985.825 ;
  END
END rasterizer_m
END LIBRARY

