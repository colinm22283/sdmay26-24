magic
tech sky130A
magscale 1 2
timestamp 1759434007
<< viali >>
rect 45017 57477 45051 57511
rect 2789 57409 2823 57443
rect 1593 57341 1627 57375
rect 45845 57341 45879 57375
rect 3065 57205 3099 57239
rect 2789 55709 2823 55743
rect 1593 55641 1627 55675
rect 3157 55573 3191 55607
rect 2789 54145 2823 54179
rect 1593 54077 1627 54111
rect 3065 53941 3099 53975
rect 58541 53057 58575 53091
rect 58357 52853 58391 52887
rect 58357 52649 58391 52683
rect 1593 52445 1627 52479
rect 2697 52445 2731 52479
rect 58449 52377 58483 52411
rect 58449 51289 58483 51323
rect 58357 51221 58391 51255
rect 2697 50881 2731 50915
rect 1593 50813 1627 50847
rect 58449 49793 58483 49827
rect 58265 49725 58299 49759
rect 2605 49181 2639 49215
rect 58541 49181 58575 49215
rect 1593 49113 1627 49147
rect 58357 49045 58391 49079
rect 58541 48093 58575 48127
rect 58357 47957 58391 47991
rect 2605 47617 2639 47651
rect 58541 47617 58575 47651
rect 1593 47549 1627 47583
rect 58357 47413 58391 47447
rect 58541 46529 58575 46563
rect 58357 46325 58391 46359
rect 2697 45917 2731 45951
rect 58541 45917 58575 45951
rect 1593 45849 1627 45883
rect 58357 45781 58391 45815
rect 58541 44829 58575 44863
rect 58357 44693 58391 44727
rect 2789 44353 2823 44387
rect 58541 44353 58575 44387
rect 1593 44285 1627 44319
rect 58357 44149 58391 44183
rect 58081 43945 58115 43979
rect 58081 43809 58115 43843
rect 58173 43741 58207 43775
rect 57897 43673 57931 43707
rect 58357 43605 58391 43639
rect 57161 43401 57195 43435
rect 57897 43333 57931 43367
rect 58081 43265 58115 43299
rect 58173 43265 58207 43299
rect 57253 43197 57287 43231
rect 57437 43197 57471 43231
rect 56333 43061 56367 43095
rect 56701 43061 56735 43095
rect 56793 43061 56827 43095
rect 58173 43061 58207 43095
rect 58357 43061 58391 43095
rect 58081 42857 58115 42891
rect 56057 42721 56091 42755
rect 56793 42721 56827 42755
rect 57713 42721 57747 42755
rect 2697 42653 2731 42687
rect 56517 42653 56551 42687
rect 57621 42653 57655 42687
rect 58265 42653 58299 42687
rect 58541 42653 58575 42687
rect 1593 42585 1627 42619
rect 56609 42585 56643 42619
rect 56149 42517 56183 42551
rect 57161 42517 57195 42551
rect 57529 42517 57563 42551
rect 58357 42517 58391 42551
rect 57345 42313 57379 42347
rect 57437 42245 57471 42279
rect 57529 42109 57563 42143
rect 56885 42041 56919 42075
rect 56977 41973 57011 42007
rect 58265 41565 58299 41599
rect 58541 41565 58575 41599
rect 58081 41429 58115 41463
rect 58357 41429 58391 41463
rect 1409 41089 1443 41123
rect 57897 41089 57931 41123
rect 58265 41089 58299 41123
rect 58449 41089 58483 41123
rect 1869 41021 1903 41055
rect 58173 41021 58207 41055
rect 57989 40953 58023 40987
rect 58081 40885 58115 40919
rect 58265 40885 58299 40919
rect 2697 40477 2731 40511
rect 57989 40477 58023 40511
rect 58081 40477 58115 40511
rect 58265 40477 58299 40511
rect 57621 40409 57655 40443
rect 3341 40341 3375 40375
rect 2145 40137 2179 40171
rect 8401 40137 8435 40171
rect 57713 40137 57747 40171
rect 57989 40137 58023 40171
rect 8217 40069 8251 40103
rect 58173 40069 58207 40103
rect 58357 40069 58391 40103
rect 1869 40001 1903 40035
rect 2237 40001 2271 40035
rect 7573 40001 7607 40035
rect 11161 40001 11195 40035
rect 57529 40001 57563 40035
rect 2145 39925 2179 39959
rect 2973 39933 3007 39967
rect 3525 39933 3559 39967
rect 9873 39933 9907 39967
rect 10149 39933 10183 39967
rect 10333 39933 10367 39967
rect 1961 39797 1995 39831
rect 2881 39797 2915 39831
rect 11713 39797 11747 39831
rect 1409 39593 1443 39627
rect 3341 39593 3375 39627
rect 9597 39593 9631 39627
rect 57437 39593 57471 39627
rect 5365 39457 5399 39491
rect 6561 39457 6595 39491
rect 7941 39457 7975 39491
rect 8125 39457 8159 39491
rect 58081 39457 58115 39491
rect 3157 39389 3191 39423
rect 3249 39389 3283 39423
rect 3433 39389 3467 39423
rect 4629 39389 4663 39423
rect 7665 39389 7699 39423
rect 7757 39389 7791 39423
rect 8677 39389 8711 39423
rect 8953 39389 8987 39423
rect 57253 39389 57287 39423
rect 57897 39389 57931 39423
rect 57989 39389 58023 39423
rect 58357 39389 58391 39423
rect 58541 39389 58575 39423
rect 2881 39321 2915 39355
rect 7941 39321 7975 39355
rect 4077 39253 4111 39287
rect 4813 39253 4847 39287
rect 7205 39253 7239 39287
rect 57161 39253 57195 39287
rect 57529 39253 57563 39287
rect 58449 39253 58483 39287
rect 3801 39049 3835 39083
rect 6469 39049 6503 39083
rect 8493 39049 8527 39083
rect 58265 38981 58299 39015
rect 1593 38913 1627 38947
rect 2789 38913 2823 38947
rect 2881 38913 2915 38947
rect 8309 38913 8343 38947
rect 8493 38913 8527 38947
rect 58081 38913 58115 38947
rect 5273 38845 5307 38879
rect 5549 38845 5583 38879
rect 7941 38845 7975 38879
rect 8217 38845 8251 38879
rect 9413 38845 9447 38879
rect 3525 38709 3559 38743
rect 10057 38709 10091 38743
rect 57621 38709 57655 38743
rect 58449 38709 58483 38743
rect 1961 38505 1995 38539
rect 4353 38505 4387 38539
rect 5181 38505 5215 38539
rect 7573 38505 7607 38539
rect 5733 38437 5767 38471
rect 7849 38437 7883 38471
rect 57621 38437 57655 38471
rect 2145 38369 2179 38403
rect 2973 38369 3007 38403
rect 3893 38369 3927 38403
rect 4077 38369 4111 38403
rect 4537 38369 4571 38403
rect 5917 38369 5951 38403
rect 6193 38369 6227 38403
rect 6837 38369 6871 38403
rect 8033 38369 8067 38403
rect 8125 38369 8159 38403
rect 10793 38369 10827 38403
rect 11069 38369 11103 38403
rect 58081 38369 58115 38403
rect 58265 38369 58299 38403
rect 1869 38301 1903 38335
rect 2237 38301 2271 38335
rect 3525 38301 3559 38335
rect 3801 38301 3835 38335
rect 4261 38301 4295 38335
rect 4445 38301 4479 38335
rect 5641 38301 5675 38335
rect 6929 38301 6963 38335
rect 7757 38301 7791 38335
rect 8677 38301 8711 38335
rect 57345 38301 57379 38335
rect 2145 38233 2179 38267
rect 4077 38233 4111 38267
rect 5917 38233 5951 38267
rect 8033 38233 8067 38267
rect 10517 38233 10551 38267
rect 57989 38233 58023 38267
rect 2881 38165 2915 38199
rect 9045 38165 9079 38199
rect 57253 38165 57287 38199
rect 57529 38165 57563 38199
rect 1501 37961 1535 37995
rect 3433 37961 3467 37995
rect 7481 37961 7515 37995
rect 8493 37961 8527 37995
rect 58449 37961 58483 37995
rect 2973 37893 3007 37927
rect 3341 37825 3375 37859
rect 3525 37825 3559 37859
rect 6653 37825 6687 37859
rect 7389 37825 7423 37859
rect 7573 37825 7607 37859
rect 8393 37825 8427 37859
rect 8585 37825 8619 37859
rect 8861 37825 8895 37859
rect 9413 37825 9447 37859
rect 57897 37825 57931 37859
rect 58265 37825 58299 37859
rect 3249 37757 3283 37791
rect 4629 37757 4663 37791
rect 4077 37621 4111 37655
rect 7297 37621 7331 37655
rect 57621 37621 57655 37655
rect 58173 37621 58207 37655
rect 5641 37417 5675 37451
rect 8677 37417 8711 37451
rect 58357 37417 58391 37451
rect 7113 37281 7147 37315
rect 9505 37281 9539 37315
rect 1593 37213 1627 37247
rect 2789 37213 2823 37247
rect 3433 37213 3467 37247
rect 3617 37213 3651 37247
rect 3893 37213 3927 37247
rect 4445 37213 4479 37247
rect 4629 37213 4663 37247
rect 7389 37213 7423 37247
rect 8125 37213 8159 37247
rect 8217 37213 8251 37247
rect 8401 37213 8435 37247
rect 58541 37213 58575 37247
rect 8309 37145 8343 37179
rect 3525 37077 3559 37111
rect 5273 37077 5307 37111
rect 7481 37077 7515 37111
rect 8953 37077 8987 37111
rect 7665 36873 7699 36907
rect 2237 36805 2271 36839
rect 5457 36805 5491 36839
rect 6929 36805 6963 36839
rect 8493 36805 8527 36839
rect 1961 36737 1995 36771
rect 2329 36737 2363 36771
rect 5733 36737 5767 36771
rect 6653 36737 6687 36771
rect 7021 36737 7055 36771
rect 10517 36737 10551 36771
rect 10793 36737 10827 36771
rect 57897 36737 57931 36771
rect 58081 36737 58115 36771
rect 58541 36737 58575 36771
rect 2237 36669 2271 36703
rect 3065 36669 3099 36703
rect 3617 36669 3651 36703
rect 3985 36669 4019 36703
rect 6929 36669 6963 36703
rect 8401 36669 8435 36703
rect 10241 36669 10275 36703
rect 2053 36533 2087 36567
rect 2973 36533 3007 36567
rect 6745 36533 6779 36567
rect 7757 36533 7791 36567
rect 57713 36533 57747 36567
rect 57989 36533 58023 36567
rect 58357 36533 58391 36567
rect 1409 36329 1443 36363
rect 3341 36329 3375 36363
rect 3985 36329 4019 36363
rect 8585 36329 8619 36363
rect 9965 36329 9999 36363
rect 57529 36261 57563 36295
rect 2881 36193 2915 36227
rect 3157 36193 3191 36227
rect 4077 36193 4111 36227
rect 8125 36193 8159 36227
rect 8309 36193 8343 36227
rect 3249 36135 3283 36169
rect 3433 36125 3467 36159
rect 3801 36125 3835 36159
rect 3893 36125 3927 36159
rect 4537 36125 4571 36159
rect 7205 36125 7239 36159
rect 8033 36125 8067 36159
rect 8493 36125 8527 36159
rect 8677 36125 8711 36159
rect 9321 36125 9355 36159
rect 57713 36125 57747 36159
rect 57805 36125 57839 36159
rect 58541 36125 58575 36159
rect 8309 36057 8343 36091
rect 57529 36057 57563 36091
rect 5181 35989 5215 36023
rect 7849 35989 7883 36023
rect 58357 35989 58391 36023
rect 3525 35785 3559 35819
rect 4353 35785 4387 35819
rect 6193 35785 6227 35819
rect 6469 35785 6503 35819
rect 4721 35717 4755 35751
rect 7941 35717 7975 35751
rect 8309 35717 8343 35751
rect 58265 35717 58299 35751
rect 1593 35649 1627 35683
rect 2789 35649 2823 35683
rect 2881 35649 2915 35683
rect 4077 35649 4111 35683
rect 4445 35649 4479 35683
rect 9229 35649 9263 35683
rect 58081 35649 58115 35683
rect 58173 35649 58207 35683
rect 58449 35649 58483 35683
rect 4353 35581 4387 35615
rect 8217 35581 8251 35615
rect 8861 35581 8895 35615
rect 4169 35445 4203 35479
rect 57621 35445 57655 35479
rect 57897 35445 57931 35479
rect 3433 35241 3467 35275
rect 3893 35241 3927 35275
rect 4721 35241 4755 35275
rect 7389 35241 7423 35275
rect 57437 35241 57471 35275
rect 58357 35241 58391 35275
rect 7297 35173 7331 35207
rect 57897 35173 57931 35207
rect 5365 35105 5399 35139
rect 5549 35105 5583 35139
rect 6285 35105 6319 35139
rect 7481 35105 7515 35139
rect 7757 35105 7791 35139
rect 8401 35105 8435 35139
rect 8585 35105 8619 35139
rect 56241 35105 56275 35139
rect 57621 35105 57655 35139
rect 2513 35037 2547 35071
rect 3341 35037 3375 35071
rect 3525 35037 3559 35071
rect 3801 35037 3835 35071
rect 3985 35037 4019 35071
rect 5457 35037 5491 35071
rect 5641 35037 5675 35071
rect 5733 35037 5767 35071
rect 7205 35037 7239 35071
rect 8493 35037 8527 35071
rect 8677 35037 8711 35071
rect 55597 35037 55631 35071
rect 55781 35037 55815 35071
rect 55873 35037 55907 35071
rect 56057 35037 56091 35071
rect 56149 35037 56183 35071
rect 56341 35037 56375 35071
rect 57069 35037 57103 35071
rect 57253 35037 57287 35071
rect 57345 35037 57379 35071
rect 57989 35037 58023 35071
rect 58173 35037 58207 35071
rect 58541 35037 58575 35071
rect 57161 34969 57195 35003
rect 3065 34901 3099 34935
rect 55597 34901 55631 34935
rect 55965 34901 55999 34935
rect 56885 34901 56919 34935
rect 57989 34901 58023 34935
rect 1409 34697 1443 34731
rect 4537 34697 4571 34731
rect 49341 34697 49375 34731
rect 55781 34697 55815 34731
rect 56517 34697 56551 34731
rect 2881 34629 2915 34663
rect 3249 34629 3283 34663
rect 57253 34629 57287 34663
rect 4077 34561 4111 34595
rect 4261 34561 4295 34595
rect 4537 34561 4571 34595
rect 4721 34561 4755 34595
rect 51181 34561 51215 34595
rect 51917 34561 51951 34595
rect 55689 34561 55723 34595
rect 55873 34561 55907 34595
rect 56333 34561 56367 34595
rect 56609 34561 56643 34595
rect 56701 34561 56735 34595
rect 56885 34561 56919 34595
rect 57437 34561 57471 34595
rect 57621 34561 57655 34595
rect 58541 34561 58575 34595
rect 3157 34493 3191 34527
rect 3801 34493 3835 34527
rect 50813 34493 50847 34527
rect 51089 34493 51123 34527
rect 57713 34493 57747 34527
rect 4169 34425 4203 34459
rect 56793 34425 56827 34459
rect 51365 34357 51399 34391
rect 52009 34357 52043 34391
rect 56333 34357 56367 34391
rect 58357 34357 58391 34391
rect 3065 34153 3099 34187
rect 7021 34153 7055 34187
rect 50813 34153 50847 34187
rect 57989 34153 58023 34187
rect 58173 34153 58207 34187
rect 3801 34085 3835 34119
rect 1593 34017 1627 34051
rect 3157 34017 3191 34051
rect 3341 34017 3375 34051
rect 4353 34017 4387 34051
rect 57345 34017 57379 34051
rect 2605 33949 2639 33983
rect 2881 33949 2915 33983
rect 2973 33949 3007 33983
rect 3249 33949 3283 33983
rect 3433 33949 3467 33983
rect 5365 33949 5399 33983
rect 5457 33949 5491 33983
rect 5641 33949 5675 33983
rect 9321 33949 9355 33983
rect 41613 33949 41647 33983
rect 45661 33949 45695 33983
rect 50169 33949 50203 33983
rect 57253 33949 57287 33983
rect 57437 33949 57471 33983
rect 5908 33881 5942 33915
rect 9566 33881 9600 33915
rect 41889 33881 41923 33915
rect 43453 33881 43487 33915
rect 44189 33881 44223 33915
rect 44741 33881 44775 33915
rect 58357 33881 58391 33915
rect 5273 33813 5307 33847
rect 7389 33813 7423 33847
rect 10701 33813 10735 33847
rect 43361 33813 43395 33847
rect 45477 33813 45511 33847
rect 46397 33813 46431 33847
rect 57805 33813 57839 33847
rect 58147 33813 58181 33847
rect 3249 33609 3283 33643
rect 4997 33609 5031 33643
rect 5923 33609 5957 33643
rect 8677 33609 8711 33643
rect 9781 33609 9815 33643
rect 42441 33609 42475 33643
rect 44281 33609 44315 33643
rect 44557 33609 44591 33643
rect 49617 33609 49651 33643
rect 50169 33609 50203 33643
rect 55689 33609 55723 33643
rect 56793 33609 56827 33643
rect 5273 33541 5307 33575
rect 5549 33541 5583 33575
rect 5825 33541 5859 33575
rect 42165 33541 42199 33575
rect 46857 33541 46891 33575
rect 50675 33541 50709 33575
rect 3341 33473 3375 33507
rect 3884 33473 3918 33507
rect 5089 33473 5123 33507
rect 5365 33473 5399 33507
rect 5457 33473 5491 33507
rect 5641 33473 5675 33507
rect 6009 33473 6043 33507
rect 6101 33473 6135 33507
rect 6377 33473 6411 33507
rect 6561 33473 6595 33507
rect 6745 33473 6779 33507
rect 7021 33473 7055 33507
rect 7205 33473 7239 33507
rect 7564 33473 7598 33507
rect 9137 33473 9171 33507
rect 9321 33473 9355 33507
rect 9413 33473 9447 33507
rect 9689 33473 9723 33507
rect 9781 33473 9815 33507
rect 9965 33473 9999 33507
rect 42257 33473 42291 33507
rect 43177 33473 43211 33507
rect 43361 33473 43395 33507
rect 43453 33473 43487 33507
rect 44189 33473 44223 33507
rect 46489 33473 46523 33507
rect 47593 33473 47627 33507
rect 49433 33473 49467 33507
rect 50353 33473 50387 33507
rect 50445 33473 50479 33507
rect 50537 33473 50571 33507
rect 51089 33473 51123 33507
rect 51273 33473 51307 33507
rect 51365 33473 51399 33507
rect 51457 33473 51491 33507
rect 51641 33473 51675 33507
rect 51733 33473 51767 33507
rect 52009 33473 52043 33507
rect 52193 33473 52227 33507
rect 55505 33473 55539 33507
rect 55781 33473 55815 33507
rect 57345 33473 57379 33507
rect 57897 33473 57931 33507
rect 58081 33473 58115 33507
rect 58541 33473 58575 33507
rect 3433 33405 3467 33439
rect 3617 33405 3651 33439
rect 6469 33405 6503 33439
rect 6837 33405 6871 33439
rect 7297 33405 7331 33439
rect 9597 33405 9631 33439
rect 41797 33405 41831 33439
rect 41981 33405 42015 33439
rect 42993 33405 43027 33439
rect 44097 33405 44131 33439
rect 46029 33405 46063 33439
rect 46305 33405 46339 33439
rect 47869 33405 47903 33439
rect 49341 33405 49375 33439
rect 50813 33405 50847 33439
rect 52101 33405 52135 33439
rect 57437 33405 57471 33439
rect 57529 33405 57563 33439
rect 5089 33337 5123 33371
rect 10333 33337 10367 33371
rect 51549 33337 51583 33371
rect 58357 33337 58391 33371
rect 7113 33269 7147 33303
rect 9137 33269 9171 33303
rect 10609 33269 10643 33303
rect 43269 33269 43303 33303
rect 50905 33269 50939 33303
rect 51825 33269 51859 33303
rect 52561 33269 52595 33303
rect 55505 33269 55539 33303
rect 56977 33269 57011 33303
rect 57989 33269 58023 33303
rect 7757 33065 7791 33099
rect 45937 33065 45971 33099
rect 46213 33065 46247 33099
rect 48145 33065 48179 33099
rect 57345 33065 57379 33099
rect 42073 32997 42107 33031
rect 44557 32997 44591 33031
rect 45109 32997 45143 33031
rect 48053 32997 48087 33031
rect 49433 32997 49467 33031
rect 56425 32997 56459 33031
rect 40325 32929 40359 32963
rect 44189 32929 44223 32963
rect 44362 32929 44396 32963
rect 2605 32861 2639 32895
rect 2881 32861 2915 32895
rect 7481 32861 7515 32895
rect 7757 32861 7791 32895
rect 42717 32861 42751 32895
rect 43545 32861 43579 32895
rect 44649 32861 44683 32895
rect 45017 32861 45051 32895
rect 45293 32861 45327 32895
rect 47869 32861 47903 32895
rect 48053 32861 48087 32895
rect 48789 32861 48823 32895
rect 48881 32861 48915 32895
rect 49065 32861 49099 32895
rect 49249 32861 49283 32895
rect 49341 32861 49375 32895
rect 49709 32861 49743 32895
rect 49985 32861 50019 32895
rect 56333 32861 56367 32895
rect 56517 32861 56551 32895
rect 56609 32861 56643 32895
rect 56793 32861 56827 32895
rect 57253 32861 57287 32895
rect 57437 32861 57471 32895
rect 58541 32861 58575 32895
rect 1593 32793 1627 32827
rect 40601 32793 40635 32827
rect 43637 32793 43671 32827
rect 44373 32793 44407 32827
rect 49433 32793 49467 32827
rect 49617 32793 49651 32827
rect 56701 32793 56735 32827
rect 3525 32725 3559 32759
rect 4905 32725 4939 32759
rect 5825 32725 5859 32759
rect 6745 32725 6779 32759
rect 7297 32725 7331 32759
rect 7573 32725 7607 32759
rect 42165 32725 42199 32759
rect 42901 32725 42935 32759
rect 49893 32725 49927 32759
rect 51273 32725 51307 32759
rect 58357 32725 58391 32759
rect 1409 32521 1443 32555
rect 3985 32521 4019 32555
rect 4813 32521 4847 32555
rect 8125 32521 8159 32555
rect 8585 32521 8619 32555
rect 38393 32521 38427 32555
rect 41337 32521 41371 32555
rect 42441 32521 42475 32555
rect 42901 32521 42935 32555
rect 44097 32453 44131 32487
rect 44189 32453 44223 32487
rect 44557 32453 44591 32487
rect 45201 32453 45235 32487
rect 58265 32453 58299 32487
rect 3985 32385 4019 32419
rect 4169 32385 4203 32419
rect 4261 32385 4295 32419
rect 4445 32385 4479 32419
rect 4537 32385 4571 32419
rect 4721 32385 4755 32419
rect 5926 32385 5960 32419
rect 8217 32385 8251 32419
rect 8401 32385 8435 32419
rect 8493 32385 8527 32419
rect 8769 32385 8803 32419
rect 9974 32385 10008 32419
rect 39037 32385 39071 32419
rect 39221 32385 39255 32419
rect 39313 32385 39347 32419
rect 39497 32385 39531 32419
rect 41521 32385 41555 32419
rect 42625 32385 42659 32419
rect 42809 32385 42843 32419
rect 42901 32385 42935 32419
rect 43085 32385 43119 32419
rect 43913 32385 43947 32419
rect 44281 32385 44315 32419
rect 44833 32385 44867 32419
rect 45109 32385 45143 32419
rect 45293 32385 45327 32419
rect 47409 32385 47443 32419
rect 47869 32385 47903 32419
rect 48881 32385 48915 32419
rect 49065 32385 49099 32419
rect 52837 32385 52871 32419
rect 53021 32385 53055 32419
rect 53849 32385 53883 32419
rect 58357 32385 58391 32419
rect 2881 32317 2915 32351
rect 3157 32317 3191 32351
rect 3801 32317 3835 32351
rect 6193 32317 6227 32351
rect 10241 32317 10275 32351
rect 40601 32317 40635 32351
rect 44649 32317 44683 32351
rect 47041 32317 47075 32351
rect 47593 32317 47627 32351
rect 52929 32317 52963 32351
rect 53665 32317 53699 32351
rect 54401 32317 54435 32351
rect 55597 32317 55631 32351
rect 8309 32249 8343 32283
rect 8769 32249 8803 32283
rect 44465 32249 44499 32283
rect 3249 32181 3283 32215
rect 4353 32181 4387 32215
rect 4629 32181 4663 32215
rect 6653 32181 6687 32215
rect 8861 32181 8895 32215
rect 10609 32181 10643 32215
rect 39129 32181 39163 32215
rect 39405 32181 39439 32215
rect 41245 32181 41279 32215
rect 44741 32181 44775 32215
rect 45017 32181 45051 32215
rect 45615 32181 45649 32215
rect 48973 32181 49007 32215
rect 53113 32181 53147 32215
rect 55045 32181 55079 32215
rect 3341 31977 3375 32011
rect 4997 31977 5031 32011
rect 6285 31977 6319 32011
rect 6469 31977 6503 32011
rect 8401 31977 8435 32011
rect 39681 31977 39715 32011
rect 42073 31977 42107 32011
rect 42441 31977 42475 32011
rect 44373 31977 44407 32011
rect 45753 31977 45787 32011
rect 46857 31977 46891 32011
rect 50629 31977 50663 32011
rect 53941 31977 53975 32011
rect 55045 31977 55079 32011
rect 2329 31909 2363 31943
rect 6653 31909 6687 31943
rect 10333 31909 10367 31943
rect 38301 31909 38335 31943
rect 43177 31909 43211 31943
rect 45845 31909 45879 31943
rect 46673 31909 46707 31943
rect 52193 31909 52227 31943
rect 2421 31841 2455 31875
rect 2697 31841 2731 31875
rect 8033 31841 8067 31875
rect 38853 31841 38887 31875
rect 39865 31841 39899 31875
rect 41337 31841 41371 31875
rect 41613 31841 41647 31875
rect 42809 31841 42843 31875
rect 42993 31841 43027 31875
rect 45937 31841 45971 31875
rect 47133 31841 47167 31875
rect 48973 31841 49007 31875
rect 49249 31841 49283 31875
rect 49433 31841 49467 31875
rect 49893 31841 49927 31875
rect 52377 31841 52411 31875
rect 55321 31841 55355 31875
rect 2145 31773 2179 31807
rect 2237 31773 2271 31807
rect 3433 31773 3467 31807
rect 3617 31773 3651 31807
rect 4721 31773 4755 31807
rect 4813 31773 4847 31807
rect 6367 31773 6401 31807
rect 6561 31773 6595 31807
rect 10057 31773 10091 31807
rect 10241 31773 10275 31807
rect 10517 31773 10551 31807
rect 10773 31773 10807 31807
rect 36277 31773 36311 31807
rect 36461 31773 36495 31807
rect 39129 31773 39163 31807
rect 39497 31773 39531 31807
rect 42533 31773 42567 31807
rect 43084 31751 43118 31785
rect 43545 31773 43579 31807
rect 43637 31773 43671 31807
rect 44005 31773 44039 31807
rect 44281 31773 44315 31807
rect 45569 31773 45603 31807
rect 45661 31773 45695 31807
rect 46029 31773 46063 31807
rect 46765 31773 46799 31807
rect 47041 31773 47075 31807
rect 47225 31773 47259 31807
rect 47317 31773 47351 31807
rect 47501 31773 47535 31807
rect 48881 31773 48915 31807
rect 49065 31773 49099 31807
rect 49525 31773 49559 31807
rect 49801 31773 49835 31807
rect 49985 31773 50019 31807
rect 52009 31773 52043 31807
rect 52101 31773 52135 31807
rect 52561 31773 52595 31807
rect 54953 31773 54987 31807
rect 55137 31773 55171 31807
rect 56793 31773 56827 31807
rect 58541 31773 58575 31807
rect 4997 31705 5031 31739
rect 7766 31705 7800 31739
rect 36737 31705 36771 31739
rect 38761 31705 38795 31739
rect 39313 31705 39347 31739
rect 39405 31705 39439 31739
rect 43177 31705 43211 31739
rect 51764 31705 51798 31739
rect 52377 31705 52411 31739
rect 52828 31705 52862 31739
rect 55566 31705 55600 31739
rect 57038 31705 57072 31739
rect 3525 31637 3559 31671
rect 11897 31637 11931 31671
rect 38209 31637 38243 31671
rect 38669 31637 38703 31671
rect 42809 31637 42843 31671
rect 47409 31637 47443 31671
rect 49249 31637 49283 31671
rect 56701 31637 56735 31671
rect 58173 31637 58207 31671
rect 58357 31637 58391 31671
rect 4905 31433 4939 31467
rect 6009 31433 6043 31467
rect 8493 31433 8527 31467
rect 36921 31433 36955 31467
rect 38301 31433 38335 31467
rect 39129 31433 39163 31467
rect 39589 31433 39623 31467
rect 47317 31433 47351 31467
rect 52469 31433 52503 31467
rect 53113 31433 53147 31467
rect 54953 31433 54987 31467
rect 56793 31433 56827 31467
rect 5089 31365 5123 31399
rect 8861 31365 8895 31399
rect 46089 31365 46123 31399
rect 46305 31365 46339 31399
rect 48237 31365 48271 31399
rect 57897 31365 57931 31399
rect 2697 31297 2731 31331
rect 3893 31297 3927 31331
rect 4077 31297 4111 31331
rect 4169 31297 4203 31331
rect 4353 31297 4387 31331
rect 5273 31297 5307 31331
rect 6009 31297 6043 31331
rect 6193 31297 6227 31331
rect 6929 31297 6963 31331
rect 7021 31297 7055 31331
rect 7205 31297 7239 31331
rect 8493 31297 8527 31331
rect 8677 31297 8711 31331
rect 8769 31297 8803 31331
rect 8953 31297 8987 31331
rect 12633 31297 12667 31331
rect 37105 31297 37139 31331
rect 38209 31297 38243 31331
rect 38485 31297 38519 31331
rect 39221 31297 39255 31331
rect 39405 31297 39439 31331
rect 40233 31297 40267 31331
rect 41245 31297 41279 31331
rect 41705 31297 41739 31331
rect 47225 31297 47259 31331
rect 48053 31297 48087 31331
rect 48329 31297 48363 31331
rect 48605 31297 48639 31331
rect 49157 31297 49191 31331
rect 51089 31297 51123 31331
rect 52837 31297 52871 31331
rect 54585 31297 54619 31331
rect 54677 31297 54711 31331
rect 55229 31297 55263 31331
rect 56241 31297 56275 31331
rect 56425 31297 56459 31331
rect 56517 31297 56551 31331
rect 58449 31297 58483 31331
rect 1593 31229 1627 31263
rect 3709 31229 3743 31263
rect 6561 31229 6595 31263
rect 13461 31229 13495 31263
rect 40969 31229 41003 31263
rect 43821 31229 43855 31263
rect 44097 31229 44131 31263
rect 45845 31229 45879 31263
rect 48881 31229 48915 31263
rect 51825 31229 51859 31263
rect 53113 31229 53147 31263
rect 54953 31229 54987 31263
rect 55873 31229 55907 31263
rect 56793 31229 56827 31263
rect 56885 31229 56919 31263
rect 57437 31229 57471 31263
rect 5641 31161 5675 31195
rect 39681 31161 39715 31195
rect 56333 31161 56367 31195
rect 3157 31093 3191 31127
rect 3985 31093 4019 31127
rect 4261 31093 4295 31127
rect 7205 31093 7239 31127
rect 9229 31093 9263 31127
rect 9597 31093 9631 31127
rect 45937 31093 45971 31127
rect 46121 31093 46155 31127
rect 47869 31093 47903 31127
rect 48697 31093 48731 31127
rect 48789 31093 48823 31127
rect 49065 31093 49099 31127
rect 51733 31093 51767 31127
rect 52929 31093 52963 31127
rect 54493 31093 54527 31127
rect 54769 31093 54803 31127
rect 56609 31093 56643 31127
rect 3433 30889 3467 30923
rect 7113 30889 7147 30923
rect 9045 30889 9079 30923
rect 9321 30889 9355 30923
rect 10701 30889 10735 30923
rect 38117 30889 38151 30923
rect 38669 30889 38703 30923
rect 39957 30889 39991 30923
rect 44649 30889 44683 30923
rect 48513 30889 48547 30923
rect 51457 30889 51491 30923
rect 42257 30821 42291 30855
rect 45753 30821 45787 30855
rect 58265 30821 58299 30855
rect 2881 30753 2915 30787
rect 3157 30753 3191 30787
rect 3525 30753 3559 30787
rect 3801 30753 3835 30787
rect 4445 30753 4479 30787
rect 39865 30753 39899 30787
rect 41337 30753 41371 30787
rect 43821 30753 43855 30787
rect 44005 30753 44039 30787
rect 48421 30753 48455 30787
rect 49065 30753 49099 30787
rect 49249 30753 49283 30787
rect 57253 30753 57287 30787
rect 57437 30753 57471 30787
rect 3249 30685 3283 30719
rect 3341 30685 3375 30719
rect 4537 30685 4571 30719
rect 6101 30685 6135 30719
rect 7021 30685 7055 30719
rect 7205 30685 7239 30719
rect 8953 30685 8987 30719
rect 9137 30685 9171 30719
rect 9229 30685 9263 30719
rect 9413 30685 9447 30719
rect 9689 30685 9723 30719
rect 9873 30685 9907 30719
rect 9965 30685 9999 30719
rect 38485 30685 38519 30719
rect 38761 30685 38795 30719
rect 40049 30685 40083 30719
rect 40141 30685 40175 30719
rect 42073 30685 42107 30719
rect 42993 30685 43027 30719
rect 43729 30685 43763 30719
rect 43913 30685 43947 30719
rect 45477 30685 45511 30719
rect 45569 30685 45603 30719
rect 46673 30685 46707 30719
rect 51365 30685 51399 30719
rect 51549 30685 51583 30719
rect 53113 30685 53147 30719
rect 53205 30685 53239 30719
rect 53297 30685 53331 30719
rect 54309 30685 54343 30719
rect 54401 30685 54435 30719
rect 56977 30685 57011 30719
rect 57069 30685 57103 30719
rect 57345 30685 57379 30719
rect 57529 30685 57563 30719
rect 57897 30685 57931 30719
rect 58357 30685 58391 30719
rect 4813 30617 4847 30651
rect 7573 30617 7607 30651
rect 8677 30617 8711 30651
rect 10149 30617 10183 30651
rect 12173 30617 12207 30651
rect 12541 30617 12575 30651
rect 15669 30617 15703 30651
rect 17417 30617 17451 30651
rect 38301 30617 38335 30651
rect 41981 30617 42015 30651
rect 45753 30617 45787 30651
rect 46949 30617 46983 30651
rect 54125 30617 54159 30651
rect 1409 30549 1443 30583
rect 5365 30549 5399 30583
rect 6193 30549 6227 30583
rect 6561 30549 6595 30583
rect 9873 30549 9907 30583
rect 10333 30549 10367 30583
rect 17693 30549 17727 30583
rect 43085 30549 43119 30583
rect 46029 30549 46063 30583
rect 49893 30549 49927 30583
rect 53481 30549 53515 30583
rect 54309 30549 54343 30583
rect 57253 30549 57287 30583
rect 58081 30549 58115 30583
rect 3341 30345 3375 30379
rect 5463 30345 5497 30379
rect 10241 30345 10275 30379
rect 10701 30345 10735 30379
rect 12909 30345 12943 30379
rect 39957 30345 39991 30379
rect 43729 30345 43763 30379
rect 46489 30345 46523 30379
rect 2605 30277 2639 30311
rect 5028 30277 5062 30311
rect 5825 30277 5859 30311
rect 10425 30277 10459 30311
rect 41981 30277 42015 30311
rect 42441 30277 42475 30311
rect 48697 30277 48731 30311
rect 50445 30277 50479 30311
rect 51825 30277 51859 30311
rect 53021 30277 53055 30311
rect 57621 30277 57655 30311
rect 2697 30209 2731 30243
rect 3433 30209 3467 30243
rect 5365 30209 5399 30243
rect 5549 30209 5583 30243
rect 5641 30209 5675 30243
rect 5733 30209 5767 30243
rect 5917 30209 5951 30243
rect 6377 30209 6411 30243
rect 6644 30209 6678 30243
rect 10149 30209 10183 30243
rect 10514 30209 10548 30243
rect 10793 30209 10827 30243
rect 10885 30199 10919 30233
rect 11069 30209 11103 30243
rect 11785 30209 11819 30243
rect 38853 30209 38887 30243
rect 39221 30209 39255 30243
rect 39405 30209 39439 30243
rect 40141 30209 40175 30243
rect 43269 30209 43303 30243
rect 43361 30209 43395 30243
rect 43637 30209 43671 30243
rect 43913 30209 43947 30243
rect 44097 30209 44131 30243
rect 44189 30209 44223 30243
rect 45661 30209 45695 30243
rect 48421 30209 48455 30243
rect 51457 30209 51491 30243
rect 51549 30209 51583 30243
rect 51641 30215 51675 30249
rect 51917 30209 51951 30243
rect 52101 30209 52135 30243
rect 52193 30209 52227 30243
rect 52377 30209 52411 30243
rect 52929 30209 52963 30243
rect 53113 30209 53147 30243
rect 53297 30209 53331 30243
rect 53481 30209 53515 30243
rect 54309 30209 54343 30243
rect 54493 30209 54527 30243
rect 54769 30209 54803 30243
rect 54953 30209 54987 30243
rect 55229 30209 55263 30243
rect 57529 30209 57563 30243
rect 57897 30209 57931 30243
rect 58173 30209 58207 30243
rect 3709 30141 3743 30175
rect 5273 30141 5307 30175
rect 11529 30141 11563 30175
rect 40509 30141 40543 30175
rect 42257 30141 42291 30175
rect 43085 30141 43119 30175
rect 45569 30141 45603 30175
rect 47041 30141 47075 30175
rect 50721 30141 50755 30175
rect 52009 30141 52043 30175
rect 3525 30073 3559 30107
rect 10425 30073 10459 30107
rect 38761 30073 38795 30107
rect 43177 30073 43211 30107
rect 45293 30073 45327 30107
rect 46305 30073 46339 30107
rect 58265 30073 58299 30107
rect 3617 30005 3651 30039
rect 3893 30005 3927 30039
rect 7757 30005 7791 30039
rect 9505 30005 9539 30039
rect 10517 30005 10551 30039
rect 10977 30005 11011 30039
rect 39405 30005 39439 30039
rect 43545 30005 43579 30039
rect 45109 30005 45143 30039
rect 45661 30005 45695 30039
rect 45937 30005 45971 30039
rect 47869 30005 47903 30039
rect 52285 30005 52319 30039
rect 53389 30005 53423 30039
rect 54401 30005 54435 30039
rect 54861 30005 54895 30039
rect 55873 30005 55907 30039
rect 58081 30005 58115 30039
rect 3801 29801 3835 29835
rect 4629 29801 4663 29835
rect 6009 29801 6043 29835
rect 6561 29801 6595 29835
rect 15853 29801 15887 29835
rect 40049 29801 40083 29835
rect 43269 29801 43303 29835
rect 43729 29801 43763 29835
rect 46765 29801 46799 29835
rect 50905 29801 50939 29835
rect 51365 29801 51399 29835
rect 55045 29801 55079 29835
rect 57529 29801 57563 29835
rect 9781 29733 9815 29767
rect 41797 29733 41831 29767
rect 47317 29733 47351 29767
rect 50169 29733 50203 29767
rect 3617 29665 3651 29699
rect 7021 29665 7055 29699
rect 8125 29665 8159 29699
rect 9137 29665 9171 29699
rect 37289 29665 37323 29699
rect 37381 29665 37415 29699
rect 39589 29665 39623 29699
rect 45017 29665 45051 29699
rect 47501 29665 47535 29699
rect 47777 29665 47811 29699
rect 50721 29665 50755 29699
rect 51181 29665 51215 29699
rect 54033 29665 54067 29699
rect 56701 29665 56735 29699
rect 2605 29597 2639 29631
rect 4445 29597 4479 29631
rect 4537 29597 4571 29631
rect 4721 29597 4755 29631
rect 6837 29597 6871 29631
rect 6929 29597 6963 29631
rect 7113 29597 7147 29631
rect 8677 29597 8711 29631
rect 9413 29597 9447 29631
rect 10609 29597 10643 29631
rect 10793 29597 10827 29631
rect 11897 29597 11931 29631
rect 15485 29597 15519 29631
rect 39497 29597 39531 29631
rect 39681 29597 39715 29631
rect 39957 29597 39991 29631
rect 40141 29597 40175 29631
rect 41981 29597 42015 29631
rect 42441 29597 42475 29631
rect 42993 29597 43027 29631
rect 43177 29597 43211 29631
rect 43361 29597 43395 29631
rect 44097 29597 44131 29631
rect 46857 29597 46891 29631
rect 47041 29597 47075 29631
rect 51089 29597 51123 29631
rect 51457 29597 51491 29631
rect 51733 29597 51767 29631
rect 52009 29597 52043 29631
rect 52193 29597 52227 29631
rect 52293 29597 52327 29631
rect 52469 29597 52503 29631
rect 53021 29597 53055 29631
rect 53205 29597 53239 29631
rect 53297 29597 53331 29631
rect 53481 29597 53515 29631
rect 53573 29597 53607 29631
rect 53757 29597 53791 29631
rect 54953 29597 54987 29631
rect 55137 29597 55171 29631
rect 56977 29597 57011 29631
rect 57161 29597 57195 29631
rect 57713 29597 57747 29631
rect 57897 29597 57931 29631
rect 1593 29529 1627 29563
rect 6561 29529 6595 29563
rect 12449 29529 12483 29563
rect 37657 29529 37691 29563
rect 43913 29529 43947 29563
rect 45293 29529 45327 29563
rect 51365 29529 51399 29563
rect 52101 29529 52135 29563
rect 53113 29529 53147 29563
rect 53665 29529 53699 29563
rect 56434 29529 56468 29563
rect 58265 29529 58299 29563
rect 2973 29461 3007 29495
rect 6745 29461 6779 29495
rect 10793 29461 10827 29495
rect 15393 29461 15427 29495
rect 39129 29461 39163 29495
rect 46949 29461 46983 29495
rect 49249 29461 49283 29495
rect 52285 29461 52319 29495
rect 52837 29461 52871 29495
rect 53389 29461 53423 29495
rect 55321 29461 55355 29495
rect 57069 29461 57103 29495
rect 1409 29257 1443 29291
rect 5825 29257 5859 29291
rect 6561 29257 6595 29291
rect 8953 29257 8987 29291
rect 10694 29257 10728 29291
rect 11621 29257 11655 29291
rect 40049 29257 40083 29291
rect 45477 29257 45511 29291
rect 48605 29257 48639 29291
rect 51457 29257 51491 29291
rect 53021 29257 53055 29291
rect 53481 29257 53515 29291
rect 55229 29257 55263 29291
rect 55965 29257 55999 29291
rect 56885 29257 56919 29291
rect 2881 29189 2915 29223
rect 4712 29189 4746 29223
rect 10180 29189 10214 29223
rect 10977 29189 11011 29223
rect 11161 29189 11195 29223
rect 37749 29189 37783 29223
rect 43545 29189 43579 29223
rect 54861 29189 54895 29223
rect 57345 29189 57379 29223
rect 3157 29121 3191 29155
rect 3341 29121 3375 29155
rect 4169 29121 4203 29155
rect 4353 29121 4387 29155
rect 6469 29121 6503 29155
rect 6745 29121 6779 29155
rect 10517 29121 10551 29155
rect 10609 29121 10643 29155
rect 10793 29121 10827 29155
rect 10885 29121 10919 29155
rect 12734 29121 12768 29155
rect 37381 29121 37415 29155
rect 39221 29121 39255 29155
rect 39405 29121 39439 29155
rect 39497 29121 39531 29155
rect 40233 29121 40267 29155
rect 44189 29121 44223 29155
rect 46673 29121 46707 29155
rect 49157 29121 49191 29155
rect 49893 29121 49927 29155
rect 51273 29121 51307 29155
rect 51457 29121 51491 29155
rect 51641 29121 51675 29155
rect 51825 29121 51859 29155
rect 53573 29121 53607 29155
rect 53757 29121 53791 29155
rect 55137 29121 55171 29155
rect 55781 29121 55815 29155
rect 56149 29121 56183 29155
rect 56241 29121 56275 29155
rect 56333 29121 56367 29155
rect 56517 29121 56551 29155
rect 56977 29121 57011 29155
rect 57161 29121 57195 29155
rect 57253 29121 57287 29155
rect 57437 29121 57471 29155
rect 58173 29121 58207 29155
rect 4445 29053 4479 29087
rect 10425 29053 10459 29087
rect 13001 29053 13035 29087
rect 37657 29053 37691 29087
rect 38301 29053 38335 29087
rect 39037 29053 39071 29087
rect 42257 29053 42291 29087
rect 42993 29053 43027 29087
rect 46765 29053 46799 29087
rect 48145 29053 48179 29087
rect 48421 29053 48455 29087
rect 49341 29053 49375 29087
rect 51733 29053 51767 29087
rect 52193 29053 52227 29087
rect 54861 29053 54895 29087
rect 55965 29053 55999 29087
rect 58265 29053 58299 29087
rect 6745 28985 6779 29019
rect 9045 28985 9079 29019
rect 11161 28985 11195 29019
rect 37473 28985 37507 29019
rect 37565 28985 37599 29019
rect 39405 28985 39439 29019
rect 39589 28985 39623 29019
rect 44097 28985 44131 29019
rect 52561 28985 52595 29019
rect 56425 28985 56459 29019
rect 57069 28985 57103 29019
rect 3893 28917 3927 28951
rect 4261 28917 4295 28951
rect 13369 28917 13403 28951
rect 38485 28917 38519 28951
rect 40496 28917 40530 28951
rect 42441 28917 42475 28951
rect 46029 28917 46063 28951
rect 47409 28917 47443 28951
rect 51181 28917 51215 28951
rect 53665 28917 53699 28951
rect 55045 28917 55079 28951
rect 3985 28713 4019 28747
rect 4813 28713 4847 28747
rect 5917 28713 5951 28747
rect 6469 28713 6503 28747
rect 9965 28713 9999 28747
rect 10609 28713 10643 28747
rect 11253 28713 11287 28747
rect 11621 28713 11655 28747
rect 36553 28713 36587 28747
rect 38669 28713 38703 28747
rect 40785 28713 40819 28747
rect 42809 28713 42843 28747
rect 44741 28713 44775 28747
rect 45569 28713 45603 28747
rect 48605 28713 48639 28747
rect 48881 28713 48915 28747
rect 49249 28713 49283 28747
rect 51549 28713 51583 28747
rect 52009 28713 52043 28747
rect 57161 28713 57195 28747
rect 57529 28713 57563 28747
rect 4261 28645 4295 28679
rect 6561 28645 6595 28679
rect 39405 28645 39439 28679
rect 41797 28645 41831 28679
rect 49525 28645 49559 28679
rect 49709 28645 49743 28679
rect 3341 28577 3375 28611
rect 7941 28577 7975 28611
rect 36737 28577 36771 28611
rect 37013 28577 37047 28611
rect 41705 28577 41739 28611
rect 42257 28577 42291 28611
rect 42441 28577 42475 28611
rect 45661 28577 45695 28611
rect 47409 28577 47443 28611
rect 47961 28577 47995 28611
rect 50169 28577 50203 28611
rect 52285 28577 52319 28611
rect 57437 28577 57471 28611
rect 57989 28577 58023 28611
rect 3249 28509 3283 28543
rect 3433 28509 3467 28543
rect 3893 28509 3927 28543
rect 4169 28509 4203 28543
rect 4353 28509 4387 28543
rect 4537 28509 4571 28543
rect 5825 28509 5859 28543
rect 6009 28509 6043 28543
rect 7674 28509 7708 28543
rect 9873 28509 9907 28543
rect 10057 28509 10091 28543
rect 10425 28509 10459 28543
rect 11253 28509 11287 28543
rect 11345 28509 11379 28543
rect 12909 28509 12943 28543
rect 38577 28509 38611 28543
rect 38761 28509 38795 28543
rect 40969 28509 41003 28543
rect 41061 28509 41095 28543
rect 42993 28509 43027 28543
rect 45109 28509 45143 28543
rect 45201 28509 45235 28543
rect 45385 28509 45419 28543
rect 49157 28509 49191 28543
rect 49617 28509 49651 28543
rect 49985 28509 50019 28543
rect 50629 28509 50663 28543
rect 51549 28509 51583 28543
rect 51641 28509 51675 28543
rect 51825 28509 51859 28543
rect 51917 28509 51951 28543
rect 52101 28509 52135 28543
rect 52377 28509 52411 28543
rect 53205 28509 53239 28543
rect 53389 28509 53423 28543
rect 57621 28509 57655 28543
rect 57713 28509 57747 28543
rect 57897 28509 57931 28543
rect 58081 28509 58115 28543
rect 58357 28509 58391 28543
rect 4813 28441 4847 28475
rect 6101 28441 6135 28475
rect 6285 28441 6319 28475
rect 10241 28441 10275 28475
rect 39037 28441 39071 28475
rect 43269 28441 43303 28475
rect 45937 28441 45971 28475
rect 48865 28441 48899 28475
rect 49065 28441 49099 28475
rect 49709 28441 49743 28475
rect 49893 28441 49927 28475
rect 58265 28441 58299 28475
rect 4629 28373 4663 28407
rect 5181 28373 5215 28407
rect 13001 28373 13035 28407
rect 38485 28373 38519 28407
rect 42165 28373 42199 28407
rect 48697 28373 48731 28407
rect 50445 28373 50479 28407
rect 50537 28373 50571 28407
rect 53297 28373 53331 28407
rect 3985 28169 4019 28203
rect 4905 28169 4939 28203
rect 8033 28169 8067 28203
rect 9045 28169 9079 28203
rect 9137 28169 9171 28203
rect 10241 28169 10275 28203
rect 10793 28169 10827 28203
rect 39129 28169 39163 28203
rect 41245 28169 41279 28203
rect 43361 28169 43395 28203
rect 43637 28169 43671 28203
rect 45293 28169 45327 28203
rect 49709 28169 49743 28203
rect 55689 28169 55723 28203
rect 57897 28169 57931 28203
rect 8585 28101 8619 28135
rect 39037 28101 39071 28135
rect 40601 28101 40635 28135
rect 46857 28101 46891 28135
rect 47317 28101 47351 28135
rect 49525 28101 49559 28135
rect 2697 28033 2731 28067
rect 3893 28033 3927 28067
rect 4077 28033 4111 28067
rect 4445 28033 4479 28067
rect 4629 28033 4663 28067
rect 8217 28033 8251 28067
rect 8493 28033 8527 28067
rect 8861 28033 8895 28067
rect 9321 28033 9355 28067
rect 9597 28033 9631 28067
rect 12633 28033 12667 28067
rect 38117 28033 38151 28067
rect 38301 28033 38335 28067
rect 38485 28033 38519 28067
rect 39865 28033 39899 28067
rect 40049 28033 40083 28067
rect 40141 28033 40175 28067
rect 40417 28033 40451 28067
rect 40785 28033 40819 28067
rect 40877 28033 40911 28067
rect 41153 28033 41187 28067
rect 41337 28033 41371 28067
rect 41981 28033 42015 28067
rect 42257 28033 42291 28067
rect 43269 28033 43303 28067
rect 43453 28033 43487 28067
rect 43729 28033 43763 28067
rect 47225 28033 47259 28067
rect 47409 28033 47443 28067
rect 47869 28033 47903 28067
rect 48513 28033 48547 28067
rect 49157 28033 49191 28067
rect 49341 28033 49375 28067
rect 49617 28033 49651 28067
rect 49801 28033 49835 28067
rect 50169 28033 50203 28067
rect 52377 28033 52411 28067
rect 52561 28033 52595 28067
rect 52745 28033 52779 28067
rect 53481 28033 53515 28067
rect 53748 28033 53782 28067
rect 55965 28033 55999 28067
rect 56149 28033 56183 28067
rect 56416 28033 56450 28067
rect 1593 27965 1627 27999
rect 3433 27965 3467 27999
rect 8401 27965 8435 27999
rect 8677 27965 8711 27999
rect 9413 27965 9447 27999
rect 12909 27965 12943 27999
rect 39681 27965 39715 27999
rect 41889 27965 41923 27999
rect 44005 27965 44039 27999
rect 44649 27965 44683 27999
rect 45385 27965 45419 27999
rect 47133 27965 47167 27999
rect 48145 27965 48179 27999
rect 48421 27965 48455 27999
rect 52285 27965 52319 27999
rect 52469 27965 52503 27999
rect 53297 27965 53331 27999
rect 54953 27965 54987 27999
rect 55689 27965 55723 27999
rect 58449 27965 58483 27999
rect 13461 27897 13495 27931
rect 47593 27897 47627 27931
rect 54861 27897 54895 27931
rect 57529 27897 57563 27931
rect 2881 27829 2915 27863
rect 4537 27829 4571 27863
rect 5365 27829 5399 27863
rect 6837 27829 6871 27863
rect 7389 27829 7423 27863
rect 8493 27829 8527 27863
rect 8861 27829 8895 27863
rect 9597 27829 9631 27863
rect 38209 27829 38243 27863
rect 40325 27829 40359 27863
rect 40601 27829 40635 27863
rect 51641 27829 51675 27863
rect 55597 27829 55631 27863
rect 55873 27829 55907 27863
rect 3341 27625 3375 27659
rect 10977 27625 11011 27659
rect 43545 27625 43579 27659
rect 44005 27625 44039 27659
rect 47317 27625 47351 27659
rect 47685 27625 47719 27659
rect 52561 27625 52595 27659
rect 53205 27625 53239 27659
rect 55413 27625 55447 27659
rect 56425 27625 56459 27659
rect 58357 27625 58391 27659
rect 4261 27557 4295 27591
rect 13461 27557 13495 27591
rect 15485 27557 15519 27591
rect 38117 27557 38151 27591
rect 38945 27557 38979 27591
rect 45109 27557 45143 27591
rect 50629 27557 50663 27591
rect 53849 27557 53883 27591
rect 56517 27557 56551 27591
rect 57989 27557 58023 27591
rect 3157 27489 3191 27523
rect 7297 27489 7331 27523
rect 9781 27489 9815 27523
rect 38209 27489 38243 27523
rect 40049 27489 40083 27523
rect 40141 27489 40175 27523
rect 40417 27489 40451 27523
rect 53757 27489 53791 27523
rect 54125 27489 54159 27523
rect 54769 27489 54803 27523
rect 54953 27489 54987 27523
rect 56333 27489 56367 27523
rect 56701 27489 56735 27523
rect 57345 27489 57379 27523
rect 57529 27489 57563 27523
rect 3249 27421 3283 27455
rect 3433 27421 3467 27455
rect 3985 27421 4019 27455
rect 5466 27421 5500 27455
rect 5733 27421 5767 27455
rect 6469 27421 6503 27455
rect 7021 27421 7055 27455
rect 7481 27421 7515 27455
rect 10057 27421 10091 27455
rect 10701 27421 10735 27455
rect 12357 27421 12391 27455
rect 12633 27421 12667 27455
rect 12817 27421 12851 27455
rect 13001 27421 13035 27455
rect 13185 27421 13219 27455
rect 14105 27421 14139 27455
rect 14361 27421 14395 27455
rect 24593 27421 24627 27455
rect 25789 27421 25823 27455
rect 37933 27421 37967 27455
rect 38025 27421 38059 27455
rect 38669 27421 38703 27455
rect 38761 27421 38795 27455
rect 39957 27421 39991 27455
rect 40325 27421 40359 27455
rect 43453 27421 43487 27455
rect 43645 27423 43679 27457
rect 44465 27421 44499 27455
rect 45017 27421 45051 27455
rect 45753 27421 45787 27455
rect 45937 27421 45971 27455
rect 46121 27421 46155 27455
rect 46489 27421 46523 27455
rect 47961 27421 47995 27455
rect 48237 27421 48271 27455
rect 48329 27421 48363 27455
rect 48513 27421 48547 27455
rect 49801 27421 49835 27455
rect 49893 27421 49927 27455
rect 50353 27421 50387 27455
rect 50997 27421 51031 27455
rect 51181 27421 51215 27455
rect 53113 27421 53147 27455
rect 53297 27421 53331 27455
rect 53941 27421 53975 27455
rect 54033 27421 54067 27455
rect 54861 27421 54895 27455
rect 55045 27421 55079 27455
rect 55321 27421 55355 27455
rect 55505 27421 55539 27455
rect 56609 27421 56643 27455
rect 57437 27421 57471 27455
rect 57621 27421 57655 27455
rect 57805 27421 57839 27455
rect 58081 27421 58115 27455
rect 58541 27421 58575 27455
rect 2881 27353 2915 27387
rect 4077 27353 4111 27387
rect 4261 27353 4295 27387
rect 6653 27353 6687 27387
rect 6837 27353 6871 27387
rect 7665 27353 7699 27387
rect 10425 27353 10459 27387
rect 12090 27353 12124 27387
rect 13093 27353 13127 27387
rect 25329 27353 25363 27387
rect 45845 27353 45879 27387
rect 48053 27353 48087 27387
rect 49617 27353 49651 27387
rect 50261 27353 50295 27387
rect 51448 27353 51482 27387
rect 1409 27285 1443 27319
rect 4353 27285 4387 27319
rect 6285 27285 6319 27319
rect 7205 27285 7239 27319
rect 8033 27285 8067 27319
rect 12449 27285 12483 27319
rect 13829 27285 13863 27319
rect 39221 27285 39255 27319
rect 39865 27285 39899 27319
rect 42165 27285 42199 27319
rect 42901 27285 42935 27319
rect 44741 27285 44775 27319
rect 48697 27285 48731 27319
rect 48973 27285 49007 27319
rect 58173 27285 58207 27319
rect 2697 27081 2731 27115
rect 3893 27081 3927 27115
rect 4629 27081 4663 27115
rect 8953 27081 8987 27115
rect 10609 27081 10643 27115
rect 11345 27081 11379 27115
rect 12817 27081 12851 27115
rect 38485 27081 38519 27115
rect 43085 27081 43119 27115
rect 46857 27081 46891 27115
rect 51457 27081 51491 27115
rect 54585 27081 54619 27115
rect 2789 27013 2823 27047
rect 4077 27013 4111 27047
rect 4813 27013 4847 27047
rect 6009 27013 6043 27047
rect 10333 27013 10367 27047
rect 11069 27013 11103 27047
rect 12081 27013 12115 27047
rect 39681 27013 39715 27047
rect 40509 27013 40543 27047
rect 43361 27013 43395 27047
rect 43453 27013 43487 27047
rect 43571 27013 43605 27047
rect 43821 27013 43855 27047
rect 44925 27013 44959 27047
rect 46213 27013 46247 27047
rect 2145 26945 2179 26979
rect 3065 26945 3099 26979
rect 3985 26945 4019 26979
rect 4169 26945 4203 26979
rect 4997 26945 5031 26979
rect 6193 26945 6227 26979
rect 6653 26945 6687 26979
rect 7021 26945 7055 26979
rect 7205 26945 7239 26979
rect 7297 26945 7331 26979
rect 7840 26945 7874 26979
rect 10149 26945 10183 26979
rect 10425 26945 10459 26979
rect 11161 26945 11195 26979
rect 11897 26945 11931 26979
rect 38669 26945 38703 26979
rect 38853 26945 38887 26979
rect 38945 26945 38979 26979
rect 39865 26945 39899 26979
rect 39957 26945 39991 26979
rect 40049 26945 40083 26979
rect 42441 26945 42475 26979
rect 42625 26945 42659 26979
rect 42809 26945 42843 26979
rect 42993 26945 43027 26979
rect 43269 26945 43303 26979
rect 44097 26945 44131 26979
rect 45753 26945 45787 26979
rect 45845 26945 45879 26979
rect 46305 26945 46339 26979
rect 46397 26945 46431 26979
rect 46581 26945 46615 26979
rect 47961 26945 47995 26979
rect 48053 26945 48087 26979
rect 48237 26945 48271 26979
rect 49433 26945 49467 26979
rect 50905 26945 50939 26979
rect 51733 26945 51767 26979
rect 53481 26945 53515 26979
rect 53665 26945 53699 26979
rect 56701 26945 56735 26979
rect 56885 26945 56919 26979
rect 57897 26945 57931 26979
rect 2789 26877 2823 26911
rect 3249 26877 3283 26911
rect 6377 26877 6411 26911
rect 7573 26877 7607 26911
rect 36921 26877 36955 26911
rect 40233 26877 40267 26911
rect 42901 26877 42935 26911
rect 43729 26877 43763 26911
rect 43821 26877 43855 26911
rect 49801 26877 49835 26911
rect 50169 26877 50203 26911
rect 51181 26877 51215 26911
rect 51457 26877 51491 26911
rect 56057 26877 56091 26911
rect 56793 26877 56827 26911
rect 57529 26877 57563 26911
rect 58541 26877 58575 26911
rect 7389 26809 7423 26843
rect 38393 26809 38427 26843
rect 44005 26809 44039 26843
rect 45937 26809 45971 26843
rect 46581 26809 46615 26843
rect 2973 26741 3007 26775
rect 5825 26741 5859 26775
rect 6469 26741 6503 26775
rect 6561 26741 6595 26775
rect 7113 26741 7147 26775
rect 9965 26741 9999 26775
rect 11713 26741 11747 26775
rect 12541 26741 12575 26775
rect 36277 26741 36311 26775
rect 37473 26741 37507 26775
rect 41981 26741 42015 26775
rect 42441 26741 42475 26775
rect 47225 26741 47259 26775
rect 48421 26741 48455 26775
rect 48789 26741 48823 26775
rect 50813 26741 50847 26775
rect 51641 26741 51675 26775
rect 53573 26741 53607 26775
rect 55413 26741 55447 26775
rect 56977 26741 57011 26775
rect 6745 26537 6779 26571
rect 7941 26537 7975 26571
rect 10057 26537 10091 26571
rect 35357 26537 35391 26571
rect 40141 26537 40175 26571
rect 42257 26537 42291 26571
rect 43085 26537 43119 26571
rect 46213 26537 46247 26571
rect 47869 26537 47903 26571
rect 48500 26537 48534 26571
rect 49985 26537 50019 26571
rect 51641 26537 51675 26571
rect 53757 26537 53791 26571
rect 53941 26537 53975 26571
rect 54585 26537 54619 26571
rect 54953 26537 54987 26571
rect 56701 26537 56735 26571
rect 58173 26537 58207 26571
rect 6377 26469 6411 26503
rect 12357 26469 12391 26503
rect 39129 26469 39163 26503
rect 39405 26469 39439 26503
rect 40509 26469 40543 26503
rect 41061 26469 41095 26503
rect 44833 26469 44867 26503
rect 8217 26401 8251 26435
rect 35449 26401 35483 26435
rect 37197 26401 37231 26435
rect 37289 26401 37323 26435
rect 41220 26401 41254 26435
rect 45385 26401 45419 26435
rect 48237 26401 48271 26435
rect 53389 26401 53423 26435
rect 55137 26401 55171 26435
rect 56793 26401 56827 26435
rect 2605 26333 2639 26367
rect 2881 26333 2915 26367
rect 3525 26333 3559 26367
rect 3801 26333 3835 26367
rect 3985 26333 4019 26367
rect 4629 26333 4663 26367
rect 4813 26333 4847 26367
rect 7665 26333 7699 26367
rect 10149 26333 10183 26367
rect 12173 26333 12207 26367
rect 13654 26333 13688 26367
rect 13921 26333 13955 26367
rect 38209 26333 38243 26367
rect 38485 26333 38519 26367
rect 38669 26333 38703 26367
rect 38853 26333 38887 26367
rect 40417 26333 40451 26367
rect 41705 26333 41739 26367
rect 42441 26333 42475 26367
rect 43177 26333 43211 26367
rect 43269 26333 43303 26367
rect 44557 26333 44591 26367
rect 44649 26333 44683 26367
rect 44833 26333 44867 26367
rect 45017 26333 45051 26367
rect 45201 26333 45235 26367
rect 45293 26333 45327 26367
rect 45489 26333 45523 26367
rect 46121 26333 46155 26367
rect 46305 26333 46339 26367
rect 46397 26333 46431 26367
rect 47225 26333 47259 26367
rect 47501 26333 47535 26367
rect 47777 26333 47811 26367
rect 52745 26333 52779 26367
rect 53757 26333 53791 26367
rect 53849 26333 53883 26367
rect 54125 26333 54159 26367
rect 54493 26333 54527 26367
rect 54677 26333 54711 26367
rect 54861 26333 54895 26367
rect 55321 26333 55355 26367
rect 58449 26333 58483 26367
rect 1593 26265 1627 26299
rect 7941 26265 7975 26299
rect 14289 26265 14323 26299
rect 35725 26265 35759 26299
rect 38025 26265 38059 26299
rect 39129 26265 39163 26299
rect 41429 26265 41463 26299
rect 42993 26265 43027 26299
rect 45109 26265 45143 26299
rect 46489 26265 46523 26299
rect 50169 26265 50203 26299
rect 53481 26265 53515 26299
rect 53665 26265 53699 26299
rect 54217 26265 54251 26299
rect 54401 26265 54435 26299
rect 55137 26265 55171 26299
rect 55566 26265 55600 26299
rect 57060 26265 57094 26299
rect 3893 26197 3927 26231
rect 4813 26197 4847 26231
rect 7757 26197 7791 26231
rect 12541 26197 12575 26231
rect 37933 26197 37967 26231
rect 38945 26197 38979 26231
rect 41337 26197 41371 26231
rect 42073 26197 42107 26231
rect 47317 26197 47351 26231
rect 47685 26197 47719 26231
rect 54309 26197 54343 26231
rect 58265 26197 58299 26231
rect 1409 25993 1443 26027
rect 5457 25993 5491 26027
rect 7389 25993 7423 26027
rect 8309 25993 8343 26027
rect 10057 25993 10091 26027
rect 10517 25993 10551 26027
rect 11529 25993 11563 26027
rect 11713 25993 11747 26027
rect 12541 25993 12575 26027
rect 35725 25993 35759 26027
rect 37289 25993 37323 26027
rect 37841 25993 37875 26027
rect 39129 25993 39163 26027
rect 46949 25993 46983 26027
rect 47869 25993 47903 26027
rect 52469 25993 52503 26027
rect 54677 25993 54711 26027
rect 55321 25993 55355 26027
rect 56977 25993 57011 26027
rect 7205 25925 7239 25959
rect 11805 25925 11839 25959
rect 12173 25925 12207 25959
rect 36829 25925 36863 25959
rect 45385 25925 45419 25959
rect 47777 25925 47811 25959
rect 48237 25925 48271 25959
rect 50905 25925 50939 25959
rect 12403 25891 12437 25925
rect 3893 25857 3927 25891
rect 4344 25857 4378 25891
rect 7481 25857 7515 25891
rect 8493 25857 8527 25891
rect 8585 25857 8619 25891
rect 8769 25857 8803 25891
rect 9321 25857 9355 25891
rect 9505 25857 9539 25891
rect 9689 25857 9723 25891
rect 10333 25857 10367 25891
rect 10517 25857 10551 25891
rect 10701 25857 10735 25891
rect 10793 25857 10827 25891
rect 11161 25857 11195 25891
rect 11345 25857 11379 25891
rect 11897 25857 11931 25891
rect 29837 25857 29871 25891
rect 35449 25857 35483 25891
rect 35633 25857 35667 25891
rect 36461 25857 36495 25891
rect 36645 25857 36679 25891
rect 36921 25857 36955 25891
rect 37289 25857 37323 25891
rect 37473 25857 37507 25891
rect 37749 25857 37783 25891
rect 37933 25857 37967 25891
rect 39221 25863 39255 25897
rect 39773 25857 39807 25891
rect 39957 25857 39991 25891
rect 45293 25857 45327 25891
rect 45477 25857 45511 25891
rect 46765 25857 46799 25891
rect 46949 25857 46983 25891
rect 48053 25857 48087 25891
rect 48513 25857 48547 25891
rect 51089 25857 51123 25891
rect 51356 25857 51390 25891
rect 53481 25857 53515 25891
rect 53665 25857 53699 25891
rect 54769 25857 54803 25891
rect 56057 25857 56091 25891
rect 56241 25857 56275 25891
rect 57161 25857 57195 25891
rect 57253 25857 57287 25891
rect 57897 25857 57931 25891
rect 58173 25857 58207 25891
rect 2881 25789 2915 25823
rect 3157 25789 3191 25823
rect 4077 25789 4111 25823
rect 9781 25789 9815 25823
rect 11253 25789 11287 25823
rect 35541 25789 35575 25823
rect 36277 25789 36311 25823
rect 48145 25789 48179 25823
rect 50169 25789 50203 25823
rect 53389 25789 53423 25823
rect 53573 25789 53607 25823
rect 55965 25789 55999 25823
rect 56149 25789 56183 25823
rect 56977 25789 57011 25823
rect 12081 25721 12115 25755
rect 31309 25721 31343 25755
rect 46305 25721 46339 25755
rect 48973 25721 49007 25755
rect 58265 25721 58299 25755
rect 3249 25653 3283 25687
rect 7205 25653 7239 25687
rect 8769 25653 8803 25687
rect 9137 25653 9171 25687
rect 9321 25653 9355 25687
rect 9873 25653 9907 25687
rect 12357 25653 12391 25687
rect 38209 25653 38243 25687
rect 39957 25653 39991 25687
rect 41337 25653 41371 25687
rect 41797 25653 41831 25687
rect 49801 25653 49835 25687
rect 52745 25653 52779 25687
rect 58081 25653 58115 25687
rect 3433 25449 3467 25483
rect 3893 25449 3927 25483
rect 4537 25449 4571 25483
rect 5733 25449 5767 25483
rect 7481 25449 7515 25483
rect 8769 25449 8803 25483
rect 10149 25449 10183 25483
rect 11805 25449 11839 25483
rect 12541 25449 12575 25483
rect 13093 25449 13127 25483
rect 13829 25449 13863 25483
rect 37105 25449 37139 25483
rect 38025 25449 38059 25483
rect 39681 25449 39715 25483
rect 40969 25449 41003 25483
rect 41429 25449 41463 25483
rect 44649 25449 44683 25483
rect 48053 25449 48087 25483
rect 48513 25449 48547 25483
rect 51365 25449 51399 25483
rect 51457 25449 51491 25483
rect 2421 25381 2455 25415
rect 5917 25381 5951 25415
rect 40325 25381 40359 25415
rect 40785 25381 40819 25415
rect 44281 25381 44315 25415
rect 58265 25381 58299 25415
rect 2605 25313 2639 25347
rect 5549 25313 5583 25347
rect 8585 25313 8619 25347
rect 9965 25313 9999 25347
rect 42533 25313 42567 25347
rect 45661 25313 45695 25347
rect 46489 25313 46523 25347
rect 46857 25313 46891 25347
rect 46949 25313 46983 25347
rect 51273 25313 51307 25347
rect 53297 25313 53331 25347
rect 53849 25313 53883 25347
rect 57437 25313 57471 25347
rect 57713 25313 57747 25347
rect 2329 25245 2363 25279
rect 2789 25245 2823 25279
rect 3801 25245 3835 25279
rect 4077 25245 4111 25279
rect 4261 25245 4295 25279
rect 4813 25245 4847 25279
rect 5273 25245 5307 25279
rect 5825 25245 5859 25279
rect 7041 25245 7075 25279
rect 7297 25245 7331 25279
rect 7389 25245 7423 25279
rect 7573 25245 7607 25279
rect 8493 25245 8527 25279
rect 9321 25245 9355 25279
rect 10149 25245 10183 25279
rect 11897 25245 11931 25279
rect 11989 25245 12023 25279
rect 12173 25245 12207 25279
rect 12909 25245 12943 25279
rect 13093 25245 13127 25279
rect 13369 25245 13403 25279
rect 36829 25245 36863 25279
rect 37013 25245 37047 25279
rect 37289 25245 37323 25279
rect 37473 25245 37507 25279
rect 37565 25245 37599 25279
rect 37657 25245 37691 25279
rect 37841 25245 37875 25279
rect 37933 25245 37967 25279
rect 38761 25245 38795 25279
rect 38945 25245 38979 25279
rect 39313 25245 39347 25279
rect 39497 25245 39531 25279
rect 39681 25245 39715 25279
rect 40049 25245 40083 25279
rect 41705 25245 41739 25279
rect 41889 25245 41923 25279
rect 42165 25245 42199 25279
rect 45753 25245 45787 25279
rect 45937 25245 45971 25279
rect 46029 25245 46063 25279
rect 46121 25245 46155 25279
rect 46673 25245 46707 25279
rect 46765 25245 46799 25279
rect 47133 25245 47167 25279
rect 47317 25245 47351 25279
rect 47961 25245 47995 25279
rect 49249 25245 49283 25279
rect 51549 25245 51583 25279
rect 53205 25245 53239 25279
rect 53389 25245 53423 25279
rect 53481 25245 53515 25279
rect 53665 25245 53699 25279
rect 53757 25245 53791 25279
rect 53941 25245 53975 25279
rect 54217 25245 54251 25279
rect 54401 25245 54435 25279
rect 54585 25245 54619 25279
rect 54769 25245 54803 25279
rect 55965 25245 55999 25279
rect 57161 25245 57195 25279
rect 57253 25245 57287 25279
rect 57621 25245 57655 25279
rect 57805 25245 57839 25279
rect 57897 25245 57931 25279
rect 58173 25245 58207 25279
rect 2605 25177 2639 25211
rect 4537 25177 4571 25211
rect 5089 25177 5123 25211
rect 8769 25177 8803 25211
rect 9873 25177 9907 25211
rect 12081 25177 12115 25211
rect 36921 25177 36955 25211
rect 37749 25177 37783 25211
rect 39957 25177 39991 25211
rect 41153 25177 41187 25211
rect 41245 25177 41279 25211
rect 41461 25177 41495 25211
rect 41797 25177 41831 25211
rect 42809 25177 42843 25211
rect 54677 25177 54711 25211
rect 4077 25109 4111 25143
rect 4721 25109 4755 25143
rect 4905 25109 4939 25143
rect 5549 25109 5583 25143
rect 8309 25109 8343 25143
rect 9045 25109 9079 25143
rect 10333 25109 10367 25143
rect 13277 25109 13311 25143
rect 13461 25109 13495 25143
rect 38945 25109 38979 25143
rect 40953 25109 40987 25143
rect 41613 25109 41647 25143
rect 45017 25109 45051 25143
rect 46397 25109 46431 25143
rect 47225 25109 47259 25143
rect 48697 25109 48731 25143
rect 53021 25109 53055 25143
rect 53481 25109 53515 25143
rect 54309 25109 54343 25143
rect 55321 25109 55355 25143
rect 57437 25109 57471 25143
rect 58081 25109 58115 25143
rect 4077 24905 4111 24939
rect 5917 24905 5951 24939
rect 11989 24905 12023 24939
rect 12633 24905 12667 24939
rect 14565 24905 14599 24939
rect 38393 24905 38427 24939
rect 38945 24905 38979 24939
rect 40509 24905 40543 24939
rect 41613 24905 41647 24939
rect 42717 24905 42751 24939
rect 42809 24905 42843 24939
rect 46765 24905 46799 24939
rect 48605 24905 48639 24939
rect 53757 24905 53791 24939
rect 12173 24837 12207 24871
rect 13452 24837 13486 24871
rect 45937 24837 45971 24871
rect 46933 24837 46967 24871
rect 47133 24837 47167 24871
rect 47317 24837 47351 24871
rect 54953 24837 54987 24871
rect 2697 24769 2731 24803
rect 12265 24769 12299 24803
rect 12541 24769 12575 24803
rect 13185 24769 13219 24803
rect 37473 24769 37507 24803
rect 37657 24769 37691 24803
rect 38209 24769 38243 24803
rect 38485 24769 38519 24803
rect 38761 24769 38795 24803
rect 39037 24769 39071 24803
rect 39773 24769 39807 24803
rect 39957 24769 39991 24803
rect 40417 24769 40451 24803
rect 40693 24769 40727 24803
rect 40877 24769 40911 24803
rect 41245 24769 41279 24803
rect 41337 24769 41371 24803
rect 41521 24769 41555 24803
rect 41705 24769 41739 24803
rect 43729 24769 43763 24803
rect 43821 24769 43855 24803
rect 44005 24769 44039 24803
rect 44097 24769 44131 24803
rect 44189 24769 44223 24803
rect 44465 24769 44499 24803
rect 44557 24769 44591 24803
rect 44649 24769 44683 24803
rect 45293 24769 45327 24803
rect 45477 24769 45511 24803
rect 46121 24769 46155 24803
rect 46397 24769 46431 24803
rect 46489 24769 46523 24803
rect 46673 24769 46707 24803
rect 47225 24769 47259 24803
rect 47409 24769 47443 24803
rect 47961 24769 47995 24803
rect 48053 24769 48087 24803
rect 48237 24769 48271 24803
rect 48329 24769 48363 24803
rect 48697 24769 48731 24803
rect 50905 24769 50939 24803
rect 51365 24769 51399 24803
rect 51641 24769 51675 24803
rect 51825 24769 51859 24803
rect 51917 24769 51951 24803
rect 52101 24769 52135 24803
rect 52745 24769 52779 24803
rect 52929 24769 52963 24803
rect 53021 24769 53055 24803
rect 53205 24769 53239 24803
rect 53297 24769 53331 24803
rect 53481 24769 53515 24803
rect 54677 24769 54711 24803
rect 55045 24769 55079 24803
rect 55301 24769 55335 24803
rect 56977 24769 57011 24803
rect 57161 24769 57195 24803
rect 58081 24769 58115 24803
rect 58173 24769 58207 24803
rect 1593 24701 1627 24735
rect 3709 24701 3743 24735
rect 37749 24701 37783 24735
rect 39865 24701 39899 24735
rect 43453 24701 43487 24735
rect 43545 24701 43579 24735
rect 48145 24701 48179 24735
rect 48605 24701 48639 24735
rect 48973 24701 49007 24735
rect 52837 24701 52871 24735
rect 54769 24701 54803 24735
rect 54953 24701 54987 24735
rect 13001 24633 13035 24667
rect 38669 24633 38703 24667
rect 40877 24633 40911 24667
rect 44327 24633 44361 24667
rect 45845 24633 45879 24667
rect 47869 24633 47903 24667
rect 52009 24633 52043 24667
rect 56793 24633 56827 24667
rect 58265 24633 58299 24667
rect 3157 24565 3191 24599
rect 10149 24565 10183 24599
rect 37013 24565 37047 24599
rect 37289 24565 37323 24599
rect 38025 24565 38059 24599
rect 42073 24565 42107 24599
rect 45477 24565 45511 24599
rect 46949 24565 46983 24599
rect 48421 24565 48455 24599
rect 50445 24565 50479 24599
rect 51733 24565 51767 24599
rect 53113 24565 53147 24599
rect 53389 24565 53423 24599
rect 56425 24565 56459 24599
rect 57069 24565 57103 24599
rect 57897 24565 57931 24599
rect 3341 24361 3375 24395
rect 3433 24361 3467 24395
rect 7941 24361 7975 24395
rect 11897 24361 11931 24395
rect 14289 24361 14323 24395
rect 37749 24361 37783 24395
rect 39589 24361 39623 24395
rect 44557 24361 44591 24395
rect 47133 24361 47167 24395
rect 48605 24361 48639 24395
rect 49433 24361 49467 24395
rect 4905 24293 4939 24327
rect 7665 24293 7699 24327
rect 8493 24293 8527 24327
rect 10425 24293 10459 24327
rect 13829 24293 13863 24327
rect 43729 24293 43763 24327
rect 44373 24293 44407 24327
rect 49709 24293 49743 24327
rect 56149 24293 56183 24327
rect 2881 24225 2915 24259
rect 3157 24225 3191 24259
rect 3525 24225 3559 24259
rect 3801 24225 3835 24259
rect 6745 24225 6779 24259
rect 9781 24225 9815 24259
rect 35081 24225 35115 24259
rect 35173 24225 35207 24259
rect 36921 24225 36955 24259
rect 38301 24225 38335 24259
rect 43085 24225 43119 24259
rect 47041 24225 47075 24259
rect 47317 24225 47351 24259
rect 48789 24225 48823 24259
rect 55965 24225 55999 24259
rect 3249 24157 3283 24191
rect 4353 24157 4387 24191
rect 4629 24157 4663 24191
rect 4721 24157 4755 24191
rect 6929 24157 6963 24191
rect 7021 24157 7055 24191
rect 7389 24157 7423 24191
rect 7481 24157 7515 24191
rect 8217 24157 8251 24191
rect 8309 24157 8343 24191
rect 9965 24157 9999 24191
rect 10057 24157 10091 24191
rect 10149 24157 10183 24191
rect 10517 24157 10551 24191
rect 10773 24157 10807 24191
rect 12449 24157 12483 24191
rect 12541 24157 12575 24191
rect 12725 24157 12759 24191
rect 13461 24157 13495 24191
rect 13553 24157 13587 24191
rect 13829 24157 13863 24191
rect 37565 24157 37599 24191
rect 39129 24157 39163 24191
rect 39221 24157 39255 24191
rect 39405 24157 39439 24191
rect 39497 24157 39531 24191
rect 39681 24157 39715 24191
rect 39865 24157 39899 24191
rect 41337 24157 41371 24191
rect 43269 24157 43303 24191
rect 44649 24157 44683 24191
rect 45017 24157 45051 24191
rect 45293 24157 45327 24191
rect 45477 24157 45511 24191
rect 47133 24157 47167 24191
rect 47225 24157 47259 24191
rect 47409 24157 47443 24191
rect 48513 24157 48547 24191
rect 48697 24157 48731 24191
rect 49617 24157 49651 24191
rect 50813 24157 50847 24191
rect 51273 24157 51307 24191
rect 51457 24157 51491 24191
rect 51549 24157 51583 24191
rect 51733 24157 51767 24191
rect 52837 24157 52871 24191
rect 53021 24157 53055 24191
rect 54861 24157 54895 24191
rect 56057 24157 56091 24191
rect 56241 24157 56275 24191
rect 56885 24157 56919 24191
rect 57069 24157 57103 24191
rect 57897 24157 57931 24191
rect 58173 24157 58207 24191
rect 4905 24089 4939 24123
rect 7665 24089 7699 24123
rect 8493 24089 8527 24123
rect 10425 24089 10459 24123
rect 12173 24089 12207 24123
rect 13185 24089 13219 24123
rect 35449 24089 35483 24123
rect 39957 24089 39991 24123
rect 41613 24089 41647 24123
rect 44005 24089 44039 24123
rect 44189 24089 44223 24123
rect 45109 24089 45143 24123
rect 55321 24089 55355 24123
rect 58265 24089 58299 24123
rect 1409 24021 1443 24055
rect 6745 24021 6779 24055
rect 9781 24021 9815 24055
rect 10241 24021 10275 24055
rect 12725 24021 12759 24055
rect 13645 24021 13679 24055
rect 37013 24021 37047 24055
rect 38485 24021 38519 24055
rect 39313 24021 39347 24055
rect 43453 24021 43487 24055
rect 46765 24021 46799 24055
rect 47777 24021 47811 24055
rect 48145 24021 48179 24055
rect 50629 24021 50663 24055
rect 51365 24021 51399 24055
rect 51733 24021 51767 24055
rect 52929 24021 52963 24055
rect 54769 24021 54803 24055
rect 56885 24021 56919 24055
rect 57989 24021 58023 24055
rect 3985 23817 4019 23851
rect 8033 23817 8067 23851
rect 10149 23817 10183 23851
rect 10517 23817 10551 23851
rect 12909 23817 12943 23851
rect 35725 23817 35759 23851
rect 38485 23817 38519 23851
rect 39589 23817 39623 23851
rect 42441 23817 42475 23851
rect 44097 23817 44131 23851
rect 53849 23817 53883 23851
rect 4169 23749 4203 23783
rect 5466 23749 5500 23783
rect 7512 23749 7546 23783
rect 8392 23749 8426 23783
rect 14114 23749 14148 23783
rect 36461 23749 36495 23783
rect 37657 23749 37691 23783
rect 38853 23749 38887 23783
rect 54769 23749 54803 23783
rect 2697 23681 2731 23715
rect 3341 23681 3375 23715
rect 3801 23681 3835 23715
rect 3985 23681 4019 23715
rect 4077 23681 4111 23715
rect 4261 23681 4295 23715
rect 5733 23681 5767 23715
rect 7757 23681 7791 23715
rect 7849 23681 7883 23715
rect 8033 23681 8067 23715
rect 10149 23681 10183 23715
rect 10333 23681 10367 23715
rect 10425 23681 10459 23715
rect 12265 23681 12299 23715
rect 12725 23681 12759 23715
rect 12909 23681 12943 23715
rect 14381 23681 14415 23715
rect 36369 23681 36403 23715
rect 36737 23681 36771 23715
rect 36829 23681 36863 23715
rect 37013 23681 37047 23715
rect 37381 23681 37415 23715
rect 38301 23681 38335 23715
rect 38485 23681 38519 23715
rect 38669 23681 38703 23715
rect 39589 23681 39623 23715
rect 39773 23681 39807 23715
rect 43361 23681 43395 23715
rect 43729 23681 43763 23715
rect 43913 23681 43947 23715
rect 44189 23681 44223 23715
rect 44281 23681 44315 23715
rect 47961 23681 47995 23715
rect 48145 23681 48179 23715
rect 49985 23681 50019 23715
rect 50169 23681 50203 23715
rect 50261 23681 50295 23715
rect 50439 23681 50473 23715
rect 50537 23681 50571 23715
rect 50721 23681 50755 23715
rect 52745 23681 52779 23715
rect 52929 23681 52963 23715
rect 54033 23681 54067 23715
rect 54217 23681 54251 23715
rect 54309 23681 54343 23715
rect 54401 23681 54435 23715
rect 54585 23681 54619 23715
rect 54677 23681 54711 23715
rect 54861 23681 54895 23715
rect 54953 23681 54987 23715
rect 55137 23681 55171 23715
rect 56508 23681 56542 23715
rect 8125 23613 8159 23647
rect 11989 23613 12023 23647
rect 36461 23613 36495 23647
rect 37657 23613 37691 23647
rect 39405 23613 39439 23647
rect 41337 23613 41371 23647
rect 41521 23613 41555 23647
rect 42165 23613 42199 23647
rect 43085 23613 43119 23647
rect 43177 23613 43211 23647
rect 43637 23613 43671 23647
rect 44373 23613 44407 23647
rect 46581 23613 46615 23647
rect 49617 23613 49651 23647
rect 49893 23613 49927 23647
rect 50077 23613 50111 23647
rect 52837 23613 52871 23647
rect 55045 23613 55079 23647
rect 56241 23613 56275 23647
rect 58449 23613 58483 23647
rect 12173 23545 12207 23579
rect 13001 23545 13035 23579
rect 36645 23545 36679 23579
rect 37473 23545 37507 23579
rect 41061 23545 41095 23579
rect 54309 23545 54343 23579
rect 57621 23545 57655 23579
rect 4353 23477 4387 23511
rect 6377 23477 6411 23511
rect 9505 23477 9539 23511
rect 10977 23477 11011 23511
rect 12081 23477 12115 23511
rect 12541 23477 12575 23511
rect 36921 23477 36955 23511
rect 37749 23477 37783 23511
rect 40877 23477 40911 23511
rect 43545 23477 43579 23511
rect 45937 23477 45971 23511
rect 48053 23477 48087 23511
rect 50261 23477 50295 23511
rect 50629 23477 50663 23511
rect 54493 23477 54527 23511
rect 57897 23477 57931 23511
rect 4721 23273 4755 23307
rect 7297 23273 7331 23307
rect 8217 23273 8251 23307
rect 12357 23273 12391 23307
rect 39221 23273 39255 23307
rect 42717 23273 42751 23307
rect 47317 23273 47351 23307
rect 48605 23273 48639 23307
rect 52837 23273 52871 23307
rect 56517 23273 56551 23307
rect 56609 23273 56643 23307
rect 58357 23273 58391 23307
rect 3893 23205 3927 23239
rect 48789 23205 48823 23239
rect 48973 23205 49007 23239
rect 51181 23205 51215 23239
rect 6653 23137 6687 23171
rect 37381 23137 37415 23171
rect 37473 23137 37507 23171
rect 46765 23137 46799 23171
rect 48513 23137 48547 23171
rect 49157 23137 49191 23171
rect 49249 23137 49283 23171
rect 49893 23137 49927 23171
rect 52561 23137 52595 23171
rect 55689 23137 55723 23171
rect 56425 23137 56459 23171
rect 56793 23137 56827 23171
rect 57805 23137 57839 23171
rect 58081 23137 58115 23171
rect 2605 23069 2639 23103
rect 2881 23069 2915 23103
rect 3801 23069 3835 23103
rect 3985 23069 4019 23103
rect 4629 23069 4663 23103
rect 4813 23069 4847 23103
rect 6837 23069 6871 23103
rect 6929 23069 6963 23103
rect 7205 23069 7239 23103
rect 7389 23069 7423 23103
rect 8309 23069 8343 23103
rect 8585 23069 8619 23103
rect 9965 23069 9999 23103
rect 10149 23069 10183 23103
rect 39497 23069 39531 23103
rect 39589 23069 39623 23103
rect 39865 23069 39899 23103
rect 45017 23069 45051 23103
rect 46857 23069 46891 23103
rect 47777 23069 47811 23103
rect 48053 23069 48087 23103
rect 48237 23069 48271 23103
rect 48881 23069 48915 23103
rect 50169 23069 50203 23103
rect 50905 23069 50939 23103
rect 51181 23069 51215 23103
rect 51365 23069 51399 23103
rect 51549 23069 51583 23103
rect 51641 23069 51675 23103
rect 51825 23069 51859 23103
rect 51917 23069 51951 23103
rect 52101 23069 52135 23103
rect 52193 23069 52227 23103
rect 52377 23069 52411 23103
rect 52469 23069 52503 23103
rect 52653 23069 52687 23103
rect 52745 23069 52779 23103
rect 52929 23069 52963 23103
rect 53481 23069 53515 23103
rect 53665 23069 53699 23103
rect 55321 23069 55355 23103
rect 55505 23069 55539 23103
rect 55597 23069 55631 23103
rect 55781 23069 55815 23103
rect 56701 23069 56735 23103
rect 57345 23069 57379 23103
rect 57529 23069 57563 23103
rect 57621 23069 57655 23103
rect 57989 23069 58023 23103
rect 58173 23069 58207 23103
rect 58265 23069 58299 23103
rect 1593 23001 1627 23035
rect 7665 23001 7699 23035
rect 37749 23001 37783 23035
rect 40141 23001 40175 23035
rect 41889 23001 41923 23035
rect 45293 23001 45327 23035
rect 47593 23001 47627 23035
rect 49157 23001 49191 23035
rect 51733 23001 51767 23035
rect 52009 23001 52043 23035
rect 55413 23001 55447 23035
rect 57805 23001 57839 23035
rect 3525 22933 3559 22967
rect 6653 22933 6687 22967
rect 10149 22933 10183 22967
rect 12909 22933 12943 22967
rect 42257 22933 42291 22967
rect 47041 22933 47075 22967
rect 47961 22933 47995 22967
rect 50813 22933 50847 22967
rect 51457 22933 51491 22967
rect 52285 22933 52319 22967
rect 53573 22933 53607 22967
rect 56057 22933 56091 22967
rect 1409 22729 1443 22763
rect 8677 22729 8711 22763
rect 9965 22729 9999 22763
rect 39405 22729 39439 22763
rect 40325 22729 40359 22763
rect 43913 22729 43947 22763
rect 45569 22729 45603 22763
rect 46673 22729 46707 22763
rect 47409 22729 47443 22763
rect 47961 22729 47995 22763
rect 49065 22729 49099 22763
rect 53297 22729 53331 22763
rect 53573 22729 53607 22763
rect 55321 22729 55355 22763
rect 57069 22729 57103 22763
rect 57437 22729 57471 22763
rect 58081 22729 58115 22763
rect 58357 22729 58391 22763
rect 9321 22661 9355 22695
rect 12633 22661 12667 22695
rect 12909 22661 12943 22695
rect 46305 22661 46339 22695
rect 48973 22661 49007 22695
rect 50537 22661 50571 22695
rect 54953 22661 54987 22695
rect 56793 22661 56827 22695
rect 3157 22593 3191 22627
rect 3985 22593 4019 22627
rect 4169 22593 4203 22627
rect 4537 22593 4571 22627
rect 4721 22593 4755 22627
rect 7941 22593 7975 22627
rect 8125 22593 8159 22627
rect 8217 22593 8251 22627
rect 9137 22593 9171 22627
rect 9781 22593 9815 22627
rect 9873 22593 9907 22627
rect 11078 22593 11112 22627
rect 12449 22593 12483 22627
rect 12725 22593 12759 22627
rect 12817 22593 12851 22627
rect 13001 22593 13035 22627
rect 40509 22593 40543 22627
rect 43361 22593 43395 22627
rect 44005 22593 44039 22627
rect 44189 22593 44223 22627
rect 46213 22593 46247 22627
rect 46581 22593 46615 22627
rect 46673 22593 46707 22627
rect 46857 22593 46891 22627
rect 47133 22593 47167 22627
rect 47225 22593 47259 22627
rect 47409 22593 47443 22627
rect 47593 22593 47627 22627
rect 47777 22593 47811 22627
rect 47869 22593 47903 22627
rect 48053 22593 48087 22627
rect 53481 22593 53515 22627
rect 53665 22593 53699 22627
rect 55137 22593 55171 22627
rect 55321 22593 55355 22627
rect 56977 22593 57011 22627
rect 57161 22593 57195 22627
rect 57253 22593 57287 22627
rect 57437 22593 57471 22627
rect 58265 22593 58299 22627
rect 58541 22593 58575 22627
rect 2881 22525 2915 22559
rect 3893 22525 3927 22559
rect 4077 22525 4111 22559
rect 9505 22525 9539 22559
rect 9597 22525 9631 22559
rect 11345 22525 11379 22559
rect 39773 22525 39807 22559
rect 42993 22525 43027 22559
rect 43637 22525 43671 22559
rect 46305 22525 46339 22559
rect 46489 22525 46523 22559
rect 50813 22525 50847 22559
rect 47041 22457 47075 22491
rect 47777 22457 47811 22491
rect 3249 22389 3283 22423
rect 4629 22389 4663 22423
rect 8033 22389 8067 22423
rect 8309 22389 8343 22423
rect 9689 22389 9723 22423
rect 11897 22389 11931 22423
rect 12449 22389 12483 22423
rect 42441 22389 42475 22423
rect 43453 22389 43487 22423
rect 44005 22389 44039 22423
rect 3341 22185 3375 22219
rect 5549 22185 5583 22219
rect 7389 22185 7423 22219
rect 9597 22185 9631 22219
rect 9965 22185 9999 22219
rect 11713 22185 11747 22219
rect 41232 22185 41266 22219
rect 43269 22185 43303 22219
rect 54769 22185 54803 22219
rect 55413 22185 55447 22219
rect 57529 22185 57563 22219
rect 2329 22117 2363 22151
rect 5733 22117 5767 22151
rect 5917 22117 5951 22151
rect 10424 22117 10458 22151
rect 55505 22117 55539 22151
rect 57621 22117 57655 22151
rect 2513 22049 2547 22083
rect 8769 22049 8803 22083
rect 11529 22049 11563 22083
rect 12081 22049 12115 22083
rect 40969 22049 41003 22083
rect 47409 22049 47443 22083
rect 49617 22049 49651 22083
rect 52561 22049 52595 22083
rect 53297 22049 53331 22083
rect 55045 22049 55079 22083
rect 55321 22049 55355 22083
rect 57069 22049 57103 22083
rect 57437 22049 57471 22083
rect 2237 21981 2271 22015
rect 2697 21981 2731 22015
rect 3433 21981 3467 22015
rect 3617 21981 3651 22015
rect 3893 21981 3927 22015
rect 3985 21981 4019 22015
rect 4169 21981 4203 22015
rect 5641 21981 5675 22015
rect 5825 21981 5859 22015
rect 7297 21981 7331 22015
rect 10149 21981 10183 22015
rect 10241 21981 10275 22015
rect 11805 21981 11839 22015
rect 12265 21981 12299 22015
rect 12357 21981 12391 22015
rect 12541 21981 12575 22015
rect 42809 21981 42843 22015
rect 44097 21981 44131 22015
rect 44281 21981 44315 22015
rect 44465 21981 44499 22015
rect 45661 21981 45695 22015
rect 45753 21981 45787 22015
rect 47133 21981 47167 22015
rect 48329 21981 48363 22015
rect 49341 21981 49375 22015
rect 51181 21981 51215 22015
rect 51733 21981 51767 22015
rect 52009 21981 52043 22015
rect 52469 21981 52503 22015
rect 52653 21981 52687 22015
rect 53573 21981 53607 22015
rect 54125 21981 54159 22015
rect 54585 21981 54619 22015
rect 54677 21981 54711 22015
rect 54861 21981 54895 22015
rect 54953 21981 54987 22015
rect 55137 21981 55171 22015
rect 55597 21981 55631 22015
rect 55965 21981 55999 22015
rect 56701 21981 56735 22015
rect 56885 21981 56919 22015
rect 56977 21981 57011 22015
rect 57161 21981 57195 22015
rect 57713 21981 57747 22015
rect 57805 21981 57839 22015
rect 57989 21981 58023 22015
rect 58081 21981 58115 22015
rect 58541 21981 58575 22015
rect 2513 21913 2547 21947
rect 4436 21913 4470 21947
rect 7030 21913 7064 21947
rect 8502 21913 8536 21947
rect 10425 21913 10459 21947
rect 12786 21913 12820 21947
rect 48605 21913 48639 21947
rect 51457 21913 51491 21947
rect 54309 21913 54343 21947
rect 54493 21913 54527 21947
rect 56609 21913 56643 21947
rect 56793 21913 56827 21947
rect 57897 21913 57931 21947
rect 3433 21845 3467 21879
rect 11529 21845 11563 21879
rect 13921 21845 13955 21879
rect 42717 21845 42751 21879
rect 42993 21845 43027 21879
rect 43545 21845 43579 21879
rect 44281 21845 44315 21879
rect 45017 21845 45051 21879
rect 46397 21845 46431 21879
rect 49249 21845 49283 21879
rect 52745 21845 52779 21879
rect 54585 21845 54619 21879
rect 58265 21845 58299 21879
rect 58357 21845 58391 21879
rect 4169 21641 4203 21675
rect 6554 21641 6588 21675
rect 7021 21641 7055 21675
rect 8039 21641 8073 21675
rect 42717 21641 42751 21675
rect 43085 21641 43119 21675
rect 43361 21641 43395 21675
rect 46673 21641 46707 21675
rect 54125 21641 54159 21675
rect 54309 21641 54343 21675
rect 55873 21641 55907 21675
rect 58541 21641 58575 21675
rect 4537 21573 4571 21607
rect 7941 21573 7975 21607
rect 44557 21573 44591 21607
rect 46121 21573 46155 21607
rect 50261 21573 50295 21607
rect 51273 21573 51307 21607
rect 2697 21505 2731 21539
rect 4721 21505 4755 21539
rect 4813 21505 4847 21539
rect 5917 21505 5951 21539
rect 6009 21505 6043 21539
rect 6377 21505 6411 21539
rect 6469 21505 6503 21539
rect 6653 21505 6687 21539
rect 8125 21505 8159 21539
rect 8217 21505 8251 21539
rect 42533 21505 42567 21539
rect 42717 21505 42751 21539
rect 42809 21505 42843 21539
rect 43913 21505 43947 21539
rect 44281 21505 44315 21539
rect 44373 21505 44407 21539
rect 46397 21505 46431 21539
rect 49157 21505 49191 21539
rect 49249 21505 49283 21539
rect 49433 21505 49467 21539
rect 49525 21505 49559 21539
rect 49617 21505 49651 21539
rect 49801 21505 49835 21539
rect 49893 21505 49927 21539
rect 50077 21505 50111 21539
rect 50169 21505 50203 21539
rect 50353 21505 50387 21539
rect 50537 21505 50571 21539
rect 50721 21505 50755 21539
rect 50813 21505 50847 21539
rect 50997 21505 51031 21539
rect 52193 21505 52227 21539
rect 52285 21505 52319 21539
rect 52745 21505 52779 21539
rect 53001 21505 53035 21539
rect 54217 21505 54251 21539
rect 54493 21505 54527 21539
rect 54760 21505 54794 21539
rect 56609 21505 56643 21539
rect 57529 21505 57563 21539
rect 1593 21437 1627 21471
rect 3709 21437 3743 21471
rect 10701 21437 10735 21471
rect 11529 21437 11563 21471
rect 43085 21437 43119 21471
rect 43637 21437 43671 21471
rect 44557 21437 44591 21471
rect 48421 21437 48455 21471
rect 48605 21437 48639 21471
rect 50905 21437 50939 21471
rect 52469 21437 52503 21471
rect 57897 21437 57931 21471
rect 4537 21369 4571 21403
rect 12541 21369 12575 21403
rect 49249 21369 49283 21403
rect 49985 21369 50019 21403
rect 52377 21369 52411 21403
rect 3157 21301 3191 21335
rect 10057 21301 10091 21335
rect 12173 21301 12207 21335
rect 42901 21301 42935 21335
rect 43821 21301 43855 21335
rect 44649 21301 44683 21335
rect 47777 21301 47811 21335
rect 49709 21301 49743 21335
rect 50629 21301 50663 21335
rect 55965 21301 55999 21335
rect 56885 21301 56919 21335
rect 3341 21097 3375 21131
rect 4629 21097 4663 21131
rect 6377 21097 6411 21131
rect 8309 21097 8343 21131
rect 9781 21097 9815 21131
rect 44741 21097 44775 21131
rect 45845 21097 45879 21131
rect 50445 21097 50479 21131
rect 51549 21097 51583 21131
rect 54861 21097 54895 21131
rect 57805 21097 57839 21131
rect 54953 21029 54987 21063
rect 56149 21029 56183 21063
rect 58081 21029 58115 21063
rect 2881 20961 2915 20995
rect 3249 20961 3283 20995
rect 3801 20961 3835 20995
rect 9873 20961 9907 20995
rect 11621 20961 11655 20995
rect 11897 20961 11931 20995
rect 43545 20961 43579 20995
rect 43821 20961 43855 20995
rect 46213 20961 46247 20995
rect 54769 20961 54803 20995
rect 56333 20961 56367 20995
rect 3157 20893 3191 20927
rect 3433 20893 3467 20927
rect 3525 20893 3559 20927
rect 4353 20893 4387 20927
rect 4997 20893 5031 20927
rect 6561 20893 6595 20927
rect 9597 20893 9631 20927
rect 9689 20893 9723 20927
rect 13737 20893 13771 20927
rect 14289 20893 14323 20927
rect 43453 20893 43487 20927
rect 44373 20893 44407 20927
rect 45017 20893 45051 20927
rect 45753 20893 45787 20927
rect 45937 20893 45971 20927
rect 47869 20893 47903 20927
rect 49157 20893 49191 20927
rect 49341 20893 49375 20927
rect 49525 20893 49559 20927
rect 49617 20893 49651 20927
rect 49801 20893 49835 20927
rect 50169 20893 50203 20927
rect 50353 20893 50387 20927
rect 50445 20893 50479 20927
rect 50629 20893 50663 20927
rect 51457 20893 51491 20927
rect 51641 20893 51675 20927
rect 55045 20893 55079 20927
rect 55965 20893 55999 20927
rect 56057 20893 56091 20927
rect 56425 20893 56459 20927
rect 57989 20893 58023 20927
rect 58173 20893 58207 20927
rect 58265 20893 58299 20927
rect 4813 20825 4847 20859
rect 6745 20825 6779 20859
rect 8493 20825 8527 20859
rect 8677 20825 8711 20859
rect 11989 20825 12023 20859
rect 44557 20825 44591 20859
rect 46480 20825 46514 20859
rect 48605 20825 48639 20859
rect 49709 20825 49743 20859
rect 50261 20825 50295 20859
rect 56333 20825 56367 20859
rect 56670 20825 56704 20859
rect 1409 20757 1443 20791
rect 10149 20757 10183 20791
rect 45201 20757 45235 20791
rect 47593 20757 47627 20791
rect 48513 20757 48547 20791
rect 49433 20757 49467 20791
rect 55321 20757 55355 20791
rect 58357 20757 58391 20791
rect 3985 20553 4019 20587
rect 6561 20553 6595 20587
rect 8125 20553 8159 20587
rect 10977 20553 11011 20587
rect 13185 20553 13219 20587
rect 19717 20553 19751 20587
rect 47317 20553 47351 20587
rect 48789 20553 48823 20587
rect 49433 20553 49467 20587
rect 51917 20553 51951 20587
rect 56333 20553 56367 20587
rect 3341 20485 3375 20519
rect 12909 20485 12943 20519
rect 47593 20485 47627 20519
rect 48329 20485 48363 20519
rect 53021 20485 53055 20519
rect 57345 20485 57379 20519
rect 2697 20417 2731 20451
rect 3525 20417 3559 20451
rect 3709 20417 3743 20451
rect 3801 20417 3835 20451
rect 3985 20417 4019 20451
rect 5374 20417 5408 20451
rect 6377 20417 6411 20451
rect 6653 20417 6687 20451
rect 6745 20417 6779 20451
rect 6929 20417 6963 20451
rect 7941 20417 7975 20451
rect 8217 20417 8251 20451
rect 8309 20417 8343 20451
rect 8493 20417 8527 20451
rect 10793 20417 10827 20451
rect 10885 20417 10919 20451
rect 11069 20417 11103 20451
rect 18245 20417 18279 20451
rect 47225 20417 47259 20451
rect 47409 20417 47443 20451
rect 48513 20417 48547 20451
rect 48605 20417 48639 20451
rect 48697 20417 48731 20451
rect 48881 20417 48915 20451
rect 51831 20417 51865 20451
rect 52009 20417 52043 20451
rect 52561 20417 52595 20451
rect 52745 20417 52779 20451
rect 56241 20417 56275 20451
rect 56425 20417 56459 20451
rect 57437 20417 57471 20451
rect 57713 20417 57747 20451
rect 5641 20349 5675 20383
rect 6837 20349 6871 20383
rect 8401 20349 8435 20383
rect 10149 20349 10183 20383
rect 12081 20349 12115 20383
rect 48145 20349 48179 20383
rect 56149 20349 56183 20383
rect 58541 20349 58575 20383
rect 4261 20281 4295 20315
rect 57529 20281 57563 20315
rect 3617 20213 3651 20247
rect 6377 20213 6411 20247
rect 7941 20213 7975 20247
rect 20361 20213 20395 20247
rect 47041 20213 47075 20247
rect 48329 20213 48363 20247
rect 55505 20213 55539 20247
rect 57897 20213 57931 20247
rect 4721 20009 4755 20043
rect 11713 20009 11747 20043
rect 49709 20009 49743 20043
rect 51181 20009 51215 20043
rect 51825 20009 51859 20043
rect 53113 20009 53147 20043
rect 56701 20009 56735 20043
rect 58173 20009 58207 20043
rect 5917 19941 5951 19975
rect 50813 19941 50847 19975
rect 53573 19941 53607 19975
rect 58357 19941 58391 19975
rect 7297 19873 7331 19907
rect 8769 19873 8803 19907
rect 47041 19873 47075 19907
rect 47961 19873 47995 19907
rect 50261 19873 50295 19907
rect 53389 19873 53423 19907
rect 55045 19873 55079 19907
rect 2605 19805 2639 19839
rect 2881 19805 2915 19839
rect 3801 19805 3835 19839
rect 3985 19805 4019 19839
rect 4077 19805 4111 19839
rect 4261 19805 4295 19839
rect 4445 19805 4479 19839
rect 4537 19805 4571 19839
rect 4721 19805 4755 19839
rect 4813 19805 4847 19839
rect 4997 19805 5031 19839
rect 7030 19805 7064 19839
rect 8502 19805 8536 19839
rect 10149 19805 10183 19839
rect 11437 19805 11471 19839
rect 11805 19805 11839 19839
rect 48605 19805 48639 19839
rect 49249 19805 49283 19839
rect 49341 19805 49375 19839
rect 49525 19805 49559 19839
rect 49617 19805 49651 19839
rect 49801 19805 49835 19839
rect 50169 19805 50203 19839
rect 50353 19805 50387 19839
rect 50445 19805 50479 19839
rect 50629 19805 50663 19839
rect 50721 19805 50755 19839
rect 50905 19805 50939 19839
rect 51733 19805 51767 19839
rect 51917 19805 51951 19839
rect 52009 19805 52043 19839
rect 52193 19805 52227 19839
rect 53297 19805 53331 19839
rect 53481 19805 53515 19839
rect 53573 19805 53607 19839
rect 54033 19805 54067 19839
rect 54125 19805 54159 19839
rect 54309 19805 54343 19839
rect 54953 19805 54987 19839
rect 55137 19805 55171 19839
rect 55321 19805 55355 19839
rect 56793 19805 56827 19839
rect 58265 19805 58299 19839
rect 1593 19737 1627 19771
rect 10793 19737 10827 19771
rect 46796 19737 46830 19771
rect 47317 19737 47351 19771
rect 48973 19737 49007 19771
rect 52101 19737 52135 19771
rect 53665 19737 53699 19771
rect 53849 19737 53883 19771
rect 55566 19737 55600 19771
rect 57060 19737 57094 19771
rect 3525 19669 3559 19703
rect 3801 19669 3835 19703
rect 4169 19669 4203 19703
rect 4813 19669 4847 19703
rect 7389 19669 7423 19703
rect 10885 19669 10919 19703
rect 12081 19669 12115 19703
rect 45661 19669 45695 19703
rect 48053 19669 48087 19703
rect 49433 19669 49467 19703
rect 50537 19669 50571 19703
rect 54033 19669 54067 19703
rect 1409 19465 1443 19499
rect 8861 19465 8895 19499
rect 9137 19465 9171 19499
rect 11805 19465 11839 19499
rect 49341 19465 49375 19499
rect 50445 19465 50479 19499
rect 51733 19465 51767 19499
rect 55045 19465 55079 19499
rect 56977 19465 57011 19499
rect 57437 19465 57471 19499
rect 10609 19397 10643 19431
rect 3157 19329 3191 19363
rect 3985 19329 4019 19363
rect 4169 19329 4203 19363
rect 8953 19329 8987 19363
rect 10885 19329 10919 19363
rect 10977 19329 11011 19363
rect 11161 19329 11195 19363
rect 47225 19329 47259 19363
rect 47409 19329 47443 19363
rect 49157 19329 49191 19363
rect 49341 19329 49375 19363
rect 49433 19329 49467 19363
rect 49617 19329 49651 19363
rect 49709 19329 49743 19363
rect 49893 19329 49927 19363
rect 50353 19329 50387 19363
rect 50537 19329 50571 19363
rect 51365 19329 51399 19363
rect 51641 19329 51675 19363
rect 51733 19329 51767 19363
rect 51917 19329 51951 19363
rect 54769 19329 54803 19363
rect 55413 19329 55447 19363
rect 55505 19329 55539 19363
rect 57253 19329 57287 19363
rect 57345 19329 57379 19363
rect 57529 19329 57563 19363
rect 2881 19261 2915 19295
rect 3893 19261 3927 19295
rect 4077 19261 4111 19295
rect 7665 19261 7699 19295
rect 8677 19261 8711 19295
rect 47317 19261 47351 19295
rect 48145 19261 48179 19295
rect 48881 19261 48915 19295
rect 49525 19261 49559 19295
rect 50261 19261 50295 19295
rect 55045 19261 55079 19295
rect 56977 19261 57011 19295
rect 57897 19261 57931 19295
rect 58449 19261 58483 19295
rect 57161 19193 57195 19227
rect 3249 19125 3283 19159
rect 8309 19125 8343 19159
rect 11069 19125 11103 19159
rect 47593 19125 47627 19159
rect 48329 19125 48363 19159
rect 49801 19125 49835 19159
rect 54861 19125 54895 19159
rect 3341 18921 3375 18955
rect 4629 18921 4663 18955
rect 6745 18921 6779 18955
rect 9781 18921 9815 18955
rect 50169 18921 50203 18955
rect 51733 18921 51767 18955
rect 57621 18921 57655 18955
rect 58357 18921 58391 18955
rect 9689 18853 9723 18887
rect 48973 18853 49007 18887
rect 57069 18853 57103 18887
rect 2421 18785 2455 18819
rect 3525 18785 3559 18819
rect 4353 18785 4387 18819
rect 4813 18785 4847 18819
rect 6837 18785 6871 18819
rect 8493 18785 8527 18819
rect 8769 18785 8803 18819
rect 9873 18785 9907 18819
rect 10517 18785 10551 18819
rect 11069 18785 11103 18819
rect 47041 18785 47075 18819
rect 47593 18785 47627 18819
rect 52285 18785 52319 18819
rect 52469 18785 52503 18819
rect 52561 18785 52595 18819
rect 54677 18785 54711 18819
rect 54861 18785 54895 18819
rect 2145 18717 2179 18751
rect 2237 18717 2271 18751
rect 2697 18717 2731 18751
rect 3433 18717 3467 18751
rect 3617 18717 3651 18751
rect 4537 18717 4571 18751
rect 5273 18717 5307 18751
rect 6561 18717 6595 18751
rect 6653 18717 6687 18751
rect 9597 18717 9631 18751
rect 47133 18717 47167 18751
rect 47317 18717 47351 18751
rect 47860 18717 47894 18751
rect 49801 18717 49835 18751
rect 50169 18717 50203 18751
rect 50353 18717 50387 18751
rect 50445 18717 50479 18751
rect 50629 18717 50663 18751
rect 51549 18717 51583 18751
rect 51733 18717 51767 18751
rect 52193 18717 52227 18751
rect 54769 18717 54803 18751
rect 54953 18717 54987 18751
rect 57253 18717 57287 18751
rect 57437 18717 57471 18751
rect 57713 18717 57747 18751
rect 57897 18717 57931 18751
rect 58081 18717 58115 18751
rect 58541 18717 58575 18751
rect 2421 18649 2455 18683
rect 4813 18649 4847 18683
rect 46796 18649 46830 18683
rect 52469 18649 52503 18683
rect 52806 18649 52840 18683
rect 54033 18649 54067 18683
rect 57345 18649 57379 18683
rect 3801 18581 3835 18615
rect 5917 18581 5951 18615
rect 7021 18581 7055 18615
rect 45661 18581 45695 18615
rect 47317 18581 47351 18615
rect 49157 18581 49191 18615
rect 50537 18581 50571 18615
rect 53941 18581 53975 18615
rect 57989 18581 58023 18615
rect 3709 18377 3743 18411
rect 7941 18377 7975 18411
rect 47225 18377 47259 18411
rect 48421 18377 48455 18411
rect 49341 18377 49375 18411
rect 51917 18377 51951 18411
rect 53021 18377 53055 18411
rect 54677 18377 54711 18411
rect 57345 18377 57379 18411
rect 58357 18377 58391 18411
rect 9873 18309 9907 18343
rect 49433 18309 49467 18343
rect 51641 18309 51675 18343
rect 52193 18309 52227 18343
rect 53757 18309 53791 18343
rect 2697 18241 2731 18275
rect 4261 18241 4295 18275
rect 6929 18241 6963 18275
rect 7113 18241 7147 18275
rect 7205 18241 7239 18275
rect 7757 18241 7791 18275
rect 9597 18241 9631 18275
rect 11529 18241 11563 18275
rect 46949 18241 46983 18275
rect 47041 18241 47075 18275
rect 47225 18241 47259 18275
rect 48145 18241 48179 18275
rect 48329 18241 48363 18275
rect 48513 18241 48547 18275
rect 49157 18241 49191 18275
rect 49341 18241 49375 18275
rect 51273 18241 51307 18275
rect 51457 18241 51491 18275
rect 51549 18241 51583 18275
rect 51733 18241 51767 18275
rect 51825 18241 51859 18275
rect 52009 18241 52043 18275
rect 52101 18241 52135 18275
rect 52285 18241 52319 18275
rect 53113 18241 53147 18275
rect 53665 18241 53699 18275
rect 53941 18241 53975 18275
rect 54033 18241 54067 18275
rect 55965 18241 55999 18275
rect 57713 18241 57747 18275
rect 57897 18241 57931 18275
rect 57989 18241 58023 18275
rect 58173 18241 58207 18275
rect 58541 18241 58575 18275
rect 1593 18173 1627 18207
rect 3525 18173 3559 18207
rect 5917 18173 5951 18207
rect 6193 18173 6227 18207
rect 8493 18173 8527 18207
rect 9873 18173 9907 18207
rect 10149 18173 10183 18207
rect 10793 18173 10827 18207
rect 46305 18173 46339 18207
rect 47593 18173 47627 18207
rect 7021 18105 7055 18139
rect 9689 18105 9723 18139
rect 57529 18105 57563 18139
rect 2973 18037 3007 18071
rect 4445 18037 4479 18071
rect 9229 18037 9263 18071
rect 12173 18037 12207 18071
rect 46121 18037 46155 18071
rect 49065 18037 49099 18071
rect 50905 18037 50939 18071
rect 51365 18037 51399 18071
rect 53665 18037 53699 18071
rect 55873 18037 55907 18071
rect 58081 18037 58115 18071
rect 1409 17833 1443 17867
rect 3341 17833 3375 17867
rect 4813 17833 4847 17867
rect 12265 17833 12299 17867
rect 49709 17833 49743 17867
rect 50169 17833 50203 17867
rect 54033 17833 54067 17867
rect 54953 17833 54987 17867
rect 58265 17833 58299 17867
rect 8585 17765 8619 17799
rect 49433 17765 49467 17799
rect 56701 17765 56735 17799
rect 57805 17765 57839 17799
rect 2881 17697 2915 17731
rect 3249 17697 3283 17731
rect 4629 17697 4663 17731
rect 5365 17697 5399 17731
rect 6101 17697 6135 17731
rect 8677 17697 8711 17731
rect 9413 17697 9447 17731
rect 11989 17697 12023 17731
rect 53389 17697 53423 17731
rect 55137 17697 55171 17731
rect 56793 17697 56827 17731
rect 3157 17629 3191 17663
rect 3433 17629 3467 17663
rect 3525 17629 3559 17663
rect 4537 17629 4571 17663
rect 4721 17629 4755 17663
rect 5549 17629 5583 17663
rect 8401 17629 8435 17663
rect 8493 17629 8527 17663
rect 9137 17629 9171 17663
rect 47869 17629 47903 17663
rect 49157 17629 49191 17663
rect 50169 17629 50203 17663
rect 50353 17629 50387 17663
rect 53297 17629 53331 17663
rect 53481 17629 53515 17663
rect 53573 17629 53607 17663
rect 53849 17629 53883 17663
rect 53941 17629 53975 17663
rect 54125 17629 54159 17663
rect 54861 17629 54895 17663
rect 55321 17629 55355 17663
rect 57529 17629 57563 17663
rect 57805 17629 57839 17663
rect 57897 17629 57931 17663
rect 58056 17631 58090 17665
rect 58173 17629 58207 17663
rect 58357 17629 58391 17663
rect 9045 17561 9079 17595
rect 11713 17561 11747 17595
rect 49433 17561 49467 17595
rect 53665 17561 53699 17595
rect 55137 17561 55171 17595
rect 55566 17561 55600 17595
rect 57713 17561 57747 17595
rect 10057 17493 10091 17527
rect 10241 17493 10275 17527
rect 47317 17493 47351 17527
rect 49249 17493 49283 17527
rect 53113 17493 53147 17527
rect 53757 17493 53791 17527
rect 57437 17493 57471 17527
rect 58081 17493 58115 17527
rect 9045 17289 9079 17323
rect 11069 17289 11103 17323
rect 47685 17289 47719 17323
rect 49157 17289 49191 17323
rect 55597 17289 55631 17323
rect 57253 17289 57287 17323
rect 58357 17289 58391 17323
rect 2697 17221 2731 17255
rect 4721 17221 4755 17255
rect 6745 17221 6779 17255
rect 48973 17221 49007 17255
rect 2421 17153 2455 17187
rect 2789 17153 2823 17187
rect 4445 17153 4479 17187
rect 4813 17153 4847 17187
rect 6469 17153 6503 17187
rect 6561 17153 6595 17187
rect 6837 17153 6871 17187
rect 8953 17153 8987 17187
rect 9781 17153 9815 17187
rect 9965 17153 9999 17187
rect 10885 17153 10919 17187
rect 10977 17153 11011 17187
rect 11161 17153 11195 17187
rect 47225 17153 47259 17187
rect 47593 17153 47627 17187
rect 47777 17153 47811 17187
rect 48605 17153 48639 17187
rect 48697 17153 48731 17187
rect 48789 17153 48823 17187
rect 49065 17153 49099 17187
rect 49249 17153 49283 17187
rect 49341 17153 49375 17187
rect 49525 17153 49559 17187
rect 56333 17153 56367 17187
rect 56517 17153 56551 17187
rect 57069 17153 57103 17187
rect 57253 17153 57287 17187
rect 57621 17153 57655 17187
rect 57989 17153 58023 17187
rect 58173 17153 58207 17187
rect 58541 17153 58575 17187
rect 2513 17085 2547 17119
rect 2697 17085 2731 17119
rect 3525 17085 3559 17119
rect 4169 17085 4203 17119
rect 4721 17085 4755 17119
rect 5549 17085 5583 17119
rect 6193 17085 6227 17119
rect 6745 17085 6779 17119
rect 7573 17085 7607 17119
rect 8125 17085 8159 17119
rect 8401 17085 8435 17119
rect 9689 17085 9723 17119
rect 9873 17085 9907 17119
rect 10241 17085 10275 17119
rect 46949 17085 46983 17119
rect 48053 17085 48087 17119
rect 48973 17085 49007 17119
rect 49433 17085 49467 17119
rect 56241 17085 56275 17119
rect 56425 17085 56459 17119
rect 58081 17017 58115 17051
rect 3433 16949 3467 16983
rect 4537 16949 4571 16983
rect 5457 16949 5491 16983
rect 7481 16949 7515 16983
rect 47041 16949 47075 16983
rect 47133 16949 47167 16983
rect 53113 16949 53147 16983
rect 3175 16745 3209 16779
rect 5837 16745 5871 16779
rect 6285 16745 6319 16779
rect 8229 16745 8263 16779
rect 10529 16745 10563 16779
rect 48053 16745 48087 16779
rect 48881 16745 48915 16779
rect 49801 16745 49835 16779
rect 52929 16745 52963 16779
rect 53665 16745 53699 16779
rect 57805 16745 57839 16779
rect 57989 16745 58023 16779
rect 51549 16677 51583 16711
rect 54217 16677 54251 16711
rect 56425 16677 56459 16711
rect 58357 16677 58391 16711
rect 3433 16609 3467 16643
rect 6101 16609 6135 16643
rect 8493 16609 8527 16643
rect 10793 16609 10827 16643
rect 46673 16609 46707 16643
rect 49985 16609 50019 16643
rect 50169 16609 50203 16643
rect 51641 16609 51675 16643
rect 3801 16541 3835 16575
rect 3985 16541 4019 16575
rect 6193 16541 6227 16575
rect 6377 16541 6411 16575
rect 46940 16541 46974 16575
rect 49709 16541 49743 16575
rect 52469 16541 52503 16575
rect 52561 16541 52595 16575
rect 52653 16541 52687 16575
rect 53205 16541 53239 16575
rect 53297 16541 53331 16575
rect 53481 16541 53515 16575
rect 53665 16541 53699 16575
rect 53757 16541 53791 16575
rect 55597 16541 55631 16575
rect 56609 16541 56643 16575
rect 58173 16541 58207 16575
rect 58541 16541 58575 16575
rect 3893 16473 3927 16507
rect 49985 16473 50019 16507
rect 50414 16473 50448 16507
rect 52929 16473 52963 16507
rect 53941 16473 53975 16507
rect 57897 16473 57931 16507
rect 58081 16473 58115 16507
rect 1685 16405 1719 16439
rect 4353 16405 4387 16439
rect 6745 16405 6779 16439
rect 9045 16405 9079 16439
rect 52285 16405 52319 16439
rect 52837 16405 52871 16439
rect 53113 16405 53147 16439
rect 53297 16405 53331 16439
rect 55505 16405 55539 16439
rect 57253 16405 57287 16439
rect 3525 16201 3559 16235
rect 6377 16201 6411 16235
rect 7297 16201 7331 16235
rect 48513 16201 48547 16235
rect 48881 16201 48915 16235
rect 49157 16201 49191 16235
rect 49709 16201 49743 16235
rect 50353 16201 50387 16235
rect 53021 16201 53055 16235
rect 53573 16201 53607 16235
rect 54125 16201 54159 16235
rect 56517 16201 56551 16235
rect 58173 16201 58207 16235
rect 44097 16133 44131 16167
rect 44189 16133 44223 16167
rect 52193 16133 52227 16167
rect 54401 16133 54435 16167
rect 57529 16133 57563 16167
rect 57989 16133 58023 16167
rect 1593 16065 1627 16099
rect 2697 16065 2731 16099
rect 7205 16065 7239 16099
rect 7389 16065 7423 16099
rect 7941 16065 7975 16099
rect 45937 16065 45971 16099
rect 47869 16065 47903 16099
rect 48053 16065 48087 16099
rect 48421 16065 48455 16099
rect 48605 16065 48639 16099
rect 48789 16065 48823 16099
rect 49065 16065 49099 16099
rect 49157 16065 49191 16099
rect 49341 16065 49375 16099
rect 51089 16065 51123 16099
rect 51273 16065 51307 16099
rect 52101 16065 52135 16099
rect 52285 16065 52319 16099
rect 52837 16065 52871 16099
rect 53021 16065 53055 16099
rect 53573 16065 53607 16099
rect 53757 16065 53791 16099
rect 54125 16065 54159 16099
rect 54217 16065 54251 16099
rect 55404 16065 55438 16099
rect 57345 16065 57379 16099
rect 57621 16065 57655 16099
rect 57897 16065 57931 16099
rect 58081 16065 58115 16099
rect 58173 16065 58207 16099
rect 58357 16065 58391 16099
rect 2881 15997 2915 16031
rect 6929 15997 6963 16031
rect 8493 15997 8527 16031
rect 50997 15997 51031 16031
rect 51181 15997 51215 16031
rect 55137 15997 55171 16031
rect 57161 15997 57195 16031
rect 57621 15929 57655 15963
rect 47961 15861 47995 15895
rect 49065 15861 49099 15895
rect 56609 15861 56643 15895
rect 49709 15657 49743 15691
rect 50261 15657 50295 15691
rect 51917 15657 51951 15691
rect 53481 15657 53515 15691
rect 53757 15657 53791 15691
rect 55505 15657 55539 15691
rect 56701 15657 56735 15691
rect 57989 15657 58023 15691
rect 58265 15657 58299 15691
rect 47409 15589 47443 15623
rect 52561 15589 52595 15623
rect 57253 15589 57287 15623
rect 46029 15521 46063 15555
rect 48053 15521 48087 15555
rect 55597 15521 55631 15555
rect 48789 15453 48823 15487
rect 49065 15453 49099 15487
rect 49249 15453 49283 15487
rect 49341 15453 49375 15487
rect 49479 15453 49513 15487
rect 50537 15453 50571 15487
rect 50629 15453 50663 15487
rect 50721 15453 50755 15487
rect 50905 15453 50939 15487
rect 51641 15453 51675 15487
rect 51917 15453 51951 15487
rect 52101 15453 52135 15487
rect 52285 15453 52319 15487
rect 53573 15453 53607 15487
rect 55321 15453 55355 15487
rect 55413 15453 55447 15487
rect 56609 15453 56643 15487
rect 56793 15453 56827 15487
rect 57529 15453 57563 15487
rect 57713 15453 57747 15487
rect 57897 15453 57931 15487
rect 58081 15453 58115 15487
rect 58173 15453 58207 15487
rect 58357 15453 58391 15487
rect 46296 15385 46330 15419
rect 53665 15385 53699 15419
rect 53849 15385 53883 15419
rect 57621 15385 57655 15419
rect 47501 15317 47535 15351
rect 48237 15317 48271 15351
rect 51733 15317 51767 15351
rect 52193 15317 52227 15351
rect 56517 15317 56551 15351
rect 46581 15113 46615 15147
rect 47869 15113 47903 15147
rect 49157 15113 49191 15147
rect 49249 15113 49283 15147
rect 50353 15113 50387 15147
rect 51089 15113 51123 15147
rect 51549 15113 51583 15147
rect 52837 15113 52871 15147
rect 53205 15113 53239 15147
rect 53573 15113 53607 15147
rect 54033 15113 54067 15147
rect 56885 15113 56919 15147
rect 57713 15113 57747 15147
rect 54125 15045 54159 15079
rect 2697 14977 2731 15011
rect 46857 14977 46891 15011
rect 47593 14977 47627 15011
rect 47685 14977 47719 15011
rect 48145 14977 48179 15011
rect 48329 14977 48363 15011
rect 48513 14977 48547 15011
rect 48697 14977 48731 15011
rect 48789 14977 48823 15011
rect 48881 14977 48915 15011
rect 49249 14977 49283 15011
rect 49433 14977 49467 15011
rect 50629 14977 50663 15011
rect 50721 14977 50755 15011
rect 50813 14977 50847 15011
rect 50997 14977 51031 15011
rect 51089 14977 51123 15011
rect 51273 14977 51307 15011
rect 51457 14977 51491 15011
rect 51641 14977 51675 15011
rect 52745 14977 52779 15011
rect 52929 14977 52963 15011
rect 53021 14977 53055 15011
rect 53205 14977 53239 15011
rect 53573 14977 53607 15011
rect 53757 14977 53791 15011
rect 54033 14977 54067 15011
rect 54309 14977 54343 15011
rect 58449 14977 58483 15011
rect 1593 14909 1627 14943
rect 46581 14909 46615 14943
rect 47869 14909 47903 14943
rect 48237 14909 48271 14943
rect 49709 14909 49743 14943
rect 50169 14909 50203 14943
rect 56149 14909 56183 14943
rect 57161 14909 57195 14943
rect 46765 14841 46799 14875
rect 55505 14773 55539 14807
rect 57897 14773 57931 14807
rect 48421 14569 48455 14603
rect 48605 14569 48639 14603
rect 49249 14569 49283 14603
rect 50537 14569 50571 14603
rect 52377 14569 52411 14603
rect 58265 14569 58299 14603
rect 50905 14501 50939 14535
rect 56701 14501 56735 14535
rect 58357 14501 58391 14535
rect 48513 14365 48547 14399
rect 48697 14365 48731 14399
rect 49157 14365 49191 14399
rect 49341 14365 49375 14399
rect 50445 14365 50479 14399
rect 50629 14365 50663 14399
rect 52285 14365 52319 14399
rect 52469 14365 52503 14399
rect 55137 14365 55171 14399
rect 55321 14365 55355 14399
rect 56885 14365 56919 14399
rect 58541 14365 58575 14399
rect 55566 14297 55600 14331
rect 57130 14297 57164 14331
rect 55045 14229 55079 14263
rect 47869 14025 47903 14059
rect 49341 14025 49375 14059
rect 51273 14025 51307 14059
rect 51457 14025 51491 14059
rect 52745 14025 52779 14059
rect 54217 14025 54251 14059
rect 55137 14025 55171 14059
rect 56333 14025 56367 14059
rect 56793 14025 56827 14059
rect 58357 14025 58391 14059
rect 47593 13889 47627 13923
rect 47685 13889 47719 13923
rect 47961 13889 47995 13923
rect 48145 13889 48179 13923
rect 48329 13889 48363 13923
rect 48421 13889 48455 13923
rect 49065 13889 49099 13923
rect 50997 13889 51031 13923
rect 51181 13889 51215 13923
rect 51273 13889 51307 13923
rect 51365 13889 51399 13923
rect 51549 13889 51583 13923
rect 51825 13889 51859 13923
rect 52929 13911 52963 13945
rect 53021 13889 53055 13923
rect 53113 13889 53147 13923
rect 53849 13889 53883 13923
rect 54033 13889 54067 13923
rect 54125 13889 54159 13923
rect 54217 13889 54251 13923
rect 54401 13889 54435 13923
rect 54861 13889 54895 13923
rect 56149 13889 56183 13923
rect 56241 13889 56275 13923
rect 56425 13889 56459 13923
rect 56517 13889 56551 13923
rect 58173 13889 58207 13923
rect 58265 13889 58299 13923
rect 58541 13889 58575 13923
rect 47869 13821 47903 13855
rect 48053 13821 48087 13855
rect 49341 13821 49375 13855
rect 51733 13821 51767 13855
rect 55137 13821 55171 13855
rect 56793 13821 56827 13855
rect 49157 13753 49191 13787
rect 54125 13753 54159 13787
rect 55505 13753 55539 13787
rect 54953 13685 54987 13719
rect 56609 13685 56643 13719
rect 48513 13481 48547 13515
rect 49433 13481 49467 13515
rect 51733 13481 51767 13515
rect 53849 13481 53883 13515
rect 54585 13481 54619 13515
rect 56425 13481 56459 13515
rect 58357 13481 58391 13515
rect 47685 13413 47719 13447
rect 57897 13413 57931 13447
rect 46305 13345 46339 13379
rect 49065 13345 49099 13379
rect 56609 13345 56643 13379
rect 2789 13277 2823 13311
rect 48329 13277 48363 13311
rect 49341 13277 49375 13311
rect 49525 13277 49559 13311
rect 51457 13277 51491 13311
rect 51641 13277 51675 13311
rect 51825 13277 51859 13311
rect 52101 13277 52135 13311
rect 52193 13277 52227 13311
rect 53573 13277 53607 13311
rect 53757 13277 53791 13311
rect 53941 13277 53975 13311
rect 54677 13277 54711 13311
rect 56333 13277 56367 13311
rect 56977 13277 57011 13311
rect 57805 13277 57839 13311
rect 58081 13277 58115 13311
rect 58541 13277 58575 13311
rect 1593 13209 1627 13243
rect 46572 13209 46606 13243
rect 52009 13209 52043 13243
rect 56885 13209 56919 13243
rect 47777 13141 47811 13175
rect 50905 13141 50939 13175
rect 52837 13141 52871 13175
rect 52929 13141 52963 13175
rect 56609 13141 56643 13175
rect 57713 13141 57747 13175
rect 46857 12937 46891 12971
rect 47869 12937 47903 12971
rect 49985 12937 50019 12971
rect 51181 12937 51215 12971
rect 52101 12937 52135 12971
rect 54125 12937 54159 12971
rect 58541 12937 58575 12971
rect 50629 12869 50663 12903
rect 52561 12869 52595 12903
rect 56497 12869 56531 12903
rect 47041 12801 47075 12835
rect 47133 12801 47167 12835
rect 47777 12801 47811 12835
rect 47961 12791 47995 12825
rect 48697 12801 48731 12835
rect 50077 12801 50111 12835
rect 50353 12801 50387 12835
rect 51089 12801 51123 12835
rect 51273 12801 51307 12835
rect 52285 12801 52319 12835
rect 53001 12801 53035 12835
rect 54217 12801 54251 12835
rect 54677 12801 54711 12835
rect 54769 12801 54803 12835
rect 56241 12801 56275 12835
rect 46857 12733 46891 12767
rect 48421 12733 48455 12767
rect 49157 12733 49191 12767
rect 49709 12733 49743 12767
rect 50629 12733 50663 12767
rect 51549 12733 51583 12767
rect 52561 12733 52595 12767
rect 52745 12733 52779 12767
rect 54309 12733 54343 12767
rect 54493 12733 54527 12767
rect 55045 12733 55079 12767
rect 55689 12733 55723 12767
rect 57897 12733 57931 12767
rect 57621 12665 57655 12699
rect 48513 12597 48547 12631
rect 48605 12597 48639 12631
rect 50445 12597 50479 12631
rect 52377 12597 52411 12631
rect 54401 12597 54435 12631
rect 49801 12393 49835 12427
rect 51641 12393 51675 12427
rect 52101 12393 52135 12427
rect 55965 12393 55999 12427
rect 56149 12393 56183 12427
rect 56793 12393 56827 12427
rect 55137 12325 55171 12359
rect 58265 12325 58299 12359
rect 48237 12257 48271 12291
rect 55321 12257 55355 12291
rect 57437 12257 57471 12291
rect 57621 12257 57655 12291
rect 48504 12189 48538 12223
rect 49709 12189 49743 12223
rect 49893 12189 49927 12223
rect 50261 12189 50295 12223
rect 52009 12189 52043 12223
rect 52193 12189 52227 12223
rect 53757 12189 53791 12223
rect 54024 12189 54058 12223
rect 56057 12189 56091 12223
rect 56241 12189 56275 12223
rect 57529 12189 57563 12223
rect 57713 12189 57747 12223
rect 57897 12189 57931 12223
rect 58173 12189 58207 12223
rect 50528 12121 50562 12155
rect 49617 12053 49651 12087
rect 58081 12053 58115 12087
rect 50353 11849 50387 11883
rect 58081 11849 58115 11883
rect 2697 11713 2731 11747
rect 49709 11713 49743 11747
rect 57897 11713 57931 11747
rect 58173 11713 58207 11747
rect 1593 11645 1627 11679
rect 58265 11577 58299 11611
rect 49249 10761 49283 10795
rect 49341 10625 49375 10659
rect 58541 10625 58575 10659
rect 58357 10489 58391 10523
rect 58357 10217 58391 10251
rect 2697 10013 2731 10047
rect 58541 10013 58575 10047
rect 1593 9945 1627 9979
rect 58357 9129 58391 9163
rect 58541 8925 58575 8959
rect 58357 8585 58391 8619
rect 2697 8449 2731 8483
rect 58541 8449 58575 8483
rect 1593 8381 1627 8415
rect 58541 7361 58575 7395
rect 58357 7157 58391 7191
rect 2697 6749 2731 6783
rect 1593 6681 1627 6715
rect 2697 5185 2731 5219
rect 1593 5117 1627 5151
rect 2697 3485 2731 3519
rect 1593 3417 1627 3451
rect 12817 2601 12851 2635
rect 42625 2601 42659 2635
rect 56149 2601 56183 2635
rect 9229 2533 9263 2567
rect 29285 2533 29319 2567
rect 22845 2465 22879 2499
rect 32505 2465 32539 2499
rect 48053 2465 48087 2499
rect 3617 2397 3651 2431
rect 8769 2397 8803 2431
rect 12633 2397 12667 2431
rect 17601 2397 17635 2431
rect 22569 2397 22603 2431
rect 28917 2397 28951 2431
rect 38669 2397 38703 2431
rect 39129 2397 39163 2431
rect 42441 2397 42475 2431
rect 47593 2397 47627 2431
rect 52745 2397 52779 2431
rect 56333 2397 56367 2431
rect 2605 2329 2639 2363
rect 7573 2329 7607 2363
rect 27721 2329 27755 2363
rect 32689 2329 32723 2363
rect 37657 2329 37691 2363
rect 57253 2329 57287 2363
rect 4077 2261 4111 2295
rect 52929 2261 52963 2295
<< metal1 >>
rect 1104 57690 58880 57712
rect 1104 57638 19574 57690
rect 19626 57638 19638 57690
rect 19690 57638 19702 57690
rect 19754 57638 19766 57690
rect 19818 57638 19830 57690
rect 19882 57638 50294 57690
rect 50346 57638 50358 57690
rect 50410 57638 50422 57690
rect 50474 57638 50486 57690
rect 50538 57638 50550 57690
rect 50602 57638 58880 57690
rect 1104 57616 58880 57638
rect 44910 57468 44916 57520
rect 44968 57508 44974 57520
rect 45005 57511 45063 57517
rect 45005 57508 45017 57511
rect 44968 57480 45017 57508
rect 44968 57468 44974 57480
rect 45005 57477 45017 57480
rect 45051 57477 45063 57511
rect 45005 57471 45063 57477
rect 2777 57443 2835 57449
rect 2777 57409 2789 57443
rect 2823 57440 2835 57443
rect 2823 57412 3096 57440
rect 2823 57409 2835 57412
rect 2777 57403 2835 57409
rect 934 57332 940 57384
rect 992 57372 998 57384
rect 1581 57375 1639 57381
rect 1581 57372 1593 57375
rect 992 57344 1593 57372
rect 992 57332 998 57344
rect 1581 57341 1593 57344
rect 1627 57341 1639 57375
rect 1581 57335 1639 57341
rect 3068 57248 3096 57412
rect 45833 57375 45891 57381
rect 45833 57341 45845 57375
rect 45879 57372 45891 57375
rect 46474 57372 46480 57384
rect 45879 57344 46480 57372
rect 45879 57341 45891 57344
rect 45833 57335 45891 57341
rect 46474 57332 46480 57344
rect 46532 57332 46538 57384
rect 3050 57196 3056 57248
rect 3108 57196 3114 57248
rect 1104 57146 58880 57168
rect 1104 57094 4214 57146
rect 4266 57094 4278 57146
rect 4330 57094 4342 57146
rect 4394 57094 4406 57146
rect 4458 57094 4470 57146
rect 4522 57094 34934 57146
rect 34986 57094 34998 57146
rect 35050 57094 35062 57146
rect 35114 57094 35126 57146
rect 35178 57094 35190 57146
rect 35242 57094 58880 57146
rect 1104 57072 58880 57094
rect 1104 56602 58880 56624
rect 1104 56550 19574 56602
rect 19626 56550 19638 56602
rect 19690 56550 19702 56602
rect 19754 56550 19766 56602
rect 19818 56550 19830 56602
rect 19882 56550 50294 56602
rect 50346 56550 50358 56602
rect 50410 56550 50422 56602
rect 50474 56550 50486 56602
rect 50538 56550 50550 56602
rect 50602 56550 58880 56602
rect 1104 56528 58880 56550
rect 1104 56058 58880 56080
rect 1104 56006 4214 56058
rect 4266 56006 4278 56058
rect 4330 56006 4342 56058
rect 4394 56006 4406 56058
rect 4458 56006 4470 56058
rect 4522 56006 34934 56058
rect 34986 56006 34998 56058
rect 35050 56006 35062 56058
rect 35114 56006 35126 56058
rect 35178 56006 35190 56058
rect 35242 56006 58880 56058
rect 1104 55984 58880 56006
rect 2777 55743 2835 55749
rect 2777 55709 2789 55743
rect 2823 55709 2835 55743
rect 2777 55703 2835 55709
rect 934 55632 940 55684
rect 992 55672 998 55684
rect 1581 55675 1639 55681
rect 1581 55672 1593 55675
rect 992 55644 1593 55672
rect 992 55632 998 55644
rect 1581 55641 1593 55644
rect 1627 55641 1639 55675
rect 1581 55635 1639 55641
rect 2792 55604 2820 55703
rect 3145 55607 3203 55613
rect 3145 55604 3157 55607
rect 2792 55576 3157 55604
rect 3145 55573 3157 55576
rect 3191 55604 3203 55607
rect 15838 55604 15844 55616
rect 3191 55576 15844 55604
rect 3191 55573 3203 55576
rect 3145 55567 3203 55573
rect 15838 55564 15844 55576
rect 15896 55564 15902 55616
rect 1104 55514 58880 55536
rect 1104 55462 19574 55514
rect 19626 55462 19638 55514
rect 19690 55462 19702 55514
rect 19754 55462 19766 55514
rect 19818 55462 19830 55514
rect 19882 55462 50294 55514
rect 50346 55462 50358 55514
rect 50410 55462 50422 55514
rect 50474 55462 50486 55514
rect 50538 55462 50550 55514
rect 50602 55462 58880 55514
rect 1104 55440 58880 55462
rect 1104 54970 58880 54992
rect 1104 54918 4214 54970
rect 4266 54918 4278 54970
rect 4330 54918 4342 54970
rect 4394 54918 4406 54970
rect 4458 54918 4470 54970
rect 4522 54918 34934 54970
rect 34986 54918 34998 54970
rect 35050 54918 35062 54970
rect 35114 54918 35126 54970
rect 35178 54918 35190 54970
rect 35242 54918 58880 54970
rect 1104 54896 58880 54918
rect 1104 54426 58880 54448
rect 1104 54374 19574 54426
rect 19626 54374 19638 54426
rect 19690 54374 19702 54426
rect 19754 54374 19766 54426
rect 19818 54374 19830 54426
rect 19882 54374 50294 54426
rect 50346 54374 50358 54426
rect 50410 54374 50422 54426
rect 50474 54374 50486 54426
rect 50538 54374 50550 54426
rect 50602 54374 58880 54426
rect 1104 54352 58880 54374
rect 2777 54179 2835 54185
rect 2777 54145 2789 54179
rect 2823 54176 2835 54179
rect 2823 54148 2912 54176
rect 2823 54145 2835 54148
rect 2777 54139 2835 54145
rect 1578 54068 1584 54120
rect 1636 54068 1642 54120
rect 2884 53984 2912 54148
rect 2866 53932 2872 53984
rect 2924 53972 2930 53984
rect 3053 53975 3111 53981
rect 3053 53972 3065 53975
rect 2924 53944 3065 53972
rect 2924 53932 2930 53944
rect 3053 53941 3065 53944
rect 3099 53941 3111 53975
rect 3053 53935 3111 53941
rect 1104 53882 58880 53904
rect 1104 53830 4214 53882
rect 4266 53830 4278 53882
rect 4330 53830 4342 53882
rect 4394 53830 4406 53882
rect 4458 53830 4470 53882
rect 4522 53830 34934 53882
rect 34986 53830 34998 53882
rect 35050 53830 35062 53882
rect 35114 53830 35126 53882
rect 35178 53830 35190 53882
rect 35242 53830 58880 53882
rect 1104 53808 58880 53830
rect 1104 53338 58880 53360
rect 1104 53286 19574 53338
rect 19626 53286 19638 53338
rect 19690 53286 19702 53338
rect 19754 53286 19766 53338
rect 19818 53286 19830 53338
rect 19882 53286 50294 53338
rect 50346 53286 50358 53338
rect 50410 53286 50422 53338
rect 50474 53286 50486 53338
rect 50538 53286 50550 53338
rect 50602 53286 58880 53338
rect 1104 53264 58880 53286
rect 58529 53091 58587 53097
rect 58529 53057 58541 53091
rect 58575 53088 58587 53091
rect 58894 53088 58900 53100
rect 58575 53060 58900 53088
rect 58575 53057 58587 53060
rect 58529 53051 58587 53057
rect 58894 53048 58900 53060
rect 58952 53048 58958 53100
rect 58345 52887 58403 52893
rect 58345 52853 58357 52887
rect 58391 52884 58403 52887
rect 58986 52884 58992 52896
rect 58391 52856 58992 52884
rect 58391 52853 58403 52856
rect 58345 52847 58403 52853
rect 58986 52844 58992 52856
rect 59044 52844 59050 52896
rect 1104 52794 58880 52816
rect 1104 52742 4214 52794
rect 4266 52742 4278 52794
rect 4330 52742 4342 52794
rect 4394 52742 4406 52794
rect 4458 52742 4470 52794
rect 4522 52742 34934 52794
rect 34986 52742 34998 52794
rect 35050 52742 35062 52794
rect 35114 52742 35126 52794
rect 35178 52742 35190 52794
rect 35242 52742 58880 52794
rect 1104 52720 58880 52742
rect 58345 52683 58403 52689
rect 58345 52649 58357 52683
rect 58391 52680 58403 52683
rect 58618 52680 58624 52692
rect 58391 52652 58624 52680
rect 58391 52649 58403 52652
rect 58345 52643 58403 52649
rect 58618 52640 58624 52652
rect 58676 52640 58682 52692
rect 1578 52436 1584 52488
rect 1636 52436 1642 52488
rect 2685 52479 2743 52485
rect 2685 52445 2697 52479
rect 2731 52476 2743 52479
rect 5534 52476 5540 52488
rect 2731 52448 5540 52476
rect 2731 52445 2743 52448
rect 2685 52439 2743 52445
rect 5534 52436 5540 52448
rect 5592 52436 5598 52488
rect 58437 52411 58495 52417
rect 58437 52377 58449 52411
rect 58483 52408 58495 52411
rect 58894 52408 58900 52420
rect 58483 52380 58900 52408
rect 58483 52377 58495 52380
rect 58437 52371 58495 52377
rect 58894 52368 58900 52380
rect 58952 52368 58958 52420
rect 1104 52250 58880 52272
rect 1104 52198 19574 52250
rect 19626 52198 19638 52250
rect 19690 52198 19702 52250
rect 19754 52198 19766 52250
rect 19818 52198 19830 52250
rect 19882 52198 50294 52250
rect 50346 52198 50358 52250
rect 50410 52198 50422 52250
rect 50474 52198 50486 52250
rect 50538 52198 50550 52250
rect 50602 52198 58880 52250
rect 1104 52176 58880 52198
rect 1104 51706 58880 51728
rect 1104 51654 4214 51706
rect 4266 51654 4278 51706
rect 4330 51654 4342 51706
rect 4394 51654 4406 51706
rect 4458 51654 4470 51706
rect 4522 51654 34934 51706
rect 34986 51654 34998 51706
rect 35050 51654 35062 51706
rect 35114 51654 35126 51706
rect 35178 51654 35190 51706
rect 35242 51654 58880 51706
rect 1104 51632 58880 51654
rect 58437 51323 58495 51329
rect 58437 51289 58449 51323
rect 58483 51320 58495 51323
rect 58894 51320 58900 51332
rect 58483 51292 58900 51320
rect 58483 51289 58495 51292
rect 58437 51283 58495 51289
rect 58894 51280 58900 51292
rect 58952 51280 58958 51332
rect 58345 51255 58403 51261
rect 58345 51221 58357 51255
rect 58391 51252 58403 51255
rect 58710 51252 58716 51264
rect 58391 51224 58716 51252
rect 58391 51221 58403 51224
rect 58345 51215 58403 51221
rect 58710 51212 58716 51224
rect 58768 51212 58774 51264
rect 1104 51162 58880 51184
rect 1104 51110 19574 51162
rect 19626 51110 19638 51162
rect 19690 51110 19702 51162
rect 19754 51110 19766 51162
rect 19818 51110 19830 51162
rect 19882 51110 50294 51162
rect 50346 51110 50358 51162
rect 50410 51110 50422 51162
rect 50474 51110 50486 51162
rect 50538 51110 50550 51162
rect 50602 51110 58880 51162
rect 1104 51088 58880 51110
rect 2682 50872 2688 50924
rect 2740 50872 2746 50924
rect 934 50804 940 50856
rect 992 50844 998 50856
rect 1581 50847 1639 50853
rect 1581 50844 1593 50847
rect 992 50816 1593 50844
rect 992 50804 998 50816
rect 1581 50813 1593 50816
rect 1627 50813 1639 50847
rect 1581 50807 1639 50813
rect 1104 50618 58880 50640
rect 1104 50566 4214 50618
rect 4266 50566 4278 50618
rect 4330 50566 4342 50618
rect 4394 50566 4406 50618
rect 4458 50566 4470 50618
rect 4522 50566 34934 50618
rect 34986 50566 34998 50618
rect 35050 50566 35062 50618
rect 35114 50566 35126 50618
rect 35178 50566 35190 50618
rect 35242 50566 58880 50618
rect 1104 50544 58880 50566
rect 1104 50074 58880 50096
rect 1104 50022 19574 50074
rect 19626 50022 19638 50074
rect 19690 50022 19702 50074
rect 19754 50022 19766 50074
rect 19818 50022 19830 50074
rect 19882 50022 50294 50074
rect 50346 50022 50358 50074
rect 50410 50022 50422 50074
rect 50474 50022 50486 50074
rect 50538 50022 50550 50074
rect 50602 50022 58880 50074
rect 1104 50000 58880 50022
rect 58437 49827 58495 49833
rect 58437 49793 58449 49827
rect 58483 49824 58495 49827
rect 58483 49796 58940 49824
rect 58483 49793 58495 49796
rect 58437 49787 58495 49793
rect 58912 49768 58940 49796
rect 58253 49759 58311 49765
rect 58253 49725 58265 49759
rect 58299 49756 58311 49759
rect 58802 49756 58808 49768
rect 58299 49728 58808 49756
rect 58299 49725 58311 49728
rect 58253 49719 58311 49725
rect 58802 49716 58808 49728
rect 58860 49716 58866 49768
rect 58894 49716 58900 49768
rect 58952 49716 58958 49768
rect 1104 49530 58880 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 58880 49530
rect 1104 49456 58880 49478
rect 2222 49172 2228 49224
rect 2280 49212 2286 49224
rect 2593 49215 2651 49221
rect 2593 49212 2605 49215
rect 2280 49184 2605 49212
rect 2280 49172 2286 49184
rect 2593 49181 2605 49184
rect 2639 49181 2651 49215
rect 2593 49175 2651 49181
rect 58529 49215 58587 49221
rect 58529 49181 58541 49215
rect 58575 49212 58587 49215
rect 58575 49184 58940 49212
rect 58575 49181 58587 49184
rect 58529 49175 58587 49181
rect 934 49104 940 49156
rect 992 49144 998 49156
rect 1581 49147 1639 49153
rect 1581 49144 1593 49147
rect 992 49116 1593 49144
rect 992 49104 998 49116
rect 1581 49113 1593 49116
rect 1627 49113 1639 49147
rect 1581 49107 1639 49113
rect 58912 49088 58940 49184
rect 58342 49036 58348 49088
rect 58400 49036 58406 49088
rect 58894 49036 58900 49088
rect 58952 49036 58958 49088
rect 1104 48986 58880 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 50294 48986
rect 50346 48934 50358 48986
rect 50410 48934 50422 48986
rect 50474 48934 50486 48986
rect 50538 48934 50550 48986
rect 50602 48934 58880 48986
rect 1104 48912 58880 48934
rect 1104 48442 58880 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 58880 48442
rect 1104 48368 58880 48390
rect 58529 48127 58587 48133
rect 58529 48093 58541 48127
rect 58575 48093 58587 48127
rect 58529 48087 58587 48093
rect 58544 48056 58572 48087
rect 58894 48056 58900 48068
rect 58544 48028 58900 48056
rect 58894 48016 58900 48028
rect 58952 48016 58958 48068
rect 57790 47948 57796 48000
rect 57848 47988 57854 48000
rect 58345 47991 58403 47997
rect 58345 47988 58357 47991
rect 57848 47960 58357 47988
rect 57848 47948 57854 47960
rect 58345 47957 58357 47960
rect 58391 47957 58403 47991
rect 58345 47951 58403 47957
rect 1104 47898 58880 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 50294 47898
rect 50346 47846 50358 47898
rect 50410 47846 50422 47898
rect 50474 47846 50486 47898
rect 50538 47846 50550 47898
rect 50602 47846 58880 47898
rect 1104 47824 58880 47846
rect 2590 47608 2596 47660
rect 2648 47608 2654 47660
rect 58529 47651 58587 47657
rect 58529 47617 58541 47651
rect 58575 47648 58587 47651
rect 58894 47648 58900 47660
rect 58575 47620 58900 47648
rect 58575 47617 58587 47620
rect 58529 47611 58587 47617
rect 58894 47608 58900 47620
rect 58952 47608 58958 47660
rect 934 47540 940 47592
rect 992 47580 998 47592
rect 1581 47583 1639 47589
rect 1581 47580 1593 47583
rect 992 47552 1593 47580
rect 992 47540 998 47552
rect 1581 47549 1593 47552
rect 1627 47549 1639 47583
rect 1581 47543 1639 47549
rect 58345 47447 58403 47453
rect 58345 47413 58357 47447
rect 58391 47444 58403 47447
rect 59078 47444 59084 47456
rect 58391 47416 59084 47444
rect 58391 47413 58403 47416
rect 58345 47407 58403 47413
rect 59078 47404 59084 47416
rect 59136 47404 59142 47456
rect 1104 47354 58880 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 58880 47354
rect 1104 47280 58880 47302
rect 1104 46810 58880 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 50294 46810
rect 50346 46758 50358 46810
rect 50410 46758 50422 46810
rect 50474 46758 50486 46810
rect 50538 46758 50550 46810
rect 50602 46758 58880 46810
rect 1104 46736 58880 46758
rect 58529 46563 58587 46569
rect 58529 46529 58541 46563
rect 58575 46560 58587 46563
rect 58575 46532 58940 46560
rect 58575 46529 58587 46532
rect 58529 46523 58587 46529
rect 58912 46436 58940 46532
rect 58894 46384 58900 46436
rect 58952 46384 58958 46436
rect 58342 46316 58348 46368
rect 58400 46316 58406 46368
rect 1104 46266 58880 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 58880 46266
rect 1104 46192 58880 46214
rect 2685 45951 2743 45957
rect 2685 45917 2697 45951
rect 2731 45948 2743 45951
rect 6546 45948 6552 45960
rect 2731 45920 6552 45948
rect 2731 45917 2743 45920
rect 2685 45911 2743 45917
rect 6546 45908 6552 45920
rect 6604 45908 6610 45960
rect 57882 45908 57888 45960
rect 57940 45948 57946 45960
rect 58529 45951 58587 45957
rect 58529 45948 58541 45951
rect 57940 45920 58541 45948
rect 57940 45908 57946 45920
rect 58529 45917 58541 45920
rect 58575 45917 58587 45951
rect 58529 45911 58587 45917
rect 1578 45840 1584 45892
rect 1636 45840 1642 45892
rect 58342 45772 58348 45824
rect 58400 45772 58406 45824
rect 1104 45722 58880 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 50294 45722
rect 50346 45670 50358 45722
rect 50410 45670 50422 45722
rect 50474 45670 50486 45722
rect 50538 45670 50550 45722
rect 50602 45670 58880 45722
rect 1104 45648 58880 45670
rect 1104 45178 58880 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 58880 45178
rect 1104 45104 58880 45126
rect 58529 44863 58587 44869
rect 58529 44829 58541 44863
rect 58575 44860 58587 44863
rect 58575 44832 59032 44860
rect 58575 44829 58587 44832
rect 58529 44823 58587 44829
rect 59004 44804 59032 44832
rect 58986 44752 58992 44804
rect 59044 44752 59050 44804
rect 57514 44684 57520 44736
rect 57572 44724 57578 44736
rect 58345 44727 58403 44733
rect 58345 44724 58357 44727
rect 57572 44696 58357 44724
rect 57572 44684 57578 44696
rect 58345 44693 58357 44696
rect 58391 44693 58403 44727
rect 58345 44687 58403 44693
rect 1104 44634 58880 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 50294 44634
rect 50346 44582 50358 44634
rect 50410 44582 50422 44634
rect 50474 44582 50486 44634
rect 50538 44582 50550 44634
rect 50602 44582 58880 44634
rect 1104 44560 58880 44582
rect 2777 44387 2835 44393
rect 2777 44353 2789 44387
rect 2823 44384 2835 44387
rect 3786 44384 3792 44396
rect 2823 44356 3792 44384
rect 2823 44353 2835 44356
rect 2777 44347 2835 44353
rect 3786 44344 3792 44356
rect 3844 44344 3850 44396
rect 58529 44387 58587 44393
rect 58529 44353 58541 44387
rect 58575 44384 58587 44387
rect 58575 44356 59032 44384
rect 58575 44353 58587 44356
rect 58529 44347 58587 44353
rect 1578 44276 1584 44328
rect 1636 44276 1642 44328
rect 59004 44192 59032 44356
rect 57974 44140 57980 44192
rect 58032 44180 58038 44192
rect 58345 44183 58403 44189
rect 58345 44180 58357 44183
rect 58032 44152 58357 44180
rect 58032 44140 58038 44152
rect 58345 44149 58357 44152
rect 58391 44149 58403 44183
rect 58345 44143 58403 44149
rect 58986 44140 58992 44192
rect 59044 44140 59050 44192
rect 1104 44090 58880 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 58880 44090
rect 1104 44016 58880 44038
rect 58066 43936 58072 43988
rect 58124 43936 58130 43988
rect 58069 43843 58127 43849
rect 58069 43809 58081 43843
rect 58115 43840 58127 43843
rect 58342 43840 58348 43852
rect 58115 43812 58348 43840
rect 58115 43809 58127 43812
rect 58069 43803 58127 43809
rect 58342 43800 58348 43812
rect 58400 43800 58406 43852
rect 58161 43775 58219 43781
rect 58161 43772 58173 43775
rect 57992 43744 58173 43772
rect 57514 43664 57520 43716
rect 57572 43704 57578 43716
rect 57885 43707 57943 43713
rect 57885 43704 57897 43707
rect 57572 43676 57897 43704
rect 57572 43664 57578 43676
rect 57885 43673 57897 43676
rect 57931 43673 57943 43707
rect 57885 43667 57943 43673
rect 57992 43648 58020 43744
rect 58161 43741 58173 43744
rect 58207 43741 58219 43775
rect 58161 43735 58219 43741
rect 57974 43596 57980 43648
rect 58032 43596 58038 43648
rect 58250 43596 58256 43648
rect 58308 43636 58314 43648
rect 58345 43639 58403 43645
rect 58345 43636 58357 43639
rect 58308 43608 58357 43636
rect 58308 43596 58314 43608
rect 58345 43605 58357 43608
rect 58391 43605 58403 43639
rect 58345 43599 58403 43605
rect 1104 43546 58880 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 50294 43546
rect 50346 43494 50358 43546
rect 50410 43494 50422 43546
rect 50474 43494 50486 43546
rect 50538 43494 50550 43546
rect 50602 43494 58880 43546
rect 1104 43472 58880 43494
rect 57149 43435 57207 43441
rect 57149 43401 57161 43435
rect 57195 43432 57207 43435
rect 58066 43432 58072 43444
rect 57195 43404 58072 43432
rect 57195 43401 57207 43404
rect 57149 43395 57207 43401
rect 58066 43392 58072 43404
rect 58124 43392 58130 43444
rect 58158 43392 58164 43444
rect 58216 43392 58222 43444
rect 57790 43324 57796 43376
rect 57848 43364 57854 43376
rect 57885 43367 57943 43373
rect 57885 43364 57897 43367
rect 57848 43336 57897 43364
rect 57848 43324 57854 43336
rect 57885 43333 57897 43336
rect 57931 43333 57943 43367
rect 58176 43364 58204 43392
rect 57885 43327 57943 43333
rect 58084 43336 58204 43364
rect 58084 43305 58112 43336
rect 58069 43299 58127 43305
rect 58069 43265 58081 43299
rect 58115 43265 58127 43299
rect 58069 43259 58127 43265
rect 58161 43299 58219 43305
rect 58161 43265 58173 43299
rect 58207 43296 58219 43299
rect 59078 43296 59084 43308
rect 58207 43268 59084 43296
rect 58207 43265 58219 43268
rect 58161 43259 58219 43265
rect 59078 43256 59084 43268
rect 59136 43256 59142 43308
rect 57241 43231 57299 43237
rect 57241 43197 57253 43231
rect 57287 43197 57299 43231
rect 57241 43191 57299 43197
rect 57256 43160 57284 43191
rect 57422 43188 57428 43240
rect 57480 43188 57486 43240
rect 58434 43188 58440 43240
rect 58492 43188 58498 43240
rect 58452 43160 58480 43188
rect 57256 43132 58480 43160
rect 56321 43095 56379 43101
rect 56321 43061 56333 43095
rect 56367 43092 56379 43095
rect 56686 43092 56692 43104
rect 56367 43064 56692 43092
rect 56367 43061 56379 43064
rect 56321 43055 56379 43061
rect 56686 43052 56692 43064
rect 56744 43052 56750 43104
rect 56778 43052 56784 43104
rect 56836 43052 56842 43104
rect 58176 43101 58204 43132
rect 58802 43120 58808 43172
rect 58860 43160 58866 43172
rect 59170 43160 59176 43172
rect 58860 43132 59176 43160
rect 58860 43120 58866 43132
rect 59170 43120 59176 43132
rect 59228 43120 59234 43172
rect 58161 43095 58219 43101
rect 58161 43061 58173 43095
rect 58207 43061 58219 43095
rect 58161 43055 58219 43061
rect 58345 43095 58403 43101
rect 58345 43061 58357 43095
rect 58391 43092 58403 43095
rect 58526 43092 58532 43104
rect 58391 43064 58532 43092
rect 58391 43061 58403 43064
rect 58345 43055 58403 43061
rect 58526 43052 58532 43064
rect 58584 43052 58590 43104
rect 1104 43002 58880 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 58880 43002
rect 1104 42928 58880 42950
rect 58066 42848 58072 42900
rect 58124 42848 58130 42900
rect 58802 42848 58808 42900
rect 58860 42848 58866 42900
rect 56045 42755 56103 42761
rect 56045 42721 56057 42755
rect 56091 42752 56103 42755
rect 56686 42752 56692 42764
rect 56091 42724 56692 42752
rect 56091 42721 56103 42724
rect 56045 42715 56103 42721
rect 56686 42712 56692 42724
rect 56744 42752 56750 42764
rect 56781 42755 56839 42761
rect 56781 42752 56793 42755
rect 56744 42724 56793 42752
rect 56744 42712 56750 42724
rect 56781 42721 56793 42724
rect 56827 42752 56839 42755
rect 57054 42752 57060 42764
rect 56827 42724 57060 42752
rect 56827 42721 56839 42724
rect 56781 42715 56839 42721
rect 57054 42712 57060 42724
rect 57112 42752 57118 42764
rect 57422 42752 57428 42764
rect 57112 42724 57428 42752
rect 57112 42712 57118 42724
rect 57422 42712 57428 42724
rect 57480 42752 57486 42764
rect 57701 42755 57759 42761
rect 57701 42752 57713 42755
rect 57480 42724 57713 42752
rect 57480 42712 57486 42724
rect 57701 42721 57713 42724
rect 57747 42721 57759 42755
rect 57701 42715 57759 42721
rect 58158 42712 58164 42764
rect 58216 42712 58222 42764
rect 58820 42752 58848 42848
rect 58268 42724 58848 42752
rect 2685 42687 2743 42693
rect 2685 42653 2697 42687
rect 2731 42684 2743 42687
rect 7558 42684 7564 42696
rect 2731 42656 7564 42684
rect 2731 42653 2743 42656
rect 2685 42647 2743 42653
rect 7558 42644 7564 42656
rect 7616 42644 7622 42696
rect 56505 42687 56563 42693
rect 56505 42653 56517 42687
rect 56551 42684 56563 42687
rect 57514 42684 57520 42696
rect 56551 42656 57520 42684
rect 56551 42653 56563 42656
rect 56505 42647 56563 42653
rect 57514 42644 57520 42656
rect 57572 42644 57578 42696
rect 57609 42687 57667 42693
rect 57609 42653 57621 42687
rect 57655 42684 57667 42687
rect 58176 42684 58204 42712
rect 58268 42693 58296 42724
rect 57655 42656 58204 42684
rect 58253 42687 58311 42693
rect 57655 42653 57667 42656
rect 57609 42647 57667 42653
rect 58253 42653 58265 42687
rect 58299 42653 58311 42687
rect 58253 42647 58311 42653
rect 58342 42644 58348 42696
rect 58400 42644 58406 42696
rect 58529 42687 58587 42693
rect 58529 42653 58541 42687
rect 58575 42684 58587 42687
rect 58986 42684 58992 42696
rect 58575 42656 58992 42684
rect 58575 42653 58587 42656
rect 58529 42647 58587 42653
rect 58986 42644 58992 42656
rect 59044 42644 59050 42696
rect 934 42576 940 42628
rect 992 42616 998 42628
rect 1581 42619 1639 42625
rect 1581 42616 1593 42619
rect 992 42588 1593 42616
rect 992 42576 998 42588
rect 1581 42585 1593 42588
rect 1627 42585 1639 42619
rect 1581 42579 1639 42585
rect 55674 42576 55680 42628
rect 55732 42616 55738 42628
rect 56597 42619 56655 42625
rect 55732 42588 56180 42616
rect 55732 42576 55738 42588
rect 56152 42557 56180 42588
rect 56597 42585 56609 42619
rect 56643 42616 56655 42619
rect 57790 42616 57796 42628
rect 56643 42588 57796 42616
rect 56643 42585 56655 42588
rect 56597 42579 56655 42585
rect 57790 42576 57796 42588
rect 57848 42576 57854 42628
rect 58360 42616 58388 42644
rect 57946 42588 58388 42616
rect 56137 42551 56195 42557
rect 56137 42517 56149 42551
rect 56183 42517 56195 42551
rect 56137 42511 56195 42517
rect 56870 42508 56876 42560
rect 56928 42548 56934 42560
rect 57149 42551 57207 42557
rect 57149 42548 57161 42551
rect 56928 42520 57161 42548
rect 56928 42508 56934 42520
rect 57149 42517 57161 42520
rect 57195 42517 57207 42551
rect 57149 42511 57207 42517
rect 57517 42551 57575 42557
rect 57517 42517 57529 42551
rect 57563 42548 57575 42551
rect 57946 42548 57974 42588
rect 57563 42520 57974 42548
rect 57563 42517 57575 42520
rect 57517 42511 57575 42517
rect 58066 42508 58072 42560
rect 58124 42548 58130 42560
rect 58345 42551 58403 42557
rect 58345 42548 58357 42551
rect 58124 42520 58357 42548
rect 58124 42508 58130 42520
rect 58345 42517 58357 42520
rect 58391 42517 58403 42551
rect 58345 42511 58403 42517
rect 1104 42458 58880 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 50294 42458
rect 50346 42406 50358 42458
rect 50410 42406 50422 42458
rect 50474 42406 50486 42458
rect 50538 42406 50550 42458
rect 50602 42406 58880 42458
rect 1104 42384 58880 42406
rect 57333 42347 57391 42353
rect 57333 42313 57345 42347
rect 57379 42344 57391 42347
rect 57974 42344 57980 42356
rect 57379 42316 57980 42344
rect 57379 42313 57391 42316
rect 57333 42307 57391 42313
rect 57974 42304 57980 42316
rect 58032 42304 58038 42356
rect 59078 42304 59084 42356
rect 59136 42304 59142 42356
rect 57425 42279 57483 42285
rect 57425 42245 57437 42279
rect 57471 42276 57483 42279
rect 59096 42276 59124 42304
rect 57471 42248 59124 42276
rect 57471 42245 57483 42248
rect 57425 42239 57483 42245
rect 57517 42143 57575 42149
rect 57517 42109 57529 42143
rect 57563 42109 57575 42143
rect 57517 42103 57575 42109
rect 56873 42075 56931 42081
rect 56873 42041 56885 42075
rect 56919 42072 56931 42075
rect 57532 42072 57560 42103
rect 56919 42044 57560 42072
rect 56919 42041 56931 42044
rect 56873 42035 56931 42041
rect 57072 42016 57100 42044
rect 56962 41964 56968 42016
rect 57020 41964 57026 42016
rect 57054 41964 57060 42016
rect 57112 41964 57118 42016
rect 1104 41914 58880 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 58880 41914
rect 1104 41840 58880 41862
rect 58253 41599 58311 41605
rect 58253 41565 58265 41599
rect 58299 41565 58311 41599
rect 58253 41559 58311 41565
rect 58529 41599 58587 41605
rect 58529 41565 58541 41599
rect 58575 41596 58587 41599
rect 58575 41568 59032 41596
rect 58575 41565 58587 41568
rect 58529 41559 58587 41565
rect 58268 41528 58296 41559
rect 58802 41528 58808 41540
rect 58268 41500 58808 41528
rect 58802 41488 58808 41500
rect 58860 41488 58866 41540
rect 59004 41472 59032 41568
rect 58069 41463 58127 41469
rect 58069 41429 58081 41463
rect 58115 41460 58127 41463
rect 58158 41460 58164 41472
rect 58115 41432 58164 41460
rect 58115 41429 58127 41432
rect 58069 41423 58127 41429
rect 58158 41420 58164 41432
rect 58216 41420 58222 41472
rect 58342 41420 58348 41472
rect 58400 41420 58406 41472
rect 58986 41420 58992 41472
rect 59044 41420 59050 41472
rect 1104 41370 58880 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 50294 41370
rect 50346 41318 50358 41370
rect 50410 41318 50422 41370
rect 50474 41318 50486 41370
rect 50538 41318 50550 41370
rect 50602 41318 58880 41370
rect 1104 41296 58880 41318
rect 58158 41256 58164 41268
rect 58084 41228 58164 41256
rect 1394 41080 1400 41132
rect 1452 41080 1458 41132
rect 57885 41123 57943 41129
rect 57885 41089 57897 41123
rect 57931 41120 57943 41123
rect 57974 41120 57980 41132
rect 57931 41092 57980 41120
rect 57931 41089 57943 41092
rect 57885 41083 57943 41089
rect 57974 41080 57980 41092
rect 58032 41080 58038 41132
rect 1210 41012 1216 41064
rect 1268 41052 1274 41064
rect 1857 41055 1915 41061
rect 1857 41052 1869 41055
rect 1268 41024 1869 41052
rect 1268 41012 1274 41024
rect 1857 41021 1869 41024
rect 1903 41021 1915 41055
rect 1857 41015 1915 41021
rect 57977 40987 58035 40993
rect 57977 40953 57989 40987
rect 58023 40984 58035 40987
rect 58084 40984 58112 41228
rect 58158 41216 58164 41228
rect 58216 41216 58222 41268
rect 58250 41080 58256 41132
rect 58308 41080 58314 41132
rect 58434 41080 58440 41132
rect 58492 41080 58498 41132
rect 58158 41012 58164 41064
rect 58216 41012 58222 41064
rect 58802 40984 58808 40996
rect 58023 40956 58808 40984
rect 58023 40953 58035 40956
rect 57977 40947 58035 40953
rect 58802 40944 58808 40956
rect 58860 40944 58866 40996
rect 58066 40876 58072 40928
rect 58124 40876 58130 40928
rect 58250 40876 58256 40928
rect 58308 40876 58314 40928
rect 1104 40826 58880 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 58880 40826
rect 1104 40752 58880 40774
rect 58066 40672 58072 40724
rect 58124 40672 58130 40724
rect 58250 40672 58256 40724
rect 58308 40672 58314 40724
rect 2682 40468 2688 40520
rect 2740 40468 2746 40520
rect 58084 40517 58112 40672
rect 58268 40576 58296 40672
rect 58176 40548 58296 40576
rect 57977 40511 58035 40517
rect 57977 40477 57989 40511
rect 58023 40477 58035 40511
rect 57977 40471 58035 40477
rect 58069 40511 58127 40517
rect 58069 40477 58081 40511
rect 58115 40477 58127 40511
rect 58069 40471 58127 40477
rect 47302 40400 47308 40452
rect 47360 40440 47366 40452
rect 57609 40443 57667 40449
rect 57609 40440 57621 40443
rect 47360 40412 57621 40440
rect 47360 40400 47366 40412
rect 57609 40409 57621 40412
rect 57655 40409 57667 40443
rect 57992 40440 58020 40471
rect 58176 40440 58204 40548
rect 58253 40511 58311 40517
rect 58253 40477 58265 40511
rect 58299 40508 58311 40511
rect 58526 40508 58532 40520
rect 58299 40480 58532 40508
rect 58299 40477 58311 40480
rect 58253 40471 58311 40477
rect 58526 40468 58532 40480
rect 58584 40468 58590 40520
rect 57992 40412 58204 40440
rect 57609 40403 57667 40409
rect 2958 40332 2964 40384
rect 3016 40372 3022 40384
rect 3329 40375 3387 40381
rect 3329 40372 3341 40375
rect 3016 40344 3341 40372
rect 3016 40332 3022 40344
rect 3329 40341 3341 40344
rect 3375 40341 3387 40375
rect 3329 40335 3387 40341
rect 1104 40282 58880 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 50294 40282
rect 50346 40230 50358 40282
rect 50410 40230 50422 40282
rect 50474 40230 50486 40282
rect 50538 40230 50550 40282
rect 50602 40230 58880 40282
rect 1104 40208 58880 40230
rect 2133 40171 2191 40177
rect 2133 40137 2145 40171
rect 2179 40168 2191 40171
rect 2682 40168 2688 40180
rect 2179 40140 2688 40168
rect 2179 40137 2191 40140
rect 2133 40131 2191 40137
rect 2682 40128 2688 40140
rect 2740 40128 2746 40180
rect 8389 40171 8447 40177
rect 8389 40168 8401 40171
rect 7576 40140 8401 40168
rect 3878 40100 3884 40112
rect 1872 40072 3884 40100
rect 1394 39992 1400 40044
rect 1452 39992 1458 40044
rect 1872 40041 1900 40072
rect 3878 40060 3884 40072
rect 3936 40060 3942 40112
rect 7576 40044 7604 40140
rect 8389 40137 8401 40140
rect 8435 40137 8447 40171
rect 8389 40131 8447 40137
rect 57701 40171 57759 40177
rect 57701 40137 57713 40171
rect 57747 40137 57759 40171
rect 57701 40131 57759 40137
rect 8205 40103 8263 40109
rect 8205 40069 8217 40103
rect 8251 40100 8263 40103
rect 8294 40100 8300 40112
rect 8251 40072 8300 40100
rect 8251 40069 8263 40072
rect 8205 40063 8263 40069
rect 8294 40060 8300 40072
rect 8352 40060 8358 40112
rect 57716 40100 57744 40131
rect 57974 40128 57980 40180
rect 58032 40128 58038 40180
rect 57882 40100 57888 40112
rect 57716 40072 57888 40100
rect 57882 40060 57888 40072
rect 57940 40100 57946 40112
rect 58161 40103 58219 40109
rect 58161 40100 58173 40103
rect 57940 40072 58173 40100
rect 57940 40060 57946 40072
rect 58161 40069 58173 40072
rect 58207 40069 58219 40103
rect 58161 40063 58219 40069
rect 58342 40060 58348 40112
rect 58400 40060 58406 40112
rect 1857 40035 1915 40041
rect 1857 40001 1869 40035
rect 1903 40001 1915 40035
rect 2225 40035 2283 40041
rect 2225 40032 2237 40035
rect 1857 39995 1915 40001
rect 1964 40004 2237 40032
rect 1412 39964 1440 39992
rect 1964 39964 1992 40004
rect 2225 40001 2237 40004
rect 2271 40001 2283 40035
rect 2225 39995 2283 40001
rect 7558 39992 7564 40044
rect 7616 39992 7622 40044
rect 8386 39992 8392 40044
rect 8444 40032 8450 40044
rect 11149 40035 11207 40041
rect 8444 40018 8786 40032
rect 8444 40004 8800 40018
rect 8444 39992 8450 40004
rect 2961 39967 3019 39973
rect 1412 39936 1992 39964
rect 2133 39959 2191 39965
rect 2961 39964 2973 39967
rect 2133 39925 2145 39959
rect 2179 39956 2191 39959
rect 2240 39956 2973 39964
rect 2179 39936 2973 39956
rect 2179 39928 2268 39936
rect 2961 39933 2973 39936
rect 3007 39933 3019 39967
rect 2179 39925 2191 39928
rect 2961 39927 3019 39933
rect 2133 39919 2191 39925
rect 3510 39924 3516 39976
rect 3568 39924 3574 39976
rect 1946 39788 1952 39840
rect 2004 39788 2010 39840
rect 2869 39831 2927 39837
rect 2869 39797 2881 39831
rect 2915 39828 2927 39831
rect 3234 39828 3240 39840
rect 2915 39800 3240 39828
rect 2915 39797 2927 39800
rect 2869 39791 2927 39797
rect 3234 39788 3240 39800
rect 3292 39788 3298 39840
rect 8772 39828 8800 40004
rect 11149 40001 11161 40035
rect 11195 40032 11207 40035
rect 57517 40035 57575 40041
rect 11195 40004 11744 40032
rect 11195 40001 11207 40004
rect 11149 39995 11207 40001
rect 9858 39924 9864 39976
rect 9916 39924 9922 39976
rect 10134 39924 10140 39976
rect 10192 39924 10198 39976
rect 10321 39967 10379 39973
rect 10321 39964 10333 39967
rect 10244 39936 10333 39964
rect 10244 39828 10272 39936
rect 10321 39933 10333 39936
rect 10367 39933 10379 39967
rect 10321 39927 10379 39933
rect 11716 39840 11744 40004
rect 57517 40001 57529 40035
rect 57563 40032 57575 40035
rect 57563 40004 57836 40032
rect 57563 40001 57575 40004
rect 57517 39995 57575 40001
rect 57808 39908 57836 40004
rect 57790 39856 57796 39908
rect 57848 39856 57854 39908
rect 8772 39800 10272 39828
rect 11698 39788 11704 39840
rect 11756 39788 11762 39840
rect 1104 39738 58880 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 58880 39738
rect 1104 39664 58880 39686
rect 1394 39584 1400 39636
rect 1452 39584 1458 39636
rect 3329 39627 3387 39633
rect 3329 39593 3341 39627
rect 3375 39624 3387 39627
rect 3510 39624 3516 39636
rect 3375 39596 3516 39624
rect 3375 39593 3387 39596
rect 3329 39587 3387 39593
rect 3510 39584 3516 39596
rect 3568 39584 3574 39636
rect 9585 39627 9643 39633
rect 9585 39593 9597 39627
rect 9631 39624 9643 39627
rect 9858 39624 9864 39636
rect 9631 39596 9864 39624
rect 9631 39593 9643 39596
rect 9585 39587 9643 39593
rect 9858 39584 9864 39596
rect 9916 39584 9922 39636
rect 57425 39627 57483 39633
rect 57425 39593 57437 39627
rect 57471 39624 57483 39627
rect 58066 39624 58072 39636
rect 57471 39596 58072 39624
rect 57471 39593 57483 39596
rect 57425 39587 57483 39593
rect 58066 39584 58072 39596
rect 58124 39584 58130 39636
rect 3786 39448 3792 39500
rect 3844 39488 3850 39500
rect 5353 39491 5411 39497
rect 5353 39488 5365 39491
rect 3844 39460 5365 39488
rect 3844 39448 3850 39460
rect 5353 39457 5365 39460
rect 5399 39457 5411 39491
rect 5353 39451 5411 39457
rect 6546 39448 6552 39500
rect 6604 39448 6610 39500
rect 7929 39491 7987 39497
rect 7929 39457 7941 39491
rect 7975 39488 7987 39491
rect 8113 39491 8171 39497
rect 8113 39488 8125 39491
rect 7975 39460 8125 39488
rect 7975 39457 7987 39460
rect 7929 39451 7987 39457
rect 8113 39457 8125 39460
rect 8159 39457 8171 39491
rect 8113 39451 8171 39457
rect 57054 39448 57060 39500
rect 57112 39488 57118 39500
rect 58069 39491 58127 39497
rect 58069 39488 58081 39491
rect 57112 39460 58081 39488
rect 57112 39448 57118 39460
rect 3145 39423 3203 39429
rect 3145 39389 3157 39423
rect 3191 39389 3203 39423
rect 3145 39383 3203 39389
rect 2406 39312 2412 39364
rect 2464 39312 2470 39364
rect 2869 39355 2927 39361
rect 2869 39321 2881 39355
rect 2915 39352 2927 39355
rect 2958 39352 2964 39364
rect 2915 39324 2964 39352
rect 2915 39321 2927 39324
rect 2869 39315 2927 39321
rect 2958 39312 2964 39324
rect 3016 39312 3022 39364
rect 3160 39352 3188 39383
rect 3234 39380 3240 39432
rect 3292 39380 3298 39432
rect 3421 39423 3479 39429
rect 3421 39420 3433 39423
rect 3344 39392 3433 39420
rect 3160 39324 3280 39352
rect 3252 39296 3280 39324
rect 3344 39296 3372 39392
rect 3421 39389 3433 39392
rect 3467 39389 3479 39423
rect 3421 39383 3479 39389
rect 4614 39380 4620 39432
rect 4672 39380 4678 39432
rect 7653 39423 7711 39429
rect 7653 39389 7665 39423
rect 7699 39389 7711 39423
rect 7653 39383 7711 39389
rect 3234 39244 3240 39296
rect 3292 39244 3298 39296
rect 3326 39244 3332 39296
rect 3384 39244 3390 39296
rect 4062 39244 4068 39296
rect 4120 39244 4126 39296
rect 4798 39244 4804 39296
rect 4856 39244 4862 39296
rect 7190 39244 7196 39296
rect 7248 39244 7254 39296
rect 7668 39284 7696 39383
rect 7742 39380 7748 39432
rect 7800 39380 7806 39432
rect 8662 39380 8668 39432
rect 8720 39380 8726 39432
rect 8941 39423 8999 39429
rect 8941 39389 8953 39423
rect 8987 39389 8999 39423
rect 8941 39383 8999 39389
rect 7929 39355 7987 39361
rect 7929 39321 7941 39355
rect 7975 39352 7987 39355
rect 8956 39352 8984 39383
rect 7975 39324 8984 39352
rect 7975 39321 7987 39324
rect 7929 39315 7987 39321
rect 9122 39284 9128 39296
rect 7668 39256 9128 39284
rect 9122 39244 9128 39256
rect 9180 39244 9186 39296
rect 57164 39293 57192 39460
rect 58069 39457 58081 39460
rect 58115 39488 58127 39491
rect 58115 39460 58572 39488
rect 58115 39457 58127 39460
rect 58069 39451 58127 39457
rect 57241 39423 57299 39429
rect 57241 39389 57253 39423
rect 57287 39389 57299 39423
rect 57241 39383 57299 39389
rect 57256 39352 57284 39383
rect 57882 39380 57888 39432
rect 57940 39380 57946 39432
rect 57977 39423 58035 39429
rect 57977 39389 57989 39423
rect 58023 39420 58035 39423
rect 58158 39420 58164 39432
rect 58023 39392 58164 39420
rect 58023 39389 58035 39392
rect 57977 39383 58035 39389
rect 58158 39380 58164 39392
rect 58216 39380 58222 39432
rect 58342 39380 58348 39432
rect 58400 39380 58406 39432
rect 58544 39429 58572 39460
rect 58529 39423 58587 39429
rect 58529 39389 58541 39423
rect 58575 39389 58587 39423
rect 58529 39383 58587 39389
rect 57256 39324 58296 39352
rect 58268 39296 58296 39324
rect 57149 39287 57207 39293
rect 57149 39253 57161 39287
rect 57195 39284 57207 39287
rect 57330 39284 57336 39296
rect 57195 39256 57336 39284
rect 57195 39253 57207 39256
rect 57149 39247 57207 39253
rect 57330 39244 57336 39256
rect 57388 39244 57394 39296
rect 57517 39287 57575 39293
rect 57517 39253 57529 39287
rect 57563 39284 57575 39287
rect 57606 39284 57612 39296
rect 57563 39256 57612 39284
rect 57563 39253 57575 39256
rect 57517 39247 57575 39253
rect 57606 39244 57612 39256
rect 57664 39244 57670 39296
rect 58250 39244 58256 39296
rect 58308 39244 58314 39296
rect 58437 39287 58495 39293
rect 58437 39253 58449 39287
rect 58483 39284 58495 39287
rect 58526 39284 58532 39296
rect 58483 39256 58532 39284
rect 58483 39253 58495 39256
rect 58437 39247 58495 39253
rect 58526 39244 58532 39256
rect 58584 39244 58590 39296
rect 1104 39194 58880 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 50294 39194
rect 50346 39142 50358 39194
rect 50410 39142 50422 39194
rect 50474 39142 50486 39194
rect 50538 39142 50550 39194
rect 50602 39142 58880 39194
rect 1104 39120 58880 39142
rect 2590 39040 2596 39092
rect 2648 39040 2654 39092
rect 3786 39040 3792 39092
rect 3844 39040 3850 39092
rect 6457 39083 6515 39089
rect 4172 39052 6408 39080
rect 2608 39012 2636 39040
rect 2608 38984 2912 39012
rect 934 38904 940 38956
rect 992 38944 998 38956
rect 2884 38953 2912 38984
rect 1581 38947 1639 38953
rect 1581 38944 1593 38947
rect 992 38916 1593 38944
rect 992 38904 998 38916
rect 1581 38913 1593 38916
rect 1627 38913 1639 38947
rect 1581 38907 1639 38913
rect 2777 38947 2835 38953
rect 2777 38913 2789 38947
rect 2823 38913 2835 38947
rect 2777 38907 2835 38913
rect 2869 38947 2927 38953
rect 2869 38913 2881 38947
rect 2915 38913 2927 38947
rect 2869 38907 2927 38913
rect 2792 38876 2820 38907
rect 3694 38876 3700 38888
rect 2792 38848 3700 38876
rect 3694 38836 3700 38848
rect 3752 38836 3758 38888
rect 2406 38768 2412 38820
rect 2464 38808 2470 38820
rect 4172 38808 4200 39052
rect 6380 39012 6408 39052
rect 6457 39049 6469 39083
rect 6503 39080 6515 39083
rect 6546 39080 6552 39092
rect 6503 39052 6552 39080
rect 6503 39049 6515 39052
rect 6457 39043 6515 39049
rect 6546 39040 6552 39052
rect 6604 39040 6610 39092
rect 8202 39080 8208 39092
rect 6656 39052 8208 39080
rect 6656 39012 6684 39052
rect 8202 39040 8208 39052
rect 8260 39040 8266 39092
rect 8294 39040 8300 39092
rect 8352 39040 8358 39092
rect 8481 39083 8539 39089
rect 8481 39049 8493 39083
rect 8527 39080 8539 39083
rect 8662 39080 8668 39092
rect 8527 39052 8668 39080
rect 8527 39049 8539 39052
rect 8481 39043 8539 39049
rect 8662 39040 8668 39052
rect 8720 39040 8726 39092
rect 58066 39040 58072 39092
rect 58124 39040 58130 39092
rect 6380 38984 6762 39012
rect 8312 38953 8340 39040
rect 58084 39012 58112 39040
rect 58253 39015 58311 39021
rect 58253 39012 58265 39015
rect 58084 38984 58265 39012
rect 58253 38981 58265 38984
rect 58299 38981 58311 39015
rect 58253 38975 58311 38981
rect 8297 38947 8355 38953
rect 8297 38913 8309 38947
rect 8343 38913 8355 38947
rect 8297 38907 8355 38913
rect 8478 38904 8484 38956
rect 8536 38904 8542 38956
rect 57974 38904 57980 38956
rect 58032 38944 58038 38956
rect 58069 38947 58127 38953
rect 58069 38944 58081 38947
rect 58032 38916 58081 38944
rect 58032 38904 58038 38916
rect 58069 38913 58081 38916
rect 58115 38913 58127 38947
rect 58069 38907 58127 38913
rect 5258 38836 5264 38888
rect 5316 38836 5322 38888
rect 5534 38836 5540 38888
rect 5592 38836 5598 38888
rect 7926 38836 7932 38888
rect 7984 38836 7990 38888
rect 8205 38879 8263 38885
rect 8205 38845 8217 38879
rect 8251 38845 8263 38879
rect 8205 38839 8263 38845
rect 2464 38780 4200 38808
rect 2464 38768 2470 38780
rect 3510 38700 3516 38752
rect 3568 38700 3574 38752
rect 5552 38740 5580 38836
rect 8220 38740 8248 38839
rect 8754 38836 8760 38888
rect 8812 38876 8818 38888
rect 9401 38879 9459 38885
rect 9401 38876 9413 38879
rect 8812 38848 9413 38876
rect 8812 38836 8818 38848
rect 9401 38845 9413 38848
rect 9447 38845 9459 38879
rect 9401 38839 9459 38845
rect 58250 38808 58256 38820
rect 57624 38780 58256 38808
rect 5552 38712 8248 38740
rect 10045 38743 10103 38749
rect 10045 38709 10057 38743
rect 10091 38740 10103 38743
rect 10226 38740 10232 38752
rect 10091 38712 10232 38740
rect 10091 38709 10103 38712
rect 10045 38703 10103 38709
rect 10226 38700 10232 38712
rect 10284 38700 10290 38752
rect 57330 38700 57336 38752
rect 57388 38740 57394 38752
rect 57624 38749 57652 38780
rect 58250 38768 58256 38780
rect 58308 38768 58314 38820
rect 57609 38743 57667 38749
rect 57609 38740 57621 38743
rect 57388 38712 57621 38740
rect 57388 38700 57394 38712
rect 57609 38709 57621 38712
rect 57655 38709 57667 38743
rect 57609 38703 57667 38709
rect 58158 38700 58164 38752
rect 58216 38740 58222 38752
rect 58437 38743 58495 38749
rect 58437 38740 58449 38743
rect 58216 38712 58449 38740
rect 58216 38700 58222 38712
rect 58437 38709 58449 38712
rect 58483 38709 58495 38743
rect 58437 38703 58495 38709
rect 1104 38650 58880 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 58880 38650
rect 1104 38576 58880 38598
rect 1946 38496 1952 38548
rect 2004 38536 2010 38548
rect 2682 38536 2688 38548
rect 2004 38508 2688 38536
rect 2004 38496 2010 38508
rect 2682 38496 2688 38508
rect 2740 38496 2746 38548
rect 4062 38496 4068 38548
rect 4120 38496 4126 38548
rect 4341 38539 4399 38545
rect 4341 38505 4353 38539
rect 4387 38536 4399 38539
rect 4614 38536 4620 38548
rect 4387 38508 4620 38536
rect 4387 38505 4399 38508
rect 4341 38499 4399 38505
rect 4614 38496 4620 38508
rect 4672 38496 4678 38548
rect 5169 38539 5227 38545
rect 5169 38505 5181 38539
rect 5215 38536 5227 38539
rect 5258 38536 5264 38548
rect 5215 38508 5264 38536
rect 5215 38505 5227 38508
rect 5169 38499 5227 38505
rect 5258 38496 5264 38508
rect 5316 38496 5322 38548
rect 7561 38539 7619 38545
rect 7561 38505 7573 38539
rect 7607 38536 7619 38539
rect 7926 38536 7932 38548
rect 7607 38508 7932 38536
rect 7607 38505 7619 38508
rect 7561 38499 7619 38505
rect 7926 38496 7932 38508
rect 7984 38496 7990 38548
rect 8386 38496 8392 38548
rect 8444 38496 8450 38548
rect 4080 38409 4108 38496
rect 5721 38471 5779 38477
rect 5721 38468 5733 38471
rect 4172 38440 5733 38468
rect 2133 38403 2191 38409
rect 2133 38369 2145 38403
rect 2179 38400 2191 38403
rect 2961 38403 3019 38409
rect 2961 38400 2973 38403
rect 2179 38372 2973 38400
rect 2179 38369 2191 38372
rect 2133 38363 2191 38369
rect 2961 38369 2973 38372
rect 3007 38369 3019 38403
rect 3881 38403 3939 38409
rect 3881 38400 3893 38403
rect 2961 38363 3019 38369
rect 3344 38372 3893 38400
rect 1854 38292 1860 38344
rect 1912 38292 1918 38344
rect 2225 38335 2283 38341
rect 2225 38332 2237 38335
rect 2148 38304 2237 38332
rect 2148 38273 2176 38304
rect 2225 38301 2237 38304
rect 2271 38301 2283 38335
rect 2225 38295 2283 38301
rect 2682 38292 2688 38344
rect 2740 38332 2746 38344
rect 3344 38332 3372 38372
rect 3881 38369 3893 38372
rect 3927 38369 3939 38403
rect 3881 38363 3939 38369
rect 4065 38403 4123 38409
rect 4065 38369 4077 38403
rect 4111 38369 4123 38403
rect 4065 38363 4123 38369
rect 2740 38304 3372 38332
rect 2740 38292 2746 38304
rect 3418 38292 3424 38344
rect 3476 38332 3482 38344
rect 3513 38335 3571 38341
rect 3513 38332 3525 38335
rect 3476 38304 3525 38332
rect 3476 38292 3482 38304
rect 3513 38301 3525 38304
rect 3559 38301 3571 38335
rect 3513 38295 3571 38301
rect 3786 38292 3792 38344
rect 3844 38292 3850 38344
rect 3896 38332 3924 38363
rect 4172 38332 4200 38440
rect 5721 38437 5733 38440
rect 5767 38468 5779 38471
rect 7742 38468 7748 38480
rect 5767 38440 7748 38468
rect 5767 38437 5779 38440
rect 5721 38431 5779 38437
rect 7742 38428 7748 38440
rect 7800 38468 7806 38480
rect 7837 38471 7895 38477
rect 7837 38468 7849 38471
rect 7800 38440 7849 38468
rect 7800 38428 7806 38440
rect 7837 38437 7849 38440
rect 7883 38437 7895 38471
rect 7837 38431 7895 38437
rect 4525 38403 4583 38409
rect 4525 38400 4537 38403
rect 4356 38372 4537 38400
rect 3896 38304 4200 38332
rect 4246 38292 4252 38344
rect 4304 38292 4310 38344
rect 2133 38267 2191 38273
rect 2133 38233 2145 38267
rect 2179 38233 2191 38267
rect 2133 38227 2191 38233
rect 2498 38224 2504 38276
rect 2556 38264 2562 38276
rect 4065 38267 4123 38273
rect 2556 38236 4016 38264
rect 2556 38224 2562 38236
rect 2866 38156 2872 38208
rect 2924 38156 2930 38208
rect 3988 38196 4016 38236
rect 4065 38233 4077 38267
rect 4111 38264 4123 38267
rect 4356 38264 4384 38372
rect 4525 38369 4537 38372
rect 4571 38369 4583 38403
rect 4525 38363 4583 38369
rect 5905 38403 5963 38409
rect 5905 38369 5917 38403
rect 5951 38400 5963 38403
rect 6181 38403 6239 38409
rect 6181 38400 6193 38403
rect 5951 38372 6193 38400
rect 5951 38369 5963 38372
rect 5905 38363 5963 38369
rect 6181 38369 6193 38372
rect 6227 38369 6239 38403
rect 6181 38363 6239 38369
rect 6825 38403 6883 38409
rect 6825 38369 6837 38403
rect 6871 38400 6883 38403
rect 7466 38400 7472 38412
rect 6871 38372 7472 38400
rect 6871 38369 6883 38372
rect 6825 38363 6883 38369
rect 7466 38360 7472 38372
rect 7524 38360 7530 38412
rect 8021 38403 8079 38409
rect 8021 38369 8033 38403
rect 8067 38400 8079 38403
rect 8113 38403 8171 38409
rect 8113 38400 8125 38403
rect 8067 38372 8125 38400
rect 8067 38369 8079 38372
rect 8021 38363 8079 38369
rect 8113 38369 8125 38372
rect 8159 38369 8171 38403
rect 8404 38400 8432 38496
rect 57238 38428 57244 38480
rect 57296 38468 57302 38480
rect 57609 38471 57667 38477
rect 57609 38468 57621 38471
rect 57296 38440 57621 38468
rect 57296 38428 57302 38440
rect 57609 38437 57621 38440
rect 57655 38437 57667 38471
rect 58802 38468 58808 38480
rect 57609 38431 57667 38437
rect 58084 38440 58808 38468
rect 8404 38372 9444 38400
rect 8113 38363 8171 38369
rect 4433 38335 4491 38341
rect 4433 38301 4445 38335
rect 4479 38301 4491 38335
rect 4433 38295 4491 38301
rect 4111 38236 4384 38264
rect 4448 38264 4476 38295
rect 4798 38292 4804 38344
rect 4856 38292 4862 38344
rect 5626 38292 5632 38344
rect 5684 38292 5690 38344
rect 6917 38335 6975 38341
rect 6917 38301 6929 38335
rect 6963 38301 6975 38335
rect 6917 38295 6975 38301
rect 4816 38264 4844 38292
rect 4448 38236 4844 38264
rect 5905 38267 5963 38273
rect 4111 38233 4123 38236
rect 4065 38227 4123 38233
rect 5905 38233 5917 38267
rect 5951 38264 5963 38267
rect 6932 38264 6960 38295
rect 7742 38292 7748 38344
rect 7800 38292 7806 38344
rect 8662 38292 8668 38344
rect 8720 38292 8726 38344
rect 8754 38292 8760 38344
rect 8812 38292 8818 38344
rect 9416 38332 9444 38372
rect 10502 38360 10508 38412
rect 10560 38400 10566 38412
rect 58084 38409 58112 38440
rect 58802 38428 58808 38440
rect 58860 38428 58866 38480
rect 10781 38403 10839 38409
rect 10781 38400 10793 38403
rect 10560 38372 10793 38400
rect 10560 38360 10566 38372
rect 10781 38369 10793 38372
rect 10827 38400 10839 38403
rect 11057 38403 11115 38409
rect 11057 38400 11069 38403
rect 10827 38372 11069 38400
rect 10827 38369 10839 38372
rect 10781 38363 10839 38369
rect 11057 38369 11069 38372
rect 11103 38369 11115 38403
rect 11057 38363 11115 38369
rect 58069 38403 58127 38409
rect 58069 38369 58081 38403
rect 58115 38369 58127 38403
rect 58069 38363 58127 38369
rect 58250 38360 58256 38412
rect 58308 38360 58314 38412
rect 9490 38332 9496 38344
rect 9416 38318 9496 38332
rect 9430 38304 9496 38318
rect 9490 38292 9496 38304
rect 9548 38292 9554 38344
rect 57333 38335 57391 38341
rect 57333 38301 57345 38335
rect 57379 38332 57391 38335
rect 57379 38304 58388 38332
rect 57379 38301 57391 38304
rect 57333 38295 57391 38301
rect 5951 38236 6960 38264
rect 8021 38267 8079 38273
rect 5951 38233 5963 38236
rect 5905 38227 5963 38233
rect 8021 38233 8033 38267
rect 8067 38264 8079 38267
rect 8772 38264 8800 38292
rect 58360 38276 58388 38304
rect 8067 38236 8800 38264
rect 8067 38233 8079 38236
rect 8021 38227 8079 38233
rect 10226 38224 10232 38276
rect 10284 38264 10290 38276
rect 10505 38267 10563 38273
rect 10505 38264 10517 38267
rect 10284 38236 10517 38264
rect 10284 38224 10290 38236
rect 10505 38233 10517 38236
rect 10551 38233 10563 38267
rect 57974 38264 57980 38276
rect 10505 38227 10563 38233
rect 57532 38236 57980 38264
rect 9030 38196 9036 38208
rect 3988 38168 9036 38196
rect 9030 38156 9036 38168
rect 9088 38156 9094 38208
rect 57241 38199 57299 38205
rect 57241 38165 57253 38199
rect 57287 38196 57299 38199
rect 57330 38196 57336 38208
rect 57287 38168 57336 38196
rect 57287 38165 57299 38168
rect 57241 38159 57299 38165
rect 57330 38156 57336 38168
rect 57388 38156 57394 38208
rect 57532 38205 57560 38236
rect 57974 38224 57980 38236
rect 58032 38224 58038 38276
rect 58342 38224 58348 38276
rect 58400 38224 58406 38276
rect 57517 38199 57575 38205
rect 57517 38165 57529 38199
rect 57563 38165 57575 38199
rect 57517 38159 57575 38165
rect 1104 38106 58880 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 50294 38106
rect 50346 38054 50358 38106
rect 50410 38054 50422 38106
rect 50474 38054 50486 38106
rect 50538 38054 50550 38106
rect 50602 38054 58880 38106
rect 1104 38032 58880 38054
rect 1489 37995 1547 38001
rect 1489 37961 1501 37995
rect 1535 37992 1547 37995
rect 2590 37992 2596 38004
rect 1535 37964 2596 37992
rect 1535 37961 1547 37964
rect 1489 37955 1547 37961
rect 2590 37952 2596 37964
rect 2648 37952 2654 38004
rect 2866 37952 2872 38004
rect 2924 37992 2930 38004
rect 2924 37964 3004 37992
rect 2924 37952 2930 37964
rect 2406 37884 2412 37936
rect 2464 37884 2470 37936
rect 2976 37933 3004 37964
rect 3418 37952 3424 38004
rect 3476 37952 3482 38004
rect 3510 37952 3516 38004
rect 3568 37952 3574 38004
rect 7190 37952 7196 38004
rect 7248 37952 7254 38004
rect 7466 37952 7472 38004
rect 7524 37952 7530 38004
rect 8481 37995 8539 38001
rect 8481 37961 8493 37995
rect 8527 37992 8539 37995
rect 8662 37992 8668 38004
rect 8527 37964 8668 37992
rect 8527 37961 8539 37964
rect 8481 37955 8539 37961
rect 8662 37952 8668 37964
rect 8720 37952 8726 38004
rect 9030 37952 9036 38004
rect 9088 37952 9094 38004
rect 58434 37952 58440 38004
rect 58492 37952 58498 38004
rect 2961 37927 3019 37933
rect 2961 37893 2973 37927
rect 3007 37893 3019 37927
rect 2961 37887 3019 37893
rect 3326 37816 3332 37868
rect 3384 37816 3390 37868
rect 3528 37865 3556 37952
rect 3513 37859 3571 37865
rect 3513 37825 3525 37859
rect 3559 37825 3571 37859
rect 3513 37819 3571 37825
rect 4246 37816 4252 37868
rect 4304 37856 4310 37868
rect 4304 37828 4743 37856
rect 4304 37816 4310 37828
rect 2958 37748 2964 37800
rect 3016 37788 3022 37800
rect 3016 37760 3188 37788
rect 3016 37748 3022 37760
rect 3160 37720 3188 37760
rect 3234 37748 3240 37800
rect 3292 37748 3298 37800
rect 3344 37788 3372 37816
rect 4264 37788 4292 37816
rect 3344 37760 4292 37788
rect 4614 37748 4620 37800
rect 4672 37748 4678 37800
rect 4715 37788 4743 37828
rect 5718 37816 5724 37868
rect 5776 37856 5782 37868
rect 6641 37859 6699 37865
rect 6641 37856 6653 37859
rect 5776 37828 6653 37856
rect 5776 37816 5782 37828
rect 6641 37825 6653 37828
rect 6687 37825 6699 37859
rect 7208 37856 7236 37952
rect 8386 37865 8392 37868
rect 7377 37859 7435 37865
rect 7377 37856 7389 37859
rect 7208 37828 7389 37856
rect 6641 37819 6699 37825
rect 7377 37825 7389 37828
rect 7423 37825 7435 37859
rect 7377 37819 7435 37825
rect 7561 37859 7619 37865
rect 7561 37825 7573 37859
rect 7607 37856 7619 37859
rect 8381 37856 8392 37865
rect 7607 37828 8392 37856
rect 7607 37825 7619 37828
rect 7561 37819 7619 37825
rect 8381 37819 8392 37828
rect 7576 37788 7604 37819
rect 8386 37816 8392 37819
rect 8444 37816 8450 37868
rect 8573 37859 8631 37865
rect 8573 37825 8585 37859
rect 8619 37856 8631 37859
rect 8849 37859 8907 37865
rect 8849 37856 8861 37859
rect 8619 37828 8861 37856
rect 8619 37825 8631 37828
rect 8573 37819 8631 37825
rect 8849 37825 8861 37828
rect 8895 37825 8907 37859
rect 9048 37856 9076 37952
rect 59170 37924 59176 37936
rect 57900 37896 59176 37924
rect 57900 37865 57928 37896
rect 59170 37884 59176 37896
rect 59228 37884 59234 37936
rect 9401 37859 9459 37865
rect 9401 37856 9413 37859
rect 9048 37828 9413 37856
rect 8849 37819 8907 37825
rect 9401 37825 9413 37828
rect 9447 37825 9459 37859
rect 57885 37859 57943 37865
rect 57885 37856 57897 37859
rect 9401 37819 9459 37825
rect 57624 37828 57897 37856
rect 4715 37760 7604 37788
rect 8662 37720 8668 37732
rect 3160 37692 8668 37720
rect 8662 37680 8668 37692
rect 8720 37680 8726 37732
rect 4062 37612 4068 37664
rect 4120 37612 4126 37664
rect 7282 37612 7288 37664
rect 7340 37612 7346 37664
rect 56778 37612 56784 37664
rect 56836 37652 56842 37664
rect 57624 37661 57652 37828
rect 57885 37825 57897 37828
rect 57931 37825 57943 37859
rect 57885 37819 57943 37825
rect 58250 37816 58256 37868
rect 58308 37816 58314 37868
rect 57609 37655 57667 37661
rect 57609 37652 57621 37655
rect 56836 37624 57621 37652
rect 56836 37612 56842 37624
rect 57609 37621 57621 37624
rect 57655 37621 57667 37655
rect 57609 37615 57667 37621
rect 58158 37612 58164 37664
rect 58216 37612 58222 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 5629 37451 5687 37457
rect 5629 37417 5641 37451
rect 5675 37448 5687 37451
rect 5718 37448 5724 37460
rect 5675 37420 5724 37448
rect 5675 37417 5687 37420
rect 5629 37411 5687 37417
rect 5718 37408 5724 37420
rect 5776 37408 5782 37460
rect 7282 37408 7288 37460
rect 7340 37408 7346 37460
rect 8662 37408 8668 37460
rect 8720 37408 8726 37460
rect 58250 37408 58256 37460
rect 58308 37448 58314 37460
rect 58345 37451 58403 37457
rect 58345 37448 58357 37451
rect 58308 37420 58357 37448
rect 58308 37408 58314 37420
rect 58345 37417 58357 37420
rect 58391 37417 58403 37451
rect 58345 37411 58403 37417
rect 7300 37380 7328 37408
rect 7300 37352 8248 37380
rect 3326 37272 3332 37324
rect 3384 37312 3390 37324
rect 3384 37284 3464 37312
rect 3384 37272 3390 37284
rect 1578 37204 1584 37256
rect 1636 37204 1642 37256
rect 2774 37204 2780 37256
rect 2832 37204 2838 37256
rect 3436 37253 3464 37284
rect 3694 37272 3700 37324
rect 3752 37312 3758 37324
rect 7101 37315 7159 37321
rect 3752 37284 4016 37312
rect 3752 37272 3758 37284
rect 3421 37247 3479 37253
rect 3421 37213 3433 37247
rect 3467 37213 3479 37247
rect 3421 37207 3479 37213
rect 3605 37247 3663 37253
rect 3605 37213 3617 37247
rect 3651 37244 3663 37247
rect 3881 37247 3939 37253
rect 3881 37244 3893 37247
rect 3651 37216 3893 37244
rect 3651 37213 3663 37216
rect 3605 37207 3663 37213
rect 3881 37213 3893 37216
rect 3927 37213 3939 37247
rect 3988 37244 4016 37284
rect 7101 37281 7113 37315
rect 7147 37312 7159 37315
rect 7650 37312 7656 37324
rect 7147 37284 7656 37312
rect 7147 37281 7159 37284
rect 7101 37275 7159 37281
rect 7650 37272 7656 37284
rect 7708 37272 7714 37324
rect 8220 37253 8248 37352
rect 8680 37312 8708 37408
rect 9493 37315 9551 37321
rect 9493 37312 9505 37315
rect 8680 37284 9505 37312
rect 9493 37281 9505 37284
rect 9539 37281 9551 37315
rect 58894 37312 58900 37324
rect 9493 37275 9551 37281
rect 58544 37284 58900 37312
rect 4433 37247 4491 37253
rect 4433 37244 4445 37247
rect 3988 37216 4445 37244
rect 3881 37207 3939 37213
rect 4433 37213 4445 37216
rect 4479 37213 4491 37247
rect 4433 37207 4491 37213
rect 4617 37247 4675 37253
rect 4617 37213 4629 37247
rect 4663 37213 4675 37247
rect 4617 37207 4675 37213
rect 7377 37247 7435 37253
rect 7377 37213 7389 37247
rect 7423 37213 7435 37247
rect 7377 37207 7435 37213
rect 8113 37247 8171 37253
rect 8113 37213 8125 37247
rect 8159 37213 8171 37247
rect 8113 37207 8171 37213
rect 8205 37247 8263 37253
rect 8205 37213 8217 37247
rect 8251 37213 8263 37247
rect 8205 37207 8263 37213
rect 3970 37136 3976 37188
rect 4028 37176 4034 37188
rect 4632 37176 4660 37207
rect 4028 37148 4660 37176
rect 4028 37136 4034 37148
rect 6086 37136 6092 37188
rect 6144 37136 6150 37188
rect 3513 37111 3571 37117
rect 3513 37077 3525 37111
rect 3559 37108 3571 37111
rect 4614 37108 4620 37120
rect 3559 37080 4620 37108
rect 3559 37077 3571 37080
rect 3513 37071 3571 37077
rect 4614 37068 4620 37080
rect 4672 37068 4678 37120
rect 5261 37111 5319 37117
rect 5261 37077 5273 37111
rect 5307 37108 5319 37111
rect 5350 37108 5356 37120
rect 5307 37080 5356 37108
rect 5307 37077 5319 37080
rect 5261 37071 5319 37077
rect 5350 37068 5356 37080
rect 5408 37068 5414 37120
rect 5534 37068 5540 37120
rect 5592 37108 5598 37120
rect 5718 37108 5724 37120
rect 5592 37080 5724 37108
rect 5592 37068 5598 37080
rect 5718 37068 5724 37080
rect 5776 37108 5782 37120
rect 7392 37108 7420 37207
rect 8128 37176 8156 37207
rect 8386 37204 8392 37256
rect 8444 37244 8450 37256
rect 58544 37253 58572 37284
rect 58894 37272 58900 37284
rect 58952 37272 58958 37324
rect 58529 37247 58587 37253
rect 8444 37216 8800 37244
rect 8444 37204 8450 37216
rect 8297 37179 8355 37185
rect 8297 37176 8309 37179
rect 8128 37148 8309 37176
rect 8297 37145 8309 37148
rect 8343 37145 8355 37179
rect 8297 37139 8355 37145
rect 8772 37120 8800 37216
rect 58529 37213 58541 37247
rect 58575 37213 58587 37247
rect 58529 37207 58587 37213
rect 5776 37080 7420 37108
rect 5776 37068 5782 37080
rect 7466 37068 7472 37120
rect 7524 37068 7530 37120
rect 8754 37068 8760 37120
rect 8812 37068 8818 37120
rect 8938 37068 8944 37120
rect 8996 37068 9002 37120
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 7466 36864 7472 36916
rect 7524 36864 7530 36916
rect 7650 36864 7656 36916
rect 7708 36864 7714 36916
rect 58250 36864 58256 36916
rect 58308 36864 58314 36916
rect 2225 36839 2283 36845
rect 2225 36805 2237 36839
rect 2271 36805 2283 36839
rect 2225 36799 2283 36805
rect 1949 36771 2007 36777
rect 1949 36737 1961 36771
rect 1995 36737 2007 36771
rect 2240 36768 2268 36799
rect 2406 36796 2412 36848
rect 2464 36836 2470 36848
rect 2464 36808 2774 36836
rect 2464 36796 2470 36808
rect 2317 36771 2375 36777
rect 2317 36768 2329 36771
rect 2240 36740 2329 36768
rect 1949 36731 2007 36737
rect 2317 36737 2329 36740
rect 2363 36737 2375 36771
rect 2746 36768 2774 36808
rect 5350 36796 5356 36848
rect 5408 36836 5414 36848
rect 5445 36839 5503 36845
rect 5445 36836 5457 36839
rect 5408 36808 5457 36836
rect 5408 36796 5414 36808
rect 5445 36805 5457 36808
rect 5491 36805 5503 36839
rect 5445 36799 5503 36805
rect 6917 36839 6975 36845
rect 6917 36805 6929 36839
rect 6963 36836 6975 36839
rect 6963 36808 7052 36836
rect 6963 36805 6975 36808
rect 6917 36799 6975 36805
rect 2746 36754 4370 36768
rect 2746 36740 4384 36754
rect 2317 36731 2375 36737
rect 1964 36632 1992 36731
rect 2225 36703 2283 36709
rect 2225 36669 2237 36703
rect 2271 36700 2283 36703
rect 3053 36703 3111 36709
rect 3053 36700 3065 36703
rect 2271 36672 3065 36700
rect 2271 36669 2283 36672
rect 2225 36663 2283 36669
rect 3053 36669 3065 36672
rect 3099 36669 3111 36703
rect 3053 36663 3111 36669
rect 3602 36660 3608 36712
rect 3660 36660 3666 36712
rect 3694 36660 3700 36712
rect 3752 36700 3758 36712
rect 3973 36703 4031 36709
rect 3973 36700 3985 36703
rect 3752 36672 3985 36700
rect 3752 36660 3758 36672
rect 3973 36669 3985 36672
rect 4019 36669 4031 36703
rect 4356 36700 4384 36740
rect 5718 36728 5724 36780
rect 5776 36728 5782 36780
rect 6086 36728 6092 36780
rect 6144 36728 6150 36780
rect 7024 36777 7052 36808
rect 6641 36771 6699 36777
rect 6641 36737 6653 36771
rect 6687 36737 6699 36771
rect 6641 36731 6699 36737
rect 7009 36771 7067 36777
rect 7009 36737 7021 36771
rect 7055 36737 7067 36771
rect 7009 36731 7067 36737
rect 6104 36700 6132 36728
rect 4356 36672 6132 36700
rect 3973 36663 4031 36669
rect 3326 36632 3332 36644
rect 1964 36604 3332 36632
rect 3326 36592 3332 36604
rect 3384 36592 3390 36644
rect 6656 36632 6684 36731
rect 6917 36703 6975 36709
rect 6917 36669 6929 36703
rect 6963 36700 6975 36703
rect 7484 36700 7512 36864
rect 8481 36839 8539 36845
rect 8481 36805 8493 36839
rect 8527 36836 8539 36839
rect 8662 36836 8668 36848
rect 8527 36808 8668 36836
rect 8527 36805 8539 36808
rect 8481 36799 8539 36805
rect 8662 36796 8668 36808
rect 8720 36796 8726 36848
rect 9490 36796 9496 36848
rect 9548 36796 9554 36848
rect 10502 36728 10508 36780
rect 10560 36768 10566 36780
rect 10781 36771 10839 36777
rect 10781 36768 10793 36771
rect 10560 36740 10793 36768
rect 10560 36728 10566 36740
rect 10781 36737 10793 36740
rect 10827 36737 10839 36771
rect 57885 36771 57943 36777
rect 57885 36768 57897 36771
rect 10781 36731 10839 36737
rect 57716 36740 57897 36768
rect 6963 36672 7512 36700
rect 6963 36669 6975 36672
rect 6917 36663 6975 36669
rect 8386 36660 8392 36712
rect 8444 36660 8450 36712
rect 10226 36660 10232 36712
rect 10284 36660 10290 36712
rect 7006 36632 7012 36644
rect 6656 36604 7012 36632
rect 7006 36592 7012 36604
rect 7064 36592 7070 36644
rect 57716 36576 57744 36740
rect 57885 36737 57897 36740
rect 57931 36737 57943 36771
rect 57885 36731 57943 36737
rect 58069 36771 58127 36777
rect 58069 36737 58081 36771
rect 58115 36768 58127 36771
rect 58268 36768 58296 36864
rect 58115 36740 58296 36768
rect 58529 36771 58587 36777
rect 58115 36737 58127 36740
rect 58069 36731 58127 36737
rect 58529 36737 58541 36771
rect 58575 36768 58587 36771
rect 58575 36740 58940 36768
rect 58575 36737 58587 36740
rect 58529 36731 58587 36737
rect 58912 36644 58940 36740
rect 58894 36592 58900 36644
rect 58952 36592 58958 36644
rect 2041 36567 2099 36573
rect 2041 36533 2053 36567
rect 2087 36564 2099 36567
rect 2682 36564 2688 36576
rect 2087 36536 2688 36564
rect 2087 36533 2099 36536
rect 2041 36527 2099 36533
rect 2682 36524 2688 36536
rect 2740 36524 2746 36576
rect 2866 36524 2872 36576
rect 2924 36564 2930 36576
rect 2961 36567 3019 36573
rect 2961 36564 2973 36567
rect 2924 36536 2973 36564
rect 2924 36524 2930 36536
rect 2961 36533 2973 36536
rect 3007 36533 3019 36567
rect 2961 36527 3019 36533
rect 6733 36567 6791 36573
rect 6733 36533 6745 36567
rect 6779 36564 6791 36567
rect 7282 36564 7288 36576
rect 6779 36536 7288 36564
rect 6779 36533 6791 36536
rect 6733 36527 6791 36533
rect 7282 36524 7288 36536
rect 7340 36524 7346 36576
rect 7745 36567 7803 36573
rect 7745 36533 7757 36567
rect 7791 36564 7803 36567
rect 8202 36564 8208 36576
rect 7791 36536 8208 36564
rect 7791 36533 7803 36536
rect 7745 36527 7803 36533
rect 8202 36524 8208 36536
rect 8260 36524 8266 36576
rect 57698 36524 57704 36576
rect 57756 36524 57762 36576
rect 57974 36524 57980 36576
rect 58032 36524 58038 36576
rect 58158 36524 58164 36576
rect 58216 36564 58222 36576
rect 58345 36567 58403 36573
rect 58345 36564 58357 36567
rect 58216 36536 58357 36564
rect 58216 36524 58222 36536
rect 58345 36533 58357 36536
rect 58391 36533 58403 36567
rect 58345 36527 58403 36533
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 1397 36363 1455 36369
rect 1397 36329 1409 36363
rect 1443 36360 1455 36363
rect 2774 36360 2780 36372
rect 1443 36332 2780 36360
rect 1443 36329 1455 36332
rect 1397 36323 1455 36329
rect 2774 36320 2780 36332
rect 2832 36320 2838 36372
rect 3329 36363 3387 36369
rect 3329 36329 3341 36363
rect 3375 36360 3387 36363
rect 3602 36360 3608 36372
rect 3375 36332 3608 36360
rect 3375 36329 3387 36332
rect 3329 36323 3387 36329
rect 3602 36320 3608 36332
rect 3660 36320 3666 36372
rect 3970 36320 3976 36372
rect 4028 36320 4034 36372
rect 4062 36320 4068 36372
rect 4120 36320 4126 36372
rect 8202 36320 8208 36372
rect 8260 36320 8266 36372
rect 8386 36320 8392 36372
rect 8444 36360 8450 36372
rect 8573 36363 8631 36369
rect 8573 36360 8585 36363
rect 8444 36332 8585 36360
rect 8444 36320 8450 36332
rect 8573 36329 8585 36332
rect 8619 36329 8631 36363
rect 8573 36323 8631 36329
rect 8938 36320 8944 36372
rect 8996 36320 9002 36372
rect 9953 36363 10011 36369
rect 9953 36329 9965 36363
rect 9999 36360 10011 36363
rect 10226 36360 10232 36372
rect 9999 36332 10232 36360
rect 9999 36329 10011 36332
rect 9953 36323 10011 36329
rect 10226 36320 10232 36332
rect 10284 36320 10290 36372
rect 57974 36320 57980 36372
rect 58032 36320 58038 36372
rect 58526 36320 58532 36372
rect 58584 36320 58590 36372
rect 3234 36252 3240 36304
rect 3292 36252 3298 36304
rect 2866 36184 2872 36236
rect 2924 36184 2930 36236
rect 3145 36227 3203 36233
rect 3145 36193 3157 36227
rect 3191 36193 3203 36227
rect 3145 36187 3203 36193
rect 3160 36100 3188 36187
rect 3252 36175 3280 36252
rect 4080 36233 4108 36320
rect 4065 36227 4123 36233
rect 4065 36193 4077 36227
rect 4111 36193 4123 36227
rect 8113 36227 8171 36233
rect 8113 36224 8125 36227
rect 4065 36187 4123 36193
rect 7300 36196 8125 36224
rect 3237 36169 3295 36175
rect 3237 36135 3249 36169
rect 3283 36135 3295 36169
rect 7300 36168 7328 36196
rect 8113 36193 8125 36196
rect 8159 36193 8171 36227
rect 8220 36224 8248 36320
rect 8297 36227 8355 36233
rect 8297 36224 8309 36227
rect 8220 36196 8309 36224
rect 8113 36187 8171 36193
rect 8297 36193 8309 36196
rect 8343 36193 8355 36227
rect 8754 36224 8760 36236
rect 8297 36187 8355 36193
rect 8496 36196 8760 36224
rect 3237 36129 3295 36135
rect 3418 36116 3424 36168
rect 3476 36116 3482 36168
rect 3789 36159 3847 36165
rect 3789 36125 3801 36159
rect 3835 36125 3847 36159
rect 3789 36119 3847 36125
rect 3881 36159 3939 36165
rect 3881 36125 3893 36159
rect 3927 36156 3939 36159
rect 3970 36156 3976 36168
rect 3927 36128 3976 36156
rect 3927 36125 3939 36128
rect 3881 36119 3939 36125
rect 2406 36048 2412 36100
rect 2464 36048 2470 36100
rect 3142 36048 3148 36100
rect 3200 36048 3206 36100
rect 3804 36088 3832 36119
rect 3970 36116 3976 36128
rect 4028 36116 4034 36168
rect 4522 36116 4528 36168
rect 4580 36116 4586 36168
rect 7193 36159 7251 36165
rect 7193 36156 7205 36159
rect 6472 36128 7205 36156
rect 6472 36100 6500 36128
rect 7193 36125 7205 36128
rect 7239 36125 7251 36159
rect 7193 36119 7251 36125
rect 7282 36116 7288 36168
rect 7340 36116 7346 36168
rect 8021 36159 8079 36165
rect 8021 36125 8033 36159
rect 8067 36156 8079 36159
rect 8386 36156 8392 36168
rect 8067 36128 8392 36156
rect 8067 36125 8079 36128
rect 8021 36119 8079 36125
rect 8386 36116 8392 36128
rect 8444 36116 8450 36168
rect 8496 36165 8524 36196
rect 8754 36184 8760 36196
rect 8812 36184 8818 36236
rect 8481 36159 8539 36165
rect 8481 36125 8493 36159
rect 8527 36125 8539 36159
rect 8481 36119 8539 36125
rect 8665 36159 8723 36165
rect 8665 36125 8677 36159
rect 8711 36156 8723 36159
rect 8956 36156 8984 36320
rect 57514 36252 57520 36304
rect 57572 36252 57578 36304
rect 57992 36224 58020 36320
rect 58544 36224 58572 36320
rect 57716 36196 58020 36224
rect 58084 36196 58572 36224
rect 57716 36165 57744 36196
rect 8711 36128 8984 36156
rect 9309 36159 9367 36165
rect 8711 36125 8723 36128
rect 8665 36119 8723 36125
rect 9309 36125 9321 36159
rect 9355 36125 9367 36159
rect 9309 36119 9367 36125
rect 57701 36159 57759 36165
rect 57701 36125 57713 36159
rect 57747 36125 57759 36159
rect 57701 36119 57759 36125
rect 57793 36159 57851 36165
rect 57793 36125 57805 36159
rect 57839 36156 57851 36159
rect 58084 36156 58112 36196
rect 57839 36128 58112 36156
rect 58529 36159 58587 36165
rect 57839 36125 57851 36128
rect 57793 36119 57851 36125
rect 58529 36125 58541 36159
rect 58575 36156 58587 36159
rect 58575 36128 58940 36156
rect 58575 36125 58587 36128
rect 58529 36119 58587 36125
rect 4614 36088 4620 36100
rect 3804 36060 4620 36088
rect 4614 36048 4620 36060
rect 4672 36048 4678 36100
rect 6454 36088 6460 36100
rect 4908 36060 6460 36088
rect 2222 35980 2228 36032
rect 2280 36020 2286 36032
rect 4908 36020 4936 36060
rect 6454 36048 6460 36060
rect 6512 36048 6518 36100
rect 8297 36091 8355 36097
rect 8297 36057 8309 36091
rect 8343 36088 8355 36091
rect 9324 36088 9352 36119
rect 8343 36060 9352 36088
rect 57517 36091 57575 36097
rect 8343 36057 8355 36060
rect 8297 36051 8355 36057
rect 57517 36057 57529 36091
rect 57563 36088 57575 36091
rect 58434 36088 58440 36100
rect 57563 36060 58440 36088
rect 57563 36057 57575 36060
rect 57517 36051 57575 36057
rect 58434 36048 58440 36060
rect 58492 36048 58498 36100
rect 58912 36032 58940 36128
rect 2280 35992 4936 36020
rect 2280 35980 2286 35992
rect 4982 35980 4988 36032
rect 5040 36020 5046 36032
rect 5169 36023 5227 36029
rect 5169 36020 5181 36023
rect 5040 35992 5181 36020
rect 5040 35980 5046 35992
rect 5169 35989 5181 35992
rect 5215 35989 5227 36023
rect 5169 35983 5227 35989
rect 7837 36023 7895 36029
rect 7837 35989 7849 36023
rect 7883 36020 7895 36023
rect 8478 36020 8484 36032
rect 7883 35992 8484 36020
rect 7883 35989 7895 35992
rect 7837 35983 7895 35989
rect 8478 35980 8484 35992
rect 8536 35980 8542 36032
rect 58342 35980 58348 36032
rect 58400 35980 58406 36032
rect 58894 35980 58900 36032
rect 58952 35980 58958 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 3418 35776 3424 35828
rect 3476 35816 3482 35828
rect 3513 35819 3571 35825
rect 3513 35816 3525 35819
rect 3476 35788 3525 35816
rect 3476 35776 3482 35788
rect 3513 35785 3525 35788
rect 3559 35785 3571 35819
rect 3513 35779 3571 35785
rect 4341 35819 4399 35825
rect 4341 35785 4353 35819
rect 4387 35816 4399 35819
rect 4522 35816 4528 35828
rect 4387 35788 4528 35816
rect 4387 35785 4399 35788
rect 4341 35779 4399 35785
rect 4522 35776 4528 35788
rect 4580 35776 4586 35828
rect 6178 35816 6184 35828
rect 4632 35788 6184 35816
rect 4632 35748 4660 35788
rect 6178 35776 6184 35788
rect 6236 35776 6242 35828
rect 6454 35776 6460 35828
rect 6512 35776 6518 35828
rect 2792 35720 4660 35748
rect 4709 35751 4767 35757
rect 934 35640 940 35692
rect 992 35680 998 35692
rect 2792 35689 2820 35720
rect 4709 35717 4721 35751
rect 4755 35748 4767 35751
rect 4982 35748 4988 35760
rect 4755 35720 4988 35748
rect 4755 35717 4767 35720
rect 4709 35711 4767 35717
rect 4982 35708 4988 35720
rect 5040 35708 5046 35760
rect 6086 35748 6092 35760
rect 5934 35720 6092 35748
rect 6086 35708 6092 35720
rect 6144 35748 6150 35760
rect 7929 35751 7987 35757
rect 6144 35720 6762 35748
rect 6144 35708 6150 35720
rect 7929 35717 7941 35751
rect 7975 35748 7987 35751
rect 8297 35751 8355 35757
rect 8297 35748 8309 35751
rect 7975 35720 8309 35748
rect 7975 35717 7987 35720
rect 7929 35711 7987 35717
rect 8297 35717 8309 35720
rect 8343 35717 8355 35751
rect 8297 35711 8355 35717
rect 58253 35751 58311 35757
rect 58253 35717 58265 35751
rect 58299 35748 58311 35751
rect 58342 35748 58348 35760
rect 58299 35720 58348 35748
rect 58299 35717 58311 35720
rect 58253 35711 58311 35717
rect 58342 35708 58348 35720
rect 58400 35708 58406 35760
rect 1581 35683 1639 35689
rect 1581 35680 1593 35683
rect 992 35652 1593 35680
rect 992 35640 998 35652
rect 1581 35649 1593 35652
rect 1627 35649 1639 35683
rect 1581 35643 1639 35649
rect 2777 35683 2835 35689
rect 2777 35649 2789 35683
rect 2823 35649 2835 35683
rect 2777 35643 2835 35649
rect 2866 35640 2872 35692
rect 2924 35640 2930 35692
rect 4062 35640 4068 35692
rect 4120 35640 4126 35692
rect 4433 35683 4491 35689
rect 4433 35680 4445 35683
rect 4264 35652 4445 35680
rect 3142 35572 3148 35624
rect 3200 35612 3206 35624
rect 4264 35612 4292 35652
rect 4433 35649 4445 35652
rect 4479 35649 4491 35683
rect 9217 35683 9275 35689
rect 9217 35680 9229 35683
rect 4433 35643 4491 35649
rect 8220 35652 9229 35680
rect 3200 35584 4292 35612
rect 4341 35615 4399 35621
rect 3200 35572 3206 35584
rect 4341 35581 4353 35615
rect 4387 35581 4399 35615
rect 4448 35612 4476 35643
rect 8220 35624 8248 35652
rect 9217 35649 9229 35652
rect 9263 35680 9275 35683
rect 10502 35680 10508 35692
rect 9263 35652 10508 35680
rect 9263 35649 9275 35652
rect 9217 35643 9275 35649
rect 10502 35640 10508 35652
rect 10560 35680 10566 35692
rect 17126 35680 17132 35692
rect 10560 35652 17132 35680
rect 10560 35640 10566 35652
rect 17126 35640 17132 35652
rect 17184 35640 17190 35692
rect 58066 35640 58072 35692
rect 58124 35640 58130 35692
rect 58161 35683 58219 35689
rect 58161 35649 58173 35683
rect 58207 35649 58219 35683
rect 58161 35643 58219 35649
rect 5718 35612 5724 35624
rect 4448 35584 5724 35612
rect 4341 35575 4399 35581
rect 2682 35436 2688 35488
rect 2740 35476 2746 35488
rect 3418 35476 3424 35488
rect 2740 35448 3424 35476
rect 2740 35436 2746 35448
rect 3418 35436 3424 35448
rect 3476 35476 3482 35488
rect 3970 35476 3976 35488
rect 3476 35448 3976 35476
rect 3476 35436 3482 35448
rect 3970 35436 3976 35448
rect 4028 35476 4034 35488
rect 4157 35479 4215 35485
rect 4157 35476 4169 35479
rect 4028 35448 4169 35476
rect 4028 35436 4034 35448
rect 4157 35445 4169 35448
rect 4203 35445 4215 35479
rect 4356 35476 4384 35575
rect 5718 35572 5724 35584
rect 5776 35572 5782 35624
rect 8202 35572 8208 35624
rect 8260 35572 8266 35624
rect 8846 35572 8852 35624
rect 8904 35572 8910 35624
rect 58176 35612 58204 35643
rect 58434 35640 58440 35692
rect 58492 35640 58498 35692
rect 57624 35584 58204 35612
rect 4706 35476 4712 35488
rect 4356 35448 4712 35476
rect 4157 35439 4215 35445
rect 4706 35436 4712 35448
rect 4764 35436 4770 35488
rect 56410 35436 56416 35488
rect 56468 35476 56474 35488
rect 57624 35485 57652 35584
rect 57609 35479 57667 35485
rect 57609 35476 57621 35479
rect 56468 35448 57621 35476
rect 56468 35436 56474 35448
rect 57609 35445 57621 35448
rect 57655 35476 57667 35479
rect 57698 35476 57704 35488
rect 57655 35448 57704 35476
rect 57655 35445 57667 35448
rect 57609 35439 57667 35445
rect 57698 35436 57704 35448
rect 57756 35436 57762 35488
rect 57882 35436 57888 35488
rect 57940 35436 57946 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 3326 35232 3332 35284
rect 3384 35272 3390 35284
rect 3421 35275 3479 35281
rect 3421 35272 3433 35275
rect 3384 35244 3433 35272
rect 3384 35232 3390 35244
rect 3421 35241 3433 35244
rect 3467 35241 3479 35275
rect 3421 35235 3479 35241
rect 3878 35232 3884 35284
rect 3936 35232 3942 35284
rect 4706 35232 4712 35284
rect 4764 35232 4770 35284
rect 6178 35232 6184 35284
rect 6236 35232 6242 35284
rect 7377 35275 7435 35281
rect 7377 35241 7389 35275
rect 7423 35272 7435 35275
rect 8846 35272 8852 35284
rect 7423 35244 8852 35272
rect 7423 35241 7435 35244
rect 7377 35235 7435 35241
rect 8846 35232 8852 35244
rect 8904 35232 8910 35284
rect 57425 35275 57483 35281
rect 57425 35272 57437 35275
rect 56060 35244 57437 35272
rect 3528 35176 6132 35204
rect 2501 35071 2559 35077
rect 2501 35037 2513 35071
rect 2547 35068 2559 35071
rect 2590 35068 2596 35080
rect 2547 35040 2596 35068
rect 2547 35037 2559 35040
rect 2501 35031 2559 35037
rect 2590 35028 2596 35040
rect 2648 35028 2654 35080
rect 3528 35077 3556 35176
rect 5353 35139 5411 35145
rect 5353 35105 5365 35139
rect 5399 35136 5411 35139
rect 5537 35139 5595 35145
rect 5537 35136 5549 35139
rect 5399 35108 5549 35136
rect 5399 35105 5411 35108
rect 5353 35099 5411 35105
rect 5537 35105 5549 35108
rect 5583 35105 5595 35139
rect 5537 35099 5595 35105
rect 3329 35071 3387 35077
rect 3329 35037 3341 35071
rect 3375 35037 3387 35071
rect 3329 35031 3387 35037
rect 3513 35071 3571 35077
rect 3513 35037 3525 35071
rect 3559 35037 3571 35071
rect 3789 35071 3847 35077
rect 3789 35068 3801 35071
rect 3513 35031 3571 35037
rect 3712 35040 3801 35068
rect 3344 35000 3372 35031
rect 3712 35012 3740 35040
rect 3789 35037 3801 35040
rect 3835 35037 3847 35071
rect 3789 35031 3847 35037
rect 3973 35071 4031 35077
rect 3973 35037 3985 35071
rect 4019 35068 4031 35071
rect 4982 35068 4988 35080
rect 4019 35040 4988 35068
rect 4019 35037 4031 35040
rect 3973 35031 4031 35037
rect 4982 35028 4988 35040
rect 5040 35028 5046 35080
rect 5445 35071 5503 35077
rect 5445 35037 5457 35071
rect 5491 35037 5503 35071
rect 5445 35031 5503 35037
rect 5629 35071 5687 35077
rect 5629 35037 5641 35071
rect 5675 35068 5687 35071
rect 5721 35071 5779 35077
rect 5721 35068 5733 35071
rect 5675 35040 5733 35068
rect 5675 35037 5687 35040
rect 5629 35031 5687 35037
rect 5721 35037 5733 35040
rect 5767 35037 5779 35071
rect 6104 35068 6132 35176
rect 6196 35136 6224 35232
rect 56060 35216 56088 35244
rect 7282 35164 7288 35216
rect 7340 35164 7346 35216
rect 56042 35164 56048 35216
rect 56100 35164 56106 35216
rect 6273 35139 6331 35145
rect 6273 35136 6285 35139
rect 6196 35108 6285 35136
rect 6273 35105 6285 35108
rect 6319 35105 6331 35139
rect 6273 35099 6331 35105
rect 7469 35139 7527 35145
rect 7469 35105 7481 35139
rect 7515 35136 7527 35139
rect 7745 35139 7803 35145
rect 7745 35136 7757 35139
rect 7515 35108 7757 35136
rect 7515 35105 7527 35108
rect 7469 35099 7527 35105
rect 7745 35105 7757 35108
rect 7791 35105 7803 35139
rect 7745 35099 7803 35105
rect 8389 35139 8447 35145
rect 8389 35105 8401 35139
rect 8435 35136 8447 35139
rect 8573 35139 8631 35145
rect 8573 35136 8585 35139
rect 8435 35108 8585 35136
rect 8435 35105 8447 35108
rect 8389 35099 8447 35105
rect 8573 35105 8585 35108
rect 8619 35105 8631 35139
rect 56229 35139 56287 35145
rect 56229 35136 56241 35139
rect 8573 35099 8631 35105
rect 55968 35108 56241 35136
rect 6638 35068 6644 35080
rect 6104 35040 6644 35068
rect 5721 35031 5779 35037
rect 3694 35000 3700 35012
rect 3344 34972 3700 35000
rect 3694 34960 3700 34972
rect 3752 34960 3758 35012
rect 3050 34892 3056 34944
rect 3108 34892 3114 34944
rect 5166 34892 5172 34944
rect 5224 34932 5230 34944
rect 5460 34932 5488 35031
rect 6638 35028 6644 35040
rect 6696 35028 6702 35080
rect 7193 35071 7251 35077
rect 7193 35037 7205 35071
rect 7239 35037 7251 35071
rect 7193 35031 7251 35037
rect 7208 35000 7236 35031
rect 8478 35028 8484 35080
rect 8536 35028 8542 35080
rect 8665 35071 8723 35077
rect 8665 35037 8677 35071
rect 8711 35068 8723 35071
rect 8754 35068 8760 35080
rect 8711 35040 8760 35068
rect 8711 35037 8723 35040
rect 8665 35031 8723 35037
rect 8294 35000 8300 35012
rect 7208 34972 8300 35000
rect 8294 34960 8300 34972
rect 8352 34960 8358 35012
rect 8680 34932 8708 35031
rect 8754 35028 8760 35040
rect 8812 35068 8818 35080
rect 55585 35071 55643 35077
rect 8812 35040 9168 35068
rect 8812 35028 8818 35040
rect 9140 35012 9168 35040
rect 55585 35037 55597 35071
rect 55631 35068 55643 35071
rect 55769 35071 55827 35077
rect 55631 35040 55720 35068
rect 55631 35037 55643 35040
rect 55585 35031 55643 35037
rect 9122 34960 9128 35012
rect 9180 34960 9186 35012
rect 5224 34904 8708 34932
rect 5224 34892 5230 34904
rect 55306 34892 55312 34944
rect 55364 34932 55370 34944
rect 55585 34935 55643 34941
rect 55585 34932 55597 34935
rect 55364 34904 55597 34932
rect 55364 34892 55370 34904
rect 55585 34901 55597 34904
rect 55631 34901 55643 34935
rect 55692 34932 55720 35040
rect 55769 35037 55781 35071
rect 55815 35037 55827 35071
rect 55769 35031 55827 35037
rect 55784 35000 55812 35031
rect 55858 35028 55864 35080
rect 55916 35028 55922 35080
rect 55968 35000 55996 35108
rect 56229 35105 56241 35108
rect 56275 35105 56287 35139
rect 56229 35099 56287 35105
rect 57072 35080 57100 35244
rect 57425 35241 57437 35244
rect 57471 35241 57483 35275
rect 58345 35275 58403 35281
rect 58345 35272 58357 35275
rect 57425 35235 57483 35241
rect 57532 35244 58357 35272
rect 56045 35071 56103 35077
rect 56045 35037 56057 35071
rect 56091 35037 56103 35071
rect 56045 35031 56103 35037
rect 55784 34972 55996 35000
rect 55953 34935 56011 34941
rect 55953 34932 55965 34935
rect 55692 34904 55965 34932
rect 55585 34895 55643 34901
rect 55953 34901 55965 34904
rect 55999 34901 56011 34935
rect 56060 34932 56088 35031
rect 56134 35028 56140 35080
rect 56192 35028 56198 35080
rect 56329 35071 56387 35077
rect 56329 35037 56341 35071
rect 56375 35068 56387 35071
rect 56962 35068 56968 35080
rect 56375 35040 56968 35068
rect 56375 35037 56387 35040
rect 56329 35031 56387 35037
rect 56962 35028 56968 35040
rect 57020 35028 57026 35080
rect 57054 35028 57060 35080
rect 57112 35028 57118 35080
rect 57238 35028 57244 35080
rect 57296 35028 57302 35080
rect 57333 35071 57391 35077
rect 57333 35037 57345 35071
rect 57379 35068 57391 35071
rect 57532 35068 57560 35244
rect 58345 35241 58357 35244
rect 58391 35241 58403 35275
rect 58345 35235 58403 35241
rect 57885 35207 57943 35213
rect 57885 35173 57897 35207
rect 57931 35173 57943 35207
rect 57885 35167 57943 35173
rect 57609 35139 57667 35145
rect 57609 35105 57621 35139
rect 57655 35136 57667 35139
rect 57698 35136 57704 35148
rect 57655 35108 57704 35136
rect 57655 35105 57667 35108
rect 57609 35099 57667 35105
rect 57698 35096 57704 35108
rect 57756 35096 57762 35148
rect 57900 35136 57928 35167
rect 57900 35108 58204 35136
rect 58176 35077 58204 35108
rect 57379 35040 57560 35068
rect 57977 35071 58035 35077
rect 57379 35037 57391 35040
rect 57333 35031 57391 35037
rect 57977 35037 57989 35071
rect 58023 35037 58035 35071
rect 57977 35031 58035 35037
rect 58161 35071 58219 35077
rect 58161 35037 58173 35071
rect 58207 35037 58219 35071
rect 58161 35031 58219 35037
rect 58529 35071 58587 35077
rect 58529 35037 58541 35071
rect 58575 35037 58587 35071
rect 58529 35031 58587 35037
rect 57149 35003 57207 35009
rect 56336 34972 57008 35000
rect 56336 34932 56364 34972
rect 56060 34904 56364 34932
rect 55953 34895 56011 34901
rect 56410 34892 56416 34944
rect 56468 34932 56474 34944
rect 56873 34935 56931 34941
rect 56873 34932 56885 34935
rect 56468 34904 56885 34932
rect 56468 34892 56474 34904
rect 56873 34901 56885 34904
rect 56919 34901 56931 34935
rect 56980 34932 57008 34972
rect 57149 34969 57161 35003
rect 57195 35000 57207 35003
rect 57992 35000 58020 35031
rect 57195 34972 58020 35000
rect 58544 35000 58572 35031
rect 58894 35000 58900 35012
rect 58544 34972 58900 35000
rect 57195 34969 57207 34972
rect 57149 34963 57207 34969
rect 58894 34960 58900 34972
rect 58952 34960 58958 35012
rect 57977 34935 58035 34941
rect 57977 34932 57989 34935
rect 56980 34904 57989 34932
rect 56873 34895 56931 34901
rect 57977 34901 57989 34904
rect 58023 34901 58035 34935
rect 57977 34895 58035 34901
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 1397 34731 1455 34737
rect 1397 34697 1409 34731
rect 1443 34728 1455 34731
rect 1443 34700 2636 34728
rect 1443 34697 1455 34700
rect 1397 34691 1455 34697
rect 2608 34672 2636 34700
rect 4062 34688 4068 34740
rect 4120 34728 4126 34740
rect 4525 34731 4583 34737
rect 4525 34728 4537 34731
rect 4120 34700 4537 34728
rect 4120 34688 4126 34700
rect 4525 34697 4537 34700
rect 4571 34697 4583 34731
rect 4525 34691 4583 34697
rect 49329 34731 49387 34737
rect 49329 34697 49341 34731
rect 49375 34728 49387 34731
rect 55769 34731 55827 34737
rect 49375 34700 51074 34728
rect 49375 34697 49387 34700
rect 49329 34691 49387 34697
rect 2406 34620 2412 34672
rect 2464 34620 2470 34672
rect 2590 34620 2596 34672
rect 2648 34620 2654 34672
rect 2869 34663 2927 34669
rect 2869 34629 2881 34663
rect 2915 34660 2927 34663
rect 3237 34663 3295 34669
rect 3237 34660 3249 34663
rect 2915 34632 3249 34660
rect 2915 34629 2927 34632
rect 2869 34623 2927 34629
rect 3237 34629 3249 34632
rect 3283 34629 3295 34663
rect 51046 34660 51074 34700
rect 55769 34697 55781 34731
rect 55815 34728 55827 34731
rect 56134 34728 56140 34740
rect 55815 34700 56140 34728
rect 55815 34697 55827 34700
rect 55769 34691 55827 34697
rect 56134 34688 56140 34700
rect 56192 34728 56198 34740
rect 56505 34731 56563 34737
rect 56505 34728 56517 34731
rect 56192 34700 56517 34728
rect 56192 34688 56198 34700
rect 56505 34697 56517 34700
rect 56551 34728 56563 34731
rect 56686 34728 56692 34740
rect 56551 34700 56692 34728
rect 56551 34697 56563 34700
rect 56505 34691 56563 34697
rect 56686 34688 56692 34700
rect 56744 34688 56750 34740
rect 56042 34660 56048 34672
rect 3237 34623 3295 34629
rect 4080 34632 4568 34660
rect 51046 34632 56048 34660
rect 3878 34552 3884 34604
rect 3936 34592 3942 34604
rect 4080 34601 4108 34632
rect 4540 34601 4568 34632
rect 4065 34595 4123 34601
rect 4065 34592 4077 34595
rect 3936 34564 4077 34592
rect 3936 34552 3942 34564
rect 4065 34561 4077 34564
rect 4111 34561 4123 34595
rect 4065 34555 4123 34561
rect 4249 34595 4307 34601
rect 4249 34561 4261 34595
rect 4295 34561 4307 34595
rect 4249 34555 4307 34561
rect 4525 34595 4583 34601
rect 4525 34561 4537 34595
rect 4571 34561 4583 34595
rect 4525 34555 4583 34561
rect 4709 34595 4767 34601
rect 4709 34561 4721 34595
rect 4755 34592 4767 34595
rect 5994 34592 6000 34604
rect 4755 34564 6000 34592
rect 4755 34561 4767 34564
rect 4709 34555 4767 34561
rect 3142 34484 3148 34536
rect 3200 34484 3206 34536
rect 3418 34484 3424 34536
rect 3476 34524 3482 34536
rect 3789 34527 3847 34533
rect 3789 34524 3801 34527
rect 3476 34496 3801 34524
rect 3476 34484 3482 34496
rect 3789 34493 3801 34496
rect 3835 34493 3847 34527
rect 4264 34524 4292 34555
rect 5994 34552 6000 34564
rect 6052 34552 6058 34604
rect 49694 34552 49700 34604
rect 49752 34552 49758 34604
rect 51184 34601 51212 34632
rect 51169 34595 51227 34601
rect 51169 34561 51181 34595
rect 51215 34561 51227 34595
rect 51169 34555 51227 34561
rect 51905 34595 51963 34601
rect 51905 34561 51917 34595
rect 51951 34561 51963 34595
rect 51905 34555 51963 34561
rect 9858 34524 9864 34536
rect 4264 34496 9864 34524
rect 3789 34487 3847 34493
rect 9858 34484 9864 34496
rect 9916 34484 9922 34536
rect 50798 34484 50804 34536
rect 50856 34484 50862 34536
rect 51077 34527 51135 34533
rect 51077 34493 51089 34527
rect 51123 34524 51135 34527
rect 51442 34524 51448 34536
rect 51123 34496 51448 34524
rect 51123 34493 51135 34496
rect 51077 34487 51135 34493
rect 51442 34484 51448 34496
rect 51500 34484 51506 34536
rect 4157 34459 4215 34465
rect 4157 34425 4169 34459
rect 4203 34456 4215 34459
rect 4614 34456 4620 34468
rect 4203 34428 4620 34456
rect 4203 34425 4215 34428
rect 4157 34419 4215 34425
rect 4614 34416 4620 34428
rect 4672 34416 4678 34468
rect 51920 34456 51948 34555
rect 55490 34552 55496 34604
rect 55548 34552 55554 34604
rect 55692 34601 55720 34632
rect 56042 34620 56048 34632
rect 56100 34620 56106 34672
rect 56226 34620 56232 34672
rect 56284 34660 56290 34672
rect 57241 34663 57299 34669
rect 57241 34660 57253 34663
rect 56284 34632 56456 34660
rect 56284 34620 56290 34632
rect 55677 34595 55735 34601
rect 55677 34561 55689 34595
rect 55723 34561 55735 34595
rect 55677 34555 55735 34561
rect 55858 34552 55864 34604
rect 55916 34552 55922 34604
rect 56321 34595 56379 34601
rect 56321 34561 56333 34595
rect 56367 34561 56379 34595
rect 56428 34592 56456 34632
rect 56796 34632 57253 34660
rect 56597 34595 56655 34601
rect 56597 34592 56609 34595
rect 56428 34564 56609 34592
rect 56321 34555 56379 34561
rect 56597 34561 56609 34564
rect 56643 34561 56655 34595
rect 56597 34555 56655 34561
rect 55508 34524 55536 34552
rect 55876 34524 55904 34552
rect 55508 34496 55904 34524
rect 56336 34524 56364 34555
rect 56686 34552 56692 34604
rect 56744 34552 56750 34604
rect 56796 34524 56824 34632
rect 57241 34629 57253 34632
rect 57287 34629 57299 34663
rect 57241 34623 57299 34629
rect 56870 34552 56876 34604
rect 56928 34552 56934 34604
rect 57425 34595 57483 34601
rect 57425 34561 57437 34595
rect 57471 34561 57483 34595
rect 57425 34555 57483 34561
rect 57440 34524 57468 34555
rect 57514 34552 57520 34604
rect 57572 34592 57578 34604
rect 57609 34595 57667 34601
rect 57609 34592 57621 34595
rect 57572 34564 57621 34592
rect 57572 34552 57578 34564
rect 57609 34561 57621 34564
rect 57655 34561 57667 34595
rect 57609 34555 57667 34561
rect 58529 34595 58587 34601
rect 58529 34561 58541 34595
rect 58575 34561 58587 34595
rect 58529 34555 58587 34561
rect 56336 34496 56824 34524
rect 56888 34496 57468 34524
rect 57701 34527 57759 34533
rect 51368 34428 51948 34456
rect 55876 34456 55904 34496
rect 55876 34428 56456 34456
rect 51166 34348 51172 34400
rect 51224 34388 51230 34400
rect 51368 34397 51396 34428
rect 51353 34391 51411 34397
rect 51353 34388 51365 34391
rect 51224 34360 51365 34388
rect 51224 34348 51230 34360
rect 51353 34357 51365 34360
rect 51399 34357 51411 34391
rect 51353 34351 51411 34357
rect 51997 34391 52055 34397
rect 51997 34357 52009 34391
rect 52043 34388 52055 34391
rect 52178 34388 52184 34400
rect 52043 34360 52184 34388
rect 52043 34357 52055 34360
rect 51997 34351 52055 34357
rect 52178 34348 52184 34360
rect 52236 34348 52242 34400
rect 56318 34348 56324 34400
rect 56376 34348 56382 34400
rect 56428 34388 56456 34428
rect 56502 34416 56508 34468
rect 56560 34456 56566 34468
rect 56781 34459 56839 34465
rect 56781 34456 56793 34459
rect 56560 34428 56793 34456
rect 56560 34416 56566 34428
rect 56781 34425 56793 34428
rect 56827 34425 56839 34459
rect 56781 34419 56839 34425
rect 56888 34388 56916 34496
rect 57701 34493 57713 34527
rect 57747 34524 57759 34527
rect 57974 34524 57980 34536
rect 57747 34496 57980 34524
rect 57747 34493 57759 34496
rect 57701 34487 57759 34493
rect 57974 34484 57980 34496
rect 58032 34484 58038 34536
rect 58544 34524 58572 34555
rect 58894 34524 58900 34536
rect 58544 34496 58900 34524
rect 58894 34484 58900 34496
rect 58952 34484 58958 34536
rect 56428 34360 56916 34388
rect 58342 34348 58348 34400
rect 58400 34348 58406 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 3053 34187 3111 34193
rect 3053 34153 3065 34187
rect 3099 34184 3111 34187
rect 3418 34184 3424 34196
rect 3099 34156 3424 34184
rect 3099 34153 3111 34156
rect 3053 34147 3111 34153
rect 3418 34144 3424 34156
rect 3476 34144 3482 34196
rect 5994 34144 6000 34196
rect 6052 34184 6058 34196
rect 6546 34184 6552 34196
rect 6052 34156 6552 34184
rect 6052 34144 6058 34156
rect 6546 34144 6552 34156
rect 6604 34184 6610 34196
rect 7009 34187 7067 34193
rect 7009 34184 7021 34187
rect 6604 34156 7021 34184
rect 6604 34144 6610 34156
rect 7009 34153 7021 34156
rect 7055 34153 7067 34187
rect 7009 34147 7067 34153
rect 50798 34144 50804 34196
rect 50856 34144 50862 34196
rect 52638 34144 52644 34196
rect 52696 34184 52702 34196
rect 56410 34184 56416 34196
rect 52696 34156 56416 34184
rect 52696 34144 52702 34156
rect 56410 34144 56416 34156
rect 56468 34144 56474 34196
rect 57974 34144 57980 34196
rect 58032 34144 58038 34196
rect 58161 34187 58219 34193
rect 58161 34153 58173 34187
rect 58207 34184 58219 34187
rect 58342 34184 58348 34196
rect 58207 34156 58348 34184
rect 58207 34153 58219 34156
rect 58161 34147 58219 34153
rect 58342 34144 58348 34156
rect 58400 34144 58406 34196
rect 3789 34119 3847 34125
rect 3789 34116 3801 34119
rect 3160 34088 3801 34116
rect 934 34008 940 34060
rect 992 34048 998 34060
rect 3160 34057 3188 34088
rect 3789 34085 3801 34088
rect 3835 34085 3847 34119
rect 3789 34079 3847 34085
rect 1581 34051 1639 34057
rect 1581 34048 1593 34051
rect 992 34020 1593 34048
rect 992 34008 998 34020
rect 1581 34017 1593 34020
rect 1627 34017 1639 34051
rect 1581 34011 1639 34017
rect 3145 34051 3203 34057
rect 3145 34017 3157 34051
rect 3191 34017 3203 34051
rect 3145 34011 3203 34017
rect 3329 34051 3387 34057
rect 3329 34017 3341 34051
rect 3375 34048 3387 34051
rect 4341 34051 4399 34057
rect 4341 34048 4353 34051
rect 3375 34020 4353 34048
rect 3375 34017 3387 34020
rect 3329 34011 3387 34017
rect 4341 34017 4353 34020
rect 4387 34017 4399 34051
rect 4341 34011 4399 34017
rect 57333 34051 57391 34057
rect 57333 34017 57345 34051
rect 57379 34048 57391 34051
rect 57790 34048 57796 34060
rect 57379 34020 57796 34048
rect 57379 34017 57391 34020
rect 57333 34011 57391 34017
rect 57790 34008 57796 34020
rect 57848 34008 57854 34060
rect 2590 33940 2596 33992
rect 2648 33940 2654 33992
rect 2866 33940 2872 33992
rect 2924 33940 2930 33992
rect 2961 33983 3019 33989
rect 2961 33949 2973 33983
rect 3007 33949 3019 33983
rect 2961 33943 3019 33949
rect 2976 33912 3004 33943
rect 3050 33940 3056 33992
rect 3108 33980 3114 33992
rect 3237 33983 3295 33989
rect 3237 33980 3249 33983
rect 3108 33952 3249 33980
rect 3108 33940 3114 33952
rect 3237 33949 3249 33952
rect 3283 33949 3295 33983
rect 3237 33943 3295 33949
rect 3421 33983 3479 33989
rect 3421 33949 3433 33983
rect 3467 33980 3479 33983
rect 5166 33980 5172 33992
rect 3467 33952 5172 33980
rect 3467 33949 3479 33952
rect 3421 33943 3479 33949
rect 5166 33940 5172 33952
rect 5224 33940 5230 33992
rect 5353 33983 5411 33989
rect 5353 33949 5365 33983
rect 5399 33949 5411 33983
rect 5353 33943 5411 33949
rect 5445 33983 5503 33989
rect 5445 33949 5457 33983
rect 5491 33980 5503 33983
rect 5629 33983 5687 33989
rect 5629 33980 5641 33983
rect 5491 33952 5641 33980
rect 5491 33949 5503 33952
rect 5445 33943 5503 33949
rect 5629 33949 5641 33952
rect 5675 33949 5687 33983
rect 5629 33943 5687 33949
rect 3326 33912 3332 33924
rect 2976 33884 3332 33912
rect 3326 33872 3332 33884
rect 3384 33872 3390 33924
rect 4798 33804 4804 33856
rect 4856 33844 4862 33856
rect 5261 33847 5319 33853
rect 5261 33844 5273 33847
rect 4856 33816 5273 33844
rect 4856 33804 4862 33816
rect 5261 33813 5273 33816
rect 5307 33844 5319 33847
rect 5368 33844 5396 33943
rect 9306 33940 9312 33992
rect 9364 33940 9370 33992
rect 41598 33940 41604 33992
rect 41656 33940 41662 33992
rect 43010 33966 44220 33980
rect 42996 33952 44220 33966
rect 5902 33921 5908 33924
rect 5896 33875 5908 33921
rect 5902 33872 5908 33875
rect 5960 33872 5966 33924
rect 9398 33872 9404 33924
rect 9456 33912 9462 33924
rect 9554 33915 9612 33921
rect 9554 33912 9566 33915
rect 9456 33884 9566 33912
rect 9456 33872 9462 33884
rect 9554 33881 9566 33884
rect 9600 33881 9612 33915
rect 9554 33875 9612 33881
rect 41874 33872 41880 33924
rect 41932 33872 41938 33924
rect 6730 33844 6736 33856
rect 5307 33816 6736 33844
rect 5307 33813 5319 33816
rect 5261 33807 5319 33813
rect 6730 33804 6736 33816
rect 6788 33844 6794 33856
rect 7377 33847 7435 33853
rect 7377 33844 7389 33847
rect 6788 33816 7389 33844
rect 6788 33804 6794 33816
rect 7377 33813 7389 33816
rect 7423 33844 7435 33847
rect 9766 33844 9772 33856
rect 7423 33816 9772 33844
rect 7423 33813 7435 33816
rect 7377 33807 7435 33813
rect 9766 33804 9772 33816
rect 9824 33804 9830 33856
rect 9858 33804 9864 33856
rect 9916 33844 9922 33856
rect 10689 33847 10747 33853
rect 10689 33844 10701 33847
rect 9916 33816 10701 33844
rect 9916 33804 9922 33816
rect 10689 33813 10701 33816
rect 10735 33813 10747 33847
rect 10689 33807 10747 33813
rect 42610 33804 42616 33856
rect 42668 33844 42674 33856
rect 42996 33844 43024 33952
rect 44192 33924 44220 33952
rect 45646 33940 45652 33992
rect 45704 33940 45710 33992
rect 50154 33940 50160 33992
rect 50212 33940 50218 33992
rect 57054 33940 57060 33992
rect 57112 33980 57118 33992
rect 57241 33983 57299 33989
rect 57241 33980 57253 33983
rect 57112 33952 57253 33980
rect 57112 33940 57118 33952
rect 57241 33949 57253 33952
rect 57287 33949 57299 33983
rect 57241 33943 57299 33949
rect 57425 33983 57483 33989
rect 57425 33949 57437 33983
rect 57471 33980 57483 33983
rect 57606 33980 57612 33992
rect 57471 33952 57612 33980
rect 57471 33949 57483 33952
rect 57425 33943 57483 33949
rect 57606 33940 57612 33952
rect 57664 33940 57670 33992
rect 57882 33940 57888 33992
rect 57940 33940 57946 33992
rect 43441 33915 43499 33921
rect 43441 33881 43453 33915
rect 43487 33881 43499 33915
rect 43441 33875 43499 33881
rect 42668 33816 43024 33844
rect 42668 33804 42674 33816
rect 43254 33804 43260 33856
rect 43312 33844 43318 33856
rect 43349 33847 43407 33853
rect 43349 33844 43361 33847
rect 43312 33816 43361 33844
rect 43312 33804 43318 33816
rect 43349 33813 43361 33816
rect 43395 33813 43407 33847
rect 43456 33844 43484 33875
rect 44174 33872 44180 33924
rect 44232 33872 44238 33924
rect 44729 33915 44787 33921
rect 44729 33881 44741 33915
rect 44775 33912 44787 33915
rect 44775 33884 46428 33912
rect 44775 33881 44787 33884
rect 44729 33875 44787 33881
rect 44744 33844 44772 33875
rect 46400 33856 46428 33884
rect 51258 33872 51264 33924
rect 51316 33912 51322 33924
rect 57900 33912 57928 33940
rect 51316 33884 57928 33912
rect 51316 33872 51322 33884
rect 57974 33872 57980 33924
rect 58032 33912 58038 33924
rect 58345 33915 58403 33921
rect 58345 33912 58357 33915
rect 58032 33884 58357 33912
rect 58032 33872 58038 33884
rect 58345 33881 58357 33884
rect 58391 33912 58403 33915
rect 58434 33912 58440 33924
rect 58391 33884 58440 33912
rect 58391 33881 58403 33884
rect 58345 33875 58403 33881
rect 58434 33872 58440 33884
rect 58492 33872 58498 33924
rect 43456 33816 44772 33844
rect 43349 33807 43407 33813
rect 45462 33804 45468 33856
rect 45520 33804 45526 33856
rect 46382 33804 46388 33856
rect 46440 33804 46446 33856
rect 51534 33804 51540 33856
rect 51592 33844 51598 33856
rect 56594 33844 56600 33856
rect 51592 33816 56600 33844
rect 51592 33804 51598 33816
rect 56594 33804 56600 33816
rect 56652 33804 56658 33856
rect 57514 33804 57520 33856
rect 57572 33844 57578 33856
rect 57793 33847 57851 33853
rect 57793 33844 57805 33847
rect 57572 33816 57805 33844
rect 57572 33804 57578 33816
rect 57793 33813 57805 33816
rect 57839 33844 57851 33847
rect 58135 33847 58193 33853
rect 58135 33844 58147 33847
rect 57839 33816 58147 33844
rect 57839 33813 57851 33816
rect 57793 33807 57851 33813
rect 58135 33813 58147 33816
rect 58181 33813 58193 33847
rect 58135 33807 58193 33813
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 3237 33643 3295 33649
rect 3237 33609 3249 33643
rect 3283 33640 3295 33643
rect 4798 33640 4804 33652
rect 3283 33612 4804 33640
rect 3283 33609 3295 33612
rect 3237 33603 3295 33609
rect 3344 33513 3372 33612
rect 4798 33600 4804 33612
rect 4856 33600 4862 33652
rect 4982 33600 4988 33652
rect 5040 33600 5046 33652
rect 5092 33612 5856 33640
rect 5092 33513 5120 33612
rect 5258 33532 5264 33584
rect 5316 33532 5322 33584
rect 5828 33581 5856 33612
rect 5902 33600 5908 33652
rect 5960 33649 5966 33652
rect 5960 33640 5969 33649
rect 5960 33612 6005 33640
rect 5960 33603 5969 33612
rect 5960 33600 5966 33603
rect 6546 33600 6552 33652
rect 6604 33600 6610 33652
rect 6638 33600 6644 33652
rect 6696 33600 6702 33652
rect 8665 33643 8723 33649
rect 8665 33640 8677 33643
rect 7024 33612 8677 33640
rect 5537 33575 5595 33581
rect 5537 33572 5549 33575
rect 5368 33544 5549 33572
rect 5368 33513 5396 33544
rect 5537 33541 5549 33544
rect 5583 33541 5595 33575
rect 5537 33535 5595 33541
rect 5813 33575 5871 33581
rect 5813 33541 5825 33575
rect 5859 33572 5871 33575
rect 6454 33572 6460 33584
rect 5859 33544 6460 33572
rect 5859 33541 5871 33544
rect 5813 33535 5871 33541
rect 6454 33532 6460 33544
rect 6512 33532 6518 33584
rect 3329 33507 3387 33513
rect 3329 33473 3341 33507
rect 3375 33473 3387 33507
rect 3329 33467 3387 33473
rect 3872 33507 3930 33513
rect 3872 33473 3884 33507
rect 3918 33504 3930 33507
rect 5077 33507 5135 33513
rect 3918 33476 4660 33504
rect 3918 33473 3930 33476
rect 3872 33467 3930 33473
rect 3421 33439 3479 33445
rect 3421 33405 3433 33439
rect 3467 33436 3479 33439
rect 3605 33439 3663 33445
rect 3605 33436 3617 33439
rect 3467 33408 3617 33436
rect 3467 33405 3479 33408
rect 3421 33399 3479 33405
rect 3605 33405 3617 33408
rect 3651 33405 3663 33439
rect 3605 33399 3663 33405
rect 4632 33368 4660 33476
rect 5077 33473 5089 33507
rect 5123 33473 5135 33507
rect 5077 33467 5135 33473
rect 5353 33507 5411 33513
rect 5353 33473 5365 33507
rect 5399 33473 5411 33507
rect 5353 33467 5411 33473
rect 5445 33507 5503 33513
rect 5445 33473 5457 33507
rect 5491 33473 5503 33507
rect 5445 33467 5503 33473
rect 5629 33507 5687 33513
rect 5629 33473 5641 33507
rect 5675 33473 5687 33507
rect 5629 33467 5687 33473
rect 4982 33396 4988 33448
rect 5040 33436 5046 33448
rect 5460 33436 5488 33467
rect 5040 33408 5488 33436
rect 5040 33396 5046 33408
rect 5077 33371 5135 33377
rect 5077 33368 5089 33371
rect 4632 33340 5089 33368
rect 5077 33337 5089 33340
rect 5123 33337 5135 33371
rect 5644 33368 5672 33467
rect 5994 33464 6000 33516
rect 6052 33464 6058 33516
rect 6089 33507 6147 33513
rect 6089 33473 6101 33507
rect 6135 33473 6147 33507
rect 6089 33467 6147 33473
rect 6104 33436 6132 33467
rect 6362 33464 6368 33516
rect 6420 33464 6426 33516
rect 6564 33513 6592 33600
rect 6656 33572 6684 33600
rect 7024 33572 7052 33612
rect 8665 33609 8677 33612
rect 8711 33609 8723 33643
rect 8665 33603 8723 33609
rect 9306 33600 9312 33652
rect 9364 33600 9370 33652
rect 9769 33643 9827 33649
rect 9769 33640 9781 33643
rect 9600 33612 9781 33640
rect 7466 33572 7472 33584
rect 6656 33544 7052 33572
rect 6549 33507 6607 33513
rect 6549 33473 6561 33507
rect 6595 33473 6607 33507
rect 6549 33467 6607 33473
rect 6730 33464 6736 33516
rect 6788 33464 6794 33516
rect 7024 33513 7052 33544
rect 7208 33544 7472 33572
rect 7208 33513 7236 33544
rect 7466 33532 7472 33544
rect 7524 33532 7530 33584
rect 7742 33532 7748 33584
rect 7800 33572 7806 33584
rect 9030 33572 9036 33584
rect 7800 33544 9036 33572
rect 7800 33532 7806 33544
rect 9030 33532 9036 33544
rect 9088 33532 9094 33584
rect 9324 33572 9352 33600
rect 9232 33544 9352 33572
rect 7558 33513 7564 33516
rect 7009 33507 7067 33513
rect 7009 33473 7021 33507
rect 7055 33473 7067 33507
rect 7009 33467 7067 33473
rect 7193 33507 7251 33513
rect 7193 33473 7205 33507
rect 7239 33473 7251 33507
rect 7552 33504 7564 33513
rect 7519 33476 7564 33504
rect 7193 33467 7251 33473
rect 7552 33467 7564 33476
rect 7558 33464 7564 33467
rect 7616 33464 7622 33516
rect 7834 33464 7840 33516
rect 7892 33504 7898 33516
rect 9125 33507 9183 33513
rect 9125 33504 9137 33507
rect 7892 33476 9137 33504
rect 7892 33464 7898 33476
rect 9125 33473 9137 33476
rect 9171 33473 9183 33507
rect 9125 33467 9183 33473
rect 6457 33439 6515 33445
rect 6457 33436 6469 33439
rect 6104 33408 6469 33436
rect 6457 33405 6469 33408
rect 6503 33405 6515 33439
rect 6457 33399 6515 33405
rect 6825 33439 6883 33445
rect 6825 33405 6837 33439
rect 6871 33436 6883 33439
rect 7285 33439 7343 33445
rect 7285 33436 7297 33439
rect 6871 33408 7297 33436
rect 6871 33405 6883 33408
rect 6825 33399 6883 33405
rect 7285 33405 7297 33408
rect 7331 33405 7343 33439
rect 9232 33436 9260 33544
rect 9306 33464 9312 33516
rect 9364 33464 9370 33516
rect 9401 33507 9459 33513
rect 9401 33473 9413 33507
rect 9447 33504 9459 33507
rect 9600 33504 9628 33612
rect 9769 33609 9781 33612
rect 9815 33609 9827 33643
rect 9769 33603 9827 33609
rect 9858 33600 9864 33652
rect 9916 33600 9922 33652
rect 41874 33600 41880 33652
rect 41932 33640 41938 33652
rect 42429 33643 42487 33649
rect 42429 33640 42441 33643
rect 41932 33612 42441 33640
rect 41932 33600 41938 33612
rect 42429 33609 42441 33612
rect 42475 33609 42487 33643
rect 44269 33643 44327 33649
rect 44269 33640 44281 33643
rect 42429 33603 42487 33609
rect 43180 33612 44281 33640
rect 9876 33572 9904 33600
rect 42153 33575 42211 33581
rect 9876 33544 9996 33572
rect 9968 33513 9996 33544
rect 42153 33541 42165 33575
rect 42199 33572 42211 33575
rect 43180 33572 43208 33612
rect 44269 33609 44281 33612
rect 44315 33609 44327 33643
rect 44269 33603 44327 33609
rect 44545 33643 44603 33649
rect 44545 33609 44557 33643
rect 44591 33640 44603 33643
rect 45646 33640 45652 33652
rect 44591 33612 45652 33640
rect 44591 33609 44603 33612
rect 44545 33603 44603 33609
rect 42199 33544 43208 33572
rect 42199 33541 42211 33544
rect 42153 33535 42211 33541
rect 43254 33532 43260 33584
rect 43312 33572 43318 33584
rect 44284 33572 44312 33603
rect 45646 33600 45652 33612
rect 45704 33600 45710 33652
rect 49510 33640 49516 33652
rect 49160 33612 49516 33640
rect 44634 33572 44640 33584
rect 43312 33544 43484 33572
rect 44284 33544 44640 33572
rect 43312 33532 43318 33544
rect 9447 33476 9628 33504
rect 9677 33507 9735 33513
rect 9447 33473 9459 33476
rect 9401 33467 9459 33473
rect 9677 33473 9689 33507
rect 9723 33473 9735 33507
rect 9677 33467 9735 33473
rect 9769 33507 9827 33513
rect 9769 33473 9781 33507
rect 9815 33473 9827 33507
rect 9769 33467 9827 33473
rect 9953 33507 10011 33513
rect 9953 33473 9965 33507
rect 9999 33473 10011 33507
rect 9953 33467 10011 33473
rect 42245 33507 42303 33513
rect 42245 33473 42257 33507
rect 42291 33504 42303 33507
rect 42886 33504 42892 33516
rect 42291 33476 42892 33504
rect 42291 33473 42303 33476
rect 42245 33467 42303 33473
rect 9585 33439 9643 33445
rect 9585 33436 9597 33439
rect 9232 33408 9597 33436
rect 7285 33399 7343 33405
rect 9585 33405 9597 33408
rect 9631 33405 9643 33439
rect 9585 33399 9643 33405
rect 6362 33368 6368 33380
rect 5644 33340 6368 33368
rect 5077 33331 5135 33337
rect 6362 33328 6368 33340
rect 6420 33328 6426 33380
rect 9398 33328 9404 33380
rect 9456 33328 9462 33380
rect 5534 33260 5540 33312
rect 5592 33300 5598 33312
rect 5994 33300 6000 33312
rect 5592 33272 6000 33300
rect 5592 33260 5598 33272
rect 5994 33260 6000 33272
rect 6052 33260 6058 33312
rect 7098 33260 7104 33312
rect 7156 33260 7162 33312
rect 9125 33303 9183 33309
rect 9125 33269 9137 33303
rect 9171 33300 9183 33303
rect 9416 33300 9444 33328
rect 9171 33272 9444 33300
rect 9692 33300 9720 33467
rect 9784 33436 9812 33467
rect 42886 33464 42892 33476
rect 42944 33464 42950 33516
rect 43456 33513 43484 33544
rect 44634 33532 44640 33544
rect 44692 33532 44698 33584
rect 46845 33575 46903 33581
rect 46845 33572 46857 33575
rect 45586 33544 46857 33572
rect 46400 33516 46428 33544
rect 46845 33541 46857 33544
rect 46891 33541 46903 33575
rect 49160 33572 49188 33612
rect 49510 33600 49516 33612
rect 49568 33600 49574 33652
rect 49605 33643 49663 33649
rect 49605 33609 49617 33643
rect 49651 33609 49663 33643
rect 49605 33603 49663 33609
rect 49082 33544 49188 33572
rect 46845 33535 46903 33541
rect 49234 33532 49240 33584
rect 49292 33572 49298 33584
rect 49620 33572 49648 33603
rect 50154 33600 50160 33652
rect 50212 33600 50218 33652
rect 52638 33640 52644 33652
rect 50264 33612 51764 33640
rect 50264 33572 50292 33612
rect 49292 33544 50292 33572
rect 50663 33575 50721 33581
rect 49292 33532 49298 33544
rect 50663 33541 50675 33575
rect 50709 33572 50721 33575
rect 50890 33572 50896 33584
rect 50709 33544 50896 33572
rect 50709 33541 50721 33544
rect 50663 33535 50721 33541
rect 50890 33532 50896 33544
rect 50948 33532 50954 33584
rect 43165 33507 43223 33513
rect 43165 33473 43177 33507
rect 43211 33504 43223 33507
rect 43349 33507 43407 33513
rect 43211 33476 43300 33504
rect 43211 33473 43223 33476
rect 43165 33467 43223 33473
rect 43272 33448 43300 33476
rect 43349 33473 43361 33507
rect 43395 33473 43407 33507
rect 43349 33467 43407 33473
rect 43441 33507 43499 33513
rect 43441 33473 43453 33507
rect 43487 33473 43499 33507
rect 43441 33467 43499 33473
rect 44177 33507 44235 33513
rect 44177 33473 44189 33507
rect 44223 33473 44235 33507
rect 44177 33467 44235 33473
rect 41785 33439 41843 33445
rect 9784 33408 10364 33436
rect 10336 33380 10364 33408
rect 41785 33405 41797 33439
rect 41831 33405 41843 33439
rect 41785 33399 41843 33405
rect 41969 33439 42027 33445
rect 41969 33405 41981 33439
rect 42015 33436 42027 33439
rect 42981 33439 43039 33445
rect 42981 33436 42993 33439
rect 42015 33408 42993 33436
rect 42015 33405 42027 33408
rect 41969 33399 42027 33405
rect 42981 33405 42993 33408
rect 43027 33405 43039 33439
rect 42981 33399 43039 33405
rect 10318 33328 10324 33380
rect 10376 33328 10382 33380
rect 41800 33368 41828 33399
rect 43254 33396 43260 33448
rect 43312 33396 43318 33448
rect 43364 33436 43392 33467
rect 44085 33439 44143 33445
rect 44085 33436 44097 33439
rect 43364 33408 44097 33436
rect 44085 33405 44097 33408
rect 44131 33436 44143 33439
rect 44192 33436 44220 33467
rect 46382 33464 46388 33516
rect 46440 33464 46446 33516
rect 46474 33464 46480 33516
rect 46532 33464 46538 33516
rect 47394 33504 47400 33516
rect 46952 33476 47400 33504
rect 44131 33408 44220 33436
rect 44131 33405 44143 33408
rect 44085 33399 44143 33405
rect 46014 33396 46020 33448
rect 46072 33396 46078 33448
rect 46293 33439 46351 33445
rect 46293 33405 46305 33439
rect 46339 33436 46351 33439
rect 46952 33436 46980 33476
rect 47394 33464 47400 33476
rect 47452 33504 47458 33516
rect 47581 33507 47639 33513
rect 47581 33504 47593 33507
rect 47452 33476 47593 33504
rect 47452 33464 47458 33476
rect 47581 33473 47593 33476
rect 47627 33473 47639 33507
rect 47581 33467 47639 33473
rect 49421 33507 49479 33513
rect 49421 33473 49433 33507
rect 49467 33473 49479 33507
rect 49421 33467 49479 33473
rect 46339 33408 46980 33436
rect 46339 33405 46351 33408
rect 46293 33399 46351 33405
rect 47854 33396 47860 33448
rect 47912 33396 47918 33448
rect 49329 33439 49387 33445
rect 49329 33405 49341 33439
rect 49375 33436 49387 33439
rect 49436 33436 49464 33467
rect 49786 33464 49792 33516
rect 49844 33504 49850 33516
rect 51092 33513 51120 33612
rect 51166 33532 51172 33584
rect 51224 33572 51230 33584
rect 51224 33544 51672 33572
rect 51224 33532 51230 33544
rect 50341 33507 50399 33513
rect 50341 33504 50353 33507
rect 49844 33476 50353 33504
rect 49844 33464 49850 33476
rect 50341 33473 50353 33476
rect 50387 33473 50399 33507
rect 50341 33467 50399 33473
rect 50433 33507 50491 33513
rect 50433 33473 50445 33507
rect 50479 33473 50491 33507
rect 50433 33467 50491 33473
rect 50525 33507 50583 33513
rect 50525 33473 50537 33507
rect 50571 33504 50583 33507
rect 51077 33507 51135 33513
rect 50571 33476 50936 33504
rect 50571 33473 50583 33476
rect 50525 33467 50583 33473
rect 49375 33408 49464 33436
rect 49375 33405 49387 33408
rect 49329 33399 49387 33405
rect 50448 33380 50476 33467
rect 50798 33396 50804 33448
rect 50856 33396 50862 33448
rect 50908 33436 50936 33476
rect 51077 33473 51089 33507
rect 51123 33473 51135 33507
rect 51077 33467 51135 33473
rect 51258 33464 51264 33516
rect 51316 33464 51322 33516
rect 51353 33507 51411 33513
rect 51353 33473 51365 33507
rect 51399 33473 51411 33507
rect 51353 33467 51411 33473
rect 51445 33507 51503 33513
rect 51445 33473 51457 33507
rect 51491 33504 51503 33507
rect 51534 33504 51540 33516
rect 51491 33476 51540 33504
rect 51491 33473 51503 33476
rect 51445 33467 51503 33473
rect 51368 33436 51396 33467
rect 51534 33464 51540 33476
rect 51592 33464 51598 33516
rect 51644 33513 51672 33544
rect 51736 33513 51764 33612
rect 52012 33612 52644 33640
rect 52012 33513 52040 33612
rect 52638 33600 52644 33612
rect 52696 33600 52702 33652
rect 55674 33600 55680 33652
rect 55732 33600 55738 33652
rect 56594 33600 56600 33652
rect 56652 33640 56658 33652
rect 56781 33643 56839 33649
rect 56781 33640 56793 33643
rect 56652 33612 56793 33640
rect 56652 33600 56658 33612
rect 56781 33609 56793 33612
rect 56827 33640 56839 33643
rect 57330 33640 57336 33652
rect 56827 33612 57336 33640
rect 56827 33609 56839 33612
rect 56781 33603 56839 33609
rect 57330 33600 57336 33612
rect 57388 33600 57394 33652
rect 58158 33600 58164 33652
rect 58216 33600 58222 33652
rect 58176 33572 58204 33600
rect 52196 33544 55812 33572
rect 52196 33516 52224 33544
rect 51629 33507 51687 33513
rect 51629 33473 51641 33507
rect 51675 33473 51687 33507
rect 51629 33467 51687 33473
rect 51721 33507 51779 33513
rect 51721 33473 51733 33507
rect 51767 33473 51779 33507
rect 51721 33467 51779 33473
rect 51997 33507 52055 33513
rect 51997 33473 52009 33507
rect 52043 33473 52055 33507
rect 51997 33467 52055 33473
rect 52178 33464 52184 33516
rect 52236 33464 52242 33516
rect 55490 33464 55496 33516
rect 55548 33464 55554 33516
rect 55784 33513 55812 33544
rect 57440 33544 58204 33572
rect 55769 33507 55827 33513
rect 55769 33473 55781 33507
rect 55815 33504 55827 33507
rect 56594 33504 56600 33516
rect 55815 33476 56600 33504
rect 55815 33473 55827 33476
rect 55769 33467 55827 33473
rect 56594 33464 56600 33476
rect 56652 33464 56658 33516
rect 57333 33507 57391 33513
rect 57333 33473 57345 33507
rect 57379 33473 57391 33507
rect 57333 33467 57391 33473
rect 52089 33439 52147 33445
rect 52089 33436 52101 33439
rect 50908 33408 52101 33436
rect 52089 33405 52101 33408
rect 52135 33405 52147 33439
rect 52089 33399 52147 33405
rect 43806 33368 43812 33380
rect 41800 33340 43812 33368
rect 43806 33328 43812 33340
rect 43864 33328 43870 33380
rect 50430 33328 50436 33380
rect 50488 33368 50494 33380
rect 51537 33371 51595 33377
rect 51537 33368 51549 33371
rect 50488 33340 51549 33368
rect 50488 33328 50494 33340
rect 51537 33337 51549 33340
rect 51583 33337 51595 33371
rect 55508 33368 55536 33464
rect 51537 33331 51595 33337
rect 51828 33340 55536 33368
rect 57348 33368 57376 33467
rect 57440 33445 57468 33544
rect 57790 33464 57796 33516
rect 57848 33504 57854 33516
rect 57885 33507 57943 33513
rect 57885 33504 57897 33507
rect 57848 33476 57897 33504
rect 57848 33464 57854 33476
rect 57885 33473 57897 33476
rect 57931 33473 57943 33507
rect 57885 33467 57943 33473
rect 58069 33507 58127 33513
rect 58069 33473 58081 33507
rect 58115 33473 58127 33507
rect 58069 33467 58127 33473
rect 58529 33507 58587 33513
rect 58529 33473 58541 33507
rect 58575 33504 58587 33507
rect 58575 33476 58940 33504
rect 58575 33473 58587 33476
rect 58529 33467 58587 33473
rect 57425 33439 57483 33445
rect 57425 33405 57437 33439
rect 57471 33405 57483 33439
rect 57425 33399 57483 33405
rect 57514 33396 57520 33448
rect 57572 33396 57578 33448
rect 57698 33396 57704 33448
rect 57756 33436 57762 33448
rect 58084 33436 58112 33467
rect 57756 33408 58112 33436
rect 57756 33396 57762 33408
rect 58912 33380 58940 33476
rect 58345 33371 58403 33377
rect 58345 33368 58357 33371
rect 57348 33340 58357 33368
rect 9766 33300 9772 33312
rect 9692 33272 9772 33300
rect 9171 33269 9183 33272
rect 9125 33263 9183 33269
rect 9766 33260 9772 33272
rect 9824 33300 9830 33312
rect 10410 33300 10416 33312
rect 9824 33272 10416 33300
rect 9824 33260 9830 33272
rect 10410 33260 10416 33272
rect 10468 33300 10474 33312
rect 10597 33303 10655 33309
rect 10597 33300 10609 33303
rect 10468 33272 10609 33300
rect 10468 33260 10474 33272
rect 10597 33269 10609 33272
rect 10643 33269 10655 33303
rect 10597 33263 10655 33269
rect 43257 33303 43315 33309
rect 43257 33269 43269 33303
rect 43303 33300 43315 33303
rect 44818 33300 44824 33312
rect 43303 33272 44824 33300
rect 43303 33269 43315 33272
rect 43257 33263 43315 33269
rect 44818 33260 44824 33272
rect 44876 33260 44882 33312
rect 50890 33260 50896 33312
rect 50948 33260 50954 33312
rect 50982 33260 50988 33312
rect 51040 33300 51046 33312
rect 51828 33309 51856 33340
rect 58345 33337 58357 33340
rect 58391 33337 58403 33371
rect 58345 33331 58403 33337
rect 58894 33328 58900 33380
rect 58952 33328 58958 33380
rect 51813 33303 51871 33309
rect 51813 33300 51825 33303
rect 51040 33272 51825 33300
rect 51040 33260 51046 33272
rect 51813 33269 51825 33272
rect 51859 33269 51871 33303
rect 51813 33263 51871 33269
rect 52549 33303 52607 33309
rect 52549 33269 52561 33303
rect 52595 33300 52607 33303
rect 52638 33300 52644 33312
rect 52595 33272 52644 33300
rect 52595 33269 52607 33272
rect 52549 33263 52607 33269
rect 52638 33260 52644 33272
rect 52696 33260 52702 33312
rect 55490 33260 55496 33312
rect 55548 33260 55554 33312
rect 56962 33260 56968 33312
rect 57020 33260 57026 33312
rect 57330 33260 57336 33312
rect 57388 33300 57394 33312
rect 57977 33303 58035 33309
rect 57977 33300 57989 33303
rect 57388 33272 57989 33300
rect 57388 33260 57394 33272
rect 57977 33269 57989 33272
rect 58023 33269 58035 33303
rect 57977 33263 58035 33269
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 7558 33056 7564 33108
rect 7616 33096 7622 33108
rect 7745 33099 7803 33105
rect 7745 33096 7757 33099
rect 7616 33068 7757 33096
rect 7616 33056 7622 33068
rect 7745 33065 7757 33068
rect 7791 33065 7803 33099
rect 7745 33059 7803 33065
rect 38378 33056 38384 33108
rect 38436 33096 38442 33108
rect 44082 33096 44088 33108
rect 38436 33068 44088 33096
rect 38436 33056 38442 33068
rect 44082 33056 44088 33068
rect 44140 33056 44146 33108
rect 44266 33056 44272 33108
rect 44324 33096 44330 33108
rect 45925 33099 45983 33105
rect 44324 33068 44588 33096
rect 44324 33056 44330 33068
rect 42061 33031 42119 33037
rect 42061 32997 42073 33031
rect 42107 33028 42119 33031
rect 43254 33028 43260 33040
rect 42107 33000 43260 33028
rect 42107 32997 42119 33000
rect 42061 32991 42119 32997
rect 43254 32988 43260 33000
rect 43312 32988 43318 33040
rect 44560 33037 44588 33068
rect 45925 33065 45937 33099
rect 45971 33096 45983 33099
rect 46014 33096 46020 33108
rect 45971 33068 46020 33096
rect 45971 33065 45983 33068
rect 45925 33059 45983 33065
rect 46014 33056 46020 33068
rect 46072 33056 46078 33108
rect 46106 33056 46112 33108
rect 46164 33096 46170 33108
rect 46201 33099 46259 33105
rect 46201 33096 46213 33099
rect 46164 33068 46213 33096
rect 46164 33056 46170 33068
rect 46201 33065 46213 33068
rect 46247 33096 46259 33099
rect 46474 33096 46480 33108
rect 46247 33068 46480 33096
rect 46247 33065 46259 33068
rect 46201 33059 46259 33065
rect 46474 33056 46480 33068
rect 46532 33056 46538 33108
rect 47854 33056 47860 33108
rect 47912 33096 47918 33108
rect 48133 33099 48191 33105
rect 48133 33096 48145 33099
rect 47912 33068 48145 33096
rect 47912 33056 47918 33068
rect 48133 33065 48145 33068
rect 48179 33065 48191 33099
rect 48133 33059 48191 33065
rect 49344 33068 49556 33096
rect 44545 33031 44603 33037
rect 44545 32997 44557 33031
rect 44591 33028 44603 33031
rect 45097 33031 45155 33037
rect 45097 33028 45109 33031
rect 44591 33000 45109 33028
rect 44591 32997 44603 33000
rect 44545 32991 44603 32997
rect 45097 32997 45109 33000
rect 45143 32997 45155 33031
rect 45097 32991 45155 32997
rect 48041 33031 48099 33037
rect 48041 32997 48053 33031
rect 48087 33028 48099 33031
rect 49344 33028 49372 33068
rect 48087 33000 49372 33028
rect 49421 33031 49479 33037
rect 48087 32997 48099 33000
rect 48041 32991 48099 32997
rect 49421 32997 49433 33031
rect 49467 32997 49479 33031
rect 49421 32991 49479 32997
rect 6454 32920 6460 32972
rect 6512 32960 6518 32972
rect 6822 32960 6828 32972
rect 6512 32932 6828 32960
rect 6512 32920 6518 32932
rect 6822 32920 6828 32932
rect 6880 32960 6886 32972
rect 40313 32963 40371 32969
rect 6880 32932 7788 32960
rect 6880 32920 6886 32932
rect 2593 32895 2651 32901
rect 2593 32892 2605 32895
rect 2332 32864 2605 32892
rect 934 32784 940 32836
rect 992 32824 998 32836
rect 1581 32827 1639 32833
rect 1581 32824 1593 32827
rect 992 32796 1593 32824
rect 992 32784 998 32796
rect 1581 32793 1593 32796
rect 1627 32793 1639 32827
rect 1581 32787 1639 32793
rect 1394 32716 1400 32768
rect 1452 32756 1458 32768
rect 2332 32756 2360 32864
rect 2593 32861 2605 32864
rect 2639 32892 2651 32895
rect 2869 32895 2927 32901
rect 2869 32892 2881 32895
rect 2639 32864 2881 32892
rect 2639 32861 2651 32864
rect 2593 32855 2651 32861
rect 2869 32861 2881 32864
rect 2915 32861 2927 32895
rect 2869 32855 2927 32861
rect 7098 32852 7104 32904
rect 7156 32892 7162 32904
rect 7760 32901 7788 32932
rect 40313 32929 40325 32963
rect 40359 32960 40371 32963
rect 41598 32960 41604 32972
rect 40359 32932 41604 32960
rect 40359 32929 40371 32932
rect 40313 32923 40371 32929
rect 41598 32920 41604 32932
rect 41656 32920 41662 32972
rect 44177 32963 44235 32969
rect 44177 32960 44189 32963
rect 42904 32932 44189 32960
rect 42904 32904 42932 32932
rect 44177 32929 44189 32932
rect 44223 32929 44235 32963
rect 44350 32963 44408 32969
rect 44350 32960 44362 32963
rect 44177 32923 44235 32929
rect 44284 32932 44362 32960
rect 7469 32895 7527 32901
rect 7469 32892 7481 32895
rect 7156 32864 7481 32892
rect 7156 32852 7162 32864
rect 7469 32861 7481 32864
rect 7515 32861 7527 32895
rect 7469 32855 7527 32861
rect 7745 32895 7803 32901
rect 7745 32861 7757 32895
rect 7791 32892 7803 32895
rect 7834 32892 7840 32904
rect 7791 32864 7840 32892
rect 7791 32861 7803 32864
rect 7745 32855 7803 32861
rect 7834 32852 7840 32864
rect 7892 32852 7898 32904
rect 42610 32892 42616 32904
rect 41722 32878 42616 32892
rect 41708 32864 42616 32878
rect 40586 32784 40592 32836
rect 40644 32784 40650 32836
rect 1452 32728 2360 32756
rect 1452 32716 1458 32728
rect 3510 32716 3516 32768
rect 3568 32716 3574 32768
rect 4798 32716 4804 32768
rect 4856 32756 4862 32768
rect 4893 32759 4951 32765
rect 4893 32756 4905 32759
rect 4856 32728 4905 32756
rect 4856 32716 4862 32728
rect 4893 32725 4905 32728
rect 4939 32756 4951 32759
rect 5813 32759 5871 32765
rect 5813 32756 5825 32759
rect 4939 32728 5825 32756
rect 4939 32725 4951 32728
rect 4893 32719 4951 32725
rect 5813 32725 5825 32728
rect 5859 32756 5871 32759
rect 6362 32756 6368 32768
rect 5859 32728 6368 32756
rect 5859 32725 5871 32728
rect 5813 32719 5871 32725
rect 6362 32716 6368 32728
rect 6420 32756 6426 32768
rect 6733 32759 6791 32765
rect 6733 32756 6745 32759
rect 6420 32728 6745 32756
rect 6420 32716 6426 32728
rect 6733 32725 6745 32728
rect 6779 32756 6791 32759
rect 7282 32756 7288 32768
rect 6779 32728 7288 32756
rect 6779 32725 6791 32728
rect 6733 32719 6791 32725
rect 7282 32716 7288 32728
rect 7340 32716 7346 32768
rect 7374 32716 7380 32768
rect 7432 32756 7438 32768
rect 7561 32759 7619 32765
rect 7561 32756 7573 32759
rect 7432 32728 7573 32756
rect 7432 32716 7438 32728
rect 7561 32725 7573 32728
rect 7607 32725 7619 32759
rect 7561 32719 7619 32725
rect 41414 32716 41420 32768
rect 41472 32756 41478 32768
rect 41708 32756 41736 32864
rect 42610 32852 42616 32864
rect 42668 32852 42674 32904
rect 42702 32852 42708 32904
rect 42760 32852 42766 32904
rect 42886 32852 42892 32904
rect 42944 32852 42950 32904
rect 43254 32852 43260 32904
rect 43312 32892 43318 32904
rect 43530 32892 43536 32904
rect 43312 32864 43536 32892
rect 43312 32852 43318 32864
rect 43530 32852 43536 32864
rect 43588 32852 43594 32904
rect 43714 32852 43720 32904
rect 43772 32892 43778 32904
rect 44284 32892 44312 32932
rect 44350 32929 44362 32932
rect 44396 32929 44408 32963
rect 49436 32960 49464 32991
rect 44350 32923 44408 32929
rect 49068 32932 49464 32960
rect 49528 32960 49556 33068
rect 55582 33056 55588 33108
rect 55640 33056 55646 33108
rect 56594 33056 56600 33108
rect 56652 33056 56658 33108
rect 57333 33099 57391 33105
rect 57333 33065 57345 33099
rect 57379 33096 57391 33099
rect 57698 33096 57704 33108
rect 57379 33068 57704 33096
rect 57379 33065 57391 33068
rect 57333 33059 57391 33065
rect 57698 33056 57704 33068
rect 57756 33056 57762 33108
rect 50798 32988 50804 33040
rect 50856 32988 50862 33040
rect 50816 32960 50844 32988
rect 49528 32932 50844 32960
rect 55600 32960 55628 33056
rect 56413 33031 56471 33037
rect 56413 32997 56425 33031
rect 56459 33028 56471 33031
rect 56502 33028 56508 33040
rect 56459 33000 56508 33028
rect 56459 32997 56471 33000
rect 56413 32991 56471 32997
rect 56502 32988 56508 33000
rect 56560 32988 56566 33040
rect 56612 33028 56640 33056
rect 57882 33028 57888 33040
rect 56612 33000 57888 33028
rect 55600 32932 56640 32960
rect 43772 32864 44312 32892
rect 43772 32852 43778 32864
rect 44634 32852 44640 32904
rect 44692 32852 44698 32904
rect 44818 32852 44824 32904
rect 44876 32892 44882 32904
rect 45005 32895 45063 32901
rect 45005 32892 45017 32895
rect 44876 32864 45017 32892
rect 44876 32852 44882 32864
rect 45005 32861 45017 32864
rect 45051 32861 45063 32895
rect 45005 32855 45063 32861
rect 45281 32895 45339 32901
rect 45281 32861 45293 32895
rect 45327 32861 45339 32895
rect 45281 32855 45339 32861
rect 42794 32784 42800 32836
rect 42852 32824 42858 32836
rect 43625 32827 43683 32833
rect 43625 32824 43637 32827
rect 42852 32796 43637 32824
rect 42852 32784 42858 32796
rect 43625 32793 43637 32796
rect 43671 32793 43683 32827
rect 43625 32787 43683 32793
rect 43806 32784 43812 32836
rect 43864 32824 43870 32836
rect 44361 32827 44419 32833
rect 44361 32824 44373 32827
rect 43864 32796 44373 32824
rect 43864 32784 43870 32796
rect 44361 32793 44373 32796
rect 44407 32793 44419 32827
rect 44361 32787 44419 32793
rect 44450 32784 44456 32836
rect 44508 32824 44514 32836
rect 45296 32824 45324 32855
rect 47670 32852 47676 32904
rect 47728 32892 47734 32904
rect 47857 32895 47915 32901
rect 47857 32892 47869 32895
rect 47728 32864 47869 32892
rect 47728 32852 47734 32864
rect 47857 32861 47869 32864
rect 47903 32861 47915 32895
rect 47857 32855 47915 32861
rect 48041 32895 48099 32901
rect 48041 32861 48053 32895
rect 48087 32892 48099 32895
rect 48314 32892 48320 32904
rect 48087 32864 48320 32892
rect 48087 32861 48099 32864
rect 48041 32855 48099 32861
rect 48314 32852 48320 32864
rect 48372 32852 48378 32904
rect 49068 32901 49096 32932
rect 48777 32895 48835 32901
rect 48777 32861 48789 32895
rect 48823 32892 48835 32895
rect 48869 32895 48927 32901
rect 48869 32892 48881 32895
rect 48823 32864 48881 32892
rect 48823 32861 48835 32864
rect 48777 32855 48835 32861
rect 48869 32861 48881 32864
rect 48915 32861 48927 32895
rect 48869 32855 48927 32861
rect 49053 32895 49111 32901
rect 49053 32861 49065 32895
rect 49099 32861 49111 32895
rect 49053 32855 49111 32861
rect 49234 32852 49240 32904
rect 49292 32852 49298 32904
rect 49329 32895 49387 32901
rect 49329 32861 49341 32895
rect 49375 32892 49387 32895
rect 49528 32892 49556 32932
rect 49375 32864 49556 32892
rect 49697 32895 49755 32901
rect 49375 32861 49387 32864
rect 49329 32855 49387 32861
rect 49697 32861 49709 32895
rect 49743 32892 49755 32895
rect 49973 32895 50031 32901
rect 49973 32892 49985 32895
rect 49743 32864 49985 32892
rect 49743 32861 49755 32864
rect 49697 32855 49755 32861
rect 49973 32861 49985 32864
rect 50019 32892 50031 32895
rect 50430 32892 50436 32904
rect 50019 32864 50436 32892
rect 50019 32861 50031 32864
rect 49973 32855 50031 32861
rect 50430 32852 50436 32864
rect 50488 32852 50494 32904
rect 50982 32852 50988 32904
rect 51040 32852 51046 32904
rect 56321 32895 56379 32901
rect 56321 32861 56333 32895
rect 56367 32861 56379 32895
rect 56321 32855 56379 32861
rect 44508 32796 45324 32824
rect 44508 32784 44514 32796
rect 48958 32784 48964 32836
rect 49016 32824 49022 32836
rect 49421 32827 49479 32833
rect 49421 32824 49433 32827
rect 49016 32796 49433 32824
rect 49016 32784 49022 32796
rect 49421 32793 49433 32796
rect 49467 32793 49479 32827
rect 49421 32787 49479 32793
rect 49605 32827 49663 32833
rect 49605 32793 49617 32827
rect 49651 32824 49663 32827
rect 51000 32824 51028 32852
rect 49651 32796 51028 32824
rect 56336 32824 56364 32855
rect 56410 32852 56416 32904
rect 56468 32892 56474 32904
rect 56612 32901 56640 32932
rect 56505 32895 56563 32901
rect 56505 32892 56517 32895
rect 56468 32864 56517 32892
rect 56468 32852 56474 32864
rect 56505 32861 56517 32864
rect 56551 32861 56563 32895
rect 56505 32855 56563 32861
rect 56597 32895 56655 32901
rect 56597 32861 56609 32895
rect 56643 32861 56655 32895
rect 56597 32855 56655 32861
rect 56781 32895 56839 32901
rect 56781 32861 56793 32895
rect 56827 32861 56839 32895
rect 56781 32855 56839 32861
rect 56689 32827 56747 32833
rect 56689 32824 56701 32827
rect 56336 32796 56701 32824
rect 49651 32793 49663 32796
rect 49605 32787 49663 32793
rect 56689 32793 56701 32796
rect 56735 32793 56747 32827
rect 56796 32824 56824 32855
rect 56962 32852 56968 32904
rect 57020 32892 57026 32904
rect 57241 32895 57299 32901
rect 57241 32892 57253 32895
rect 57020 32864 57253 32892
rect 57020 32852 57026 32864
rect 57241 32861 57253 32864
rect 57287 32861 57299 32895
rect 57241 32855 57299 32861
rect 57330 32852 57336 32904
rect 57388 32852 57394 32904
rect 57440 32901 57468 33000
rect 57882 32988 57888 33000
rect 57940 32988 57946 33040
rect 57425 32895 57483 32901
rect 57425 32861 57437 32895
rect 57471 32861 57483 32895
rect 57425 32855 57483 32861
rect 58529 32895 58587 32901
rect 58529 32861 58541 32895
rect 58575 32892 58587 32895
rect 58575 32864 58940 32892
rect 58575 32861 58587 32864
rect 58529 32855 58587 32861
rect 57348 32824 57376 32852
rect 58912 32836 58940 32864
rect 56796 32796 57376 32824
rect 56689 32787 56747 32793
rect 58894 32784 58900 32836
rect 58952 32784 58958 32836
rect 41472 32728 41736 32756
rect 41472 32716 41478 32728
rect 42150 32716 42156 32768
rect 42208 32716 42214 32768
rect 42889 32759 42947 32765
rect 42889 32725 42901 32759
rect 42935 32756 42947 32759
rect 43070 32756 43076 32768
rect 42935 32728 43076 32756
rect 42935 32725 42947 32728
rect 42889 32719 42947 32725
rect 43070 32716 43076 32728
rect 43128 32716 43134 32768
rect 43530 32716 43536 32768
rect 43588 32756 43594 32768
rect 44726 32756 44732 32768
rect 43588 32728 44732 32756
rect 43588 32716 43594 32728
rect 44726 32716 44732 32728
rect 44784 32716 44790 32768
rect 49878 32716 49884 32768
rect 49936 32716 49942 32768
rect 51258 32716 51264 32768
rect 51316 32756 51322 32768
rect 51534 32756 51540 32768
rect 51316 32728 51540 32756
rect 51316 32716 51322 32728
rect 51534 32716 51540 32728
rect 51592 32716 51598 32768
rect 52730 32716 52736 32768
rect 52788 32756 52794 32768
rect 56778 32756 56784 32768
rect 52788 32728 56784 32756
rect 52788 32716 52794 32728
rect 56778 32716 56784 32728
rect 56836 32716 56842 32768
rect 58345 32759 58403 32765
rect 58345 32725 58357 32759
rect 58391 32756 58403 32759
rect 58391 32728 58940 32756
rect 58391 32725 58403 32728
rect 58345 32719 58403 32725
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 1394 32512 1400 32564
rect 1452 32512 1458 32564
rect 2866 32512 2872 32564
rect 2924 32552 2930 32564
rect 3973 32555 4031 32561
rect 3973 32552 3985 32555
rect 2924 32524 3985 32552
rect 2924 32512 2930 32524
rect 3973 32521 3985 32524
rect 4019 32521 4031 32555
rect 3973 32515 4031 32521
rect 4801 32555 4859 32561
rect 4801 32521 4813 32555
rect 4847 32521 4859 32555
rect 4801 32515 4859 32521
rect 2406 32444 2412 32496
rect 2464 32444 2470 32496
rect 4816 32484 4844 32515
rect 7282 32512 7288 32564
rect 7340 32552 7346 32564
rect 7466 32552 7472 32564
rect 7340 32524 7472 32552
rect 7340 32512 7346 32524
rect 7466 32512 7472 32524
rect 7524 32552 7530 32564
rect 8113 32555 8171 32561
rect 8113 32552 8125 32555
rect 7524 32524 8125 32552
rect 7524 32512 7530 32524
rect 8113 32521 8125 32524
rect 8159 32552 8171 32555
rect 8159 32524 8432 32552
rect 8159 32521 8171 32524
rect 8113 32515 8171 32521
rect 8404 32484 8432 32524
rect 8570 32512 8576 32564
rect 8628 32552 8634 32564
rect 9306 32552 9312 32564
rect 8628 32524 9312 32552
rect 8628 32512 8634 32524
rect 9306 32512 9312 32524
rect 9364 32512 9370 32564
rect 38378 32512 38384 32564
rect 38436 32512 38442 32564
rect 40586 32512 40592 32564
rect 40644 32552 40650 32564
rect 41325 32555 41383 32561
rect 41325 32552 41337 32555
rect 40644 32524 41337 32552
rect 40644 32512 40650 32524
rect 41325 32521 41337 32524
rect 41371 32521 41383 32555
rect 41325 32515 41383 32521
rect 42150 32512 42156 32564
rect 42208 32512 42214 32564
rect 42429 32555 42487 32561
rect 42429 32521 42441 32555
rect 42475 32552 42487 32555
rect 42702 32552 42708 32564
rect 42475 32524 42708 32552
rect 42475 32521 42487 32524
rect 42429 32515 42487 32521
rect 42702 32512 42708 32524
rect 42760 32512 42766 32564
rect 42794 32512 42800 32564
rect 42852 32512 42858 32564
rect 42886 32512 42892 32564
rect 42944 32512 42950 32564
rect 44266 32552 44272 32564
rect 44192 32524 44272 32552
rect 10318 32484 10324 32496
rect 4172 32456 4844 32484
rect 4908 32456 8248 32484
rect 4172 32425 4200 32456
rect 4540 32425 4568 32456
rect 3973 32419 4031 32425
rect 3973 32385 3985 32419
rect 4019 32385 4031 32419
rect 3973 32379 4031 32385
rect 4157 32419 4215 32425
rect 4157 32385 4169 32419
rect 4203 32385 4215 32419
rect 4157 32379 4215 32385
rect 4249 32419 4307 32425
rect 4249 32385 4261 32419
rect 4295 32385 4307 32419
rect 4249 32379 4307 32385
rect 4433 32419 4491 32425
rect 4433 32385 4445 32419
rect 4479 32385 4491 32419
rect 4433 32379 4491 32385
rect 4525 32419 4583 32425
rect 4525 32385 4537 32419
rect 4571 32385 4583 32419
rect 4525 32379 4583 32385
rect 4709 32419 4767 32425
rect 4709 32385 4721 32419
rect 4755 32416 4767 32419
rect 4798 32416 4804 32428
rect 4755 32388 4804 32416
rect 4755 32385 4767 32388
rect 4709 32379 4767 32385
rect 2866 32308 2872 32360
rect 2924 32308 2930 32360
rect 3142 32308 3148 32360
rect 3200 32348 3206 32360
rect 3200 32320 3372 32348
rect 3200 32308 3206 32320
rect 2498 32172 2504 32224
rect 2556 32212 2562 32224
rect 3237 32215 3295 32221
rect 3237 32212 3249 32215
rect 2556 32184 3249 32212
rect 2556 32172 2562 32184
rect 3237 32181 3249 32184
rect 3283 32181 3295 32215
rect 3344 32212 3372 32320
rect 3786 32308 3792 32360
rect 3844 32308 3850 32360
rect 3878 32308 3884 32360
rect 3936 32348 3942 32360
rect 3988 32348 4016 32379
rect 4264 32348 4292 32379
rect 3936 32320 4292 32348
rect 4448 32348 4476 32379
rect 4798 32376 4804 32388
rect 4856 32376 4862 32428
rect 4908 32348 4936 32456
rect 8220 32425 8248 32456
rect 8404 32456 10324 32484
rect 8404 32425 8432 32456
rect 10318 32444 10324 32456
rect 10376 32484 10382 32496
rect 12434 32484 12440 32496
rect 10376 32456 12440 32484
rect 10376 32444 10382 32456
rect 12434 32444 12440 32456
rect 12492 32444 12498 32496
rect 5914 32419 5972 32425
rect 5914 32416 5926 32419
rect 4448 32320 4936 32348
rect 5000 32388 5926 32416
rect 3936 32308 3942 32320
rect 3418 32240 3424 32292
rect 3476 32280 3482 32292
rect 3476 32252 4384 32280
rect 3476 32240 3482 32252
rect 4062 32212 4068 32224
rect 3344 32184 4068 32212
rect 3237 32175 3295 32181
rect 4062 32172 4068 32184
rect 4120 32172 4126 32224
rect 4356 32221 4384 32252
rect 5000 32224 5028 32388
rect 5914 32385 5926 32388
rect 5960 32385 5972 32419
rect 5914 32379 5972 32385
rect 8205 32419 8263 32425
rect 8205 32385 8217 32419
rect 8251 32385 8263 32419
rect 8205 32379 8263 32385
rect 8389 32419 8447 32425
rect 8389 32385 8401 32419
rect 8435 32385 8447 32419
rect 8389 32379 8447 32385
rect 8481 32419 8539 32425
rect 8481 32385 8493 32419
rect 8527 32416 8539 32419
rect 8757 32419 8815 32425
rect 8527 32388 8616 32416
rect 8527 32385 8539 32388
rect 8481 32379 8539 32385
rect 6181 32351 6239 32357
rect 6181 32317 6193 32351
rect 6227 32348 6239 32351
rect 6227 32320 6684 32348
rect 6227 32317 6239 32320
rect 6181 32311 6239 32317
rect 4341 32215 4399 32221
rect 4341 32181 4353 32215
rect 4387 32181 4399 32215
rect 4341 32175 4399 32181
rect 4614 32172 4620 32224
rect 4672 32172 4678 32224
rect 4982 32172 4988 32224
rect 5040 32172 5046 32224
rect 6656 32221 6684 32320
rect 6641 32215 6699 32221
rect 6641 32181 6653 32215
rect 6687 32212 6699 32215
rect 7834 32212 7840 32224
rect 6687 32184 7840 32212
rect 6687 32181 6699 32184
rect 6641 32175 6699 32181
rect 7834 32172 7840 32184
rect 7892 32172 7898 32224
rect 8220 32212 8248 32379
rect 8297 32283 8355 32289
rect 8297 32249 8309 32283
rect 8343 32280 8355 32283
rect 8588 32280 8616 32388
rect 8757 32385 8769 32419
rect 8803 32416 8815 32419
rect 8846 32416 8852 32428
rect 8803 32388 8852 32416
rect 8803 32385 8815 32388
rect 8757 32379 8815 32385
rect 8846 32376 8852 32388
rect 8904 32376 8910 32428
rect 9962 32419 10020 32425
rect 9962 32416 9974 32419
rect 9232 32388 9974 32416
rect 9232 32348 9260 32388
rect 9962 32385 9974 32388
rect 10008 32385 10020 32419
rect 9962 32379 10020 32385
rect 39022 32376 39028 32428
rect 39080 32376 39086 32428
rect 39206 32376 39212 32428
rect 39264 32376 39270 32428
rect 39301 32419 39359 32425
rect 39301 32385 39313 32419
rect 39347 32416 39359 32419
rect 39347 32388 39436 32416
rect 39347 32385 39359 32388
rect 39301 32379 39359 32385
rect 8772 32320 9260 32348
rect 8772 32289 8800 32320
rect 10226 32308 10232 32360
rect 10284 32348 10290 32360
rect 10284 32320 10640 32348
rect 10284 32308 10290 32320
rect 8343 32252 8616 32280
rect 8757 32283 8815 32289
rect 8343 32249 8355 32252
rect 8297 32243 8355 32249
rect 8757 32249 8769 32283
rect 8803 32249 8815 32283
rect 8757 32243 8815 32249
rect 10612 32221 10640 32320
rect 39408 32280 39436 32388
rect 39482 32376 39488 32428
rect 39540 32376 39546 32428
rect 41509 32419 41567 32425
rect 41509 32385 41521 32419
rect 41555 32416 41567 32419
rect 42168 32416 42196 32512
rect 42812 32425 42840 32512
rect 43714 32484 43720 32496
rect 42904 32456 43720 32484
rect 42904 32428 42932 32456
rect 43714 32444 43720 32456
rect 43772 32444 43778 32496
rect 43806 32444 43812 32496
rect 43864 32484 43870 32496
rect 44192 32493 44220 32524
rect 44266 32512 44272 32524
rect 44324 32512 44330 32564
rect 44376 32524 44680 32552
rect 44085 32487 44143 32493
rect 44085 32484 44097 32487
rect 43864 32456 44097 32484
rect 43864 32444 43870 32456
rect 44085 32453 44097 32456
rect 44131 32453 44143 32487
rect 44085 32447 44143 32453
rect 44177 32487 44235 32493
rect 44177 32453 44189 32487
rect 44223 32453 44235 32487
rect 44376 32484 44404 32524
rect 44177 32447 44235 32453
rect 44284 32456 44404 32484
rect 41555 32388 42196 32416
rect 42613 32419 42671 32425
rect 41555 32385 41567 32388
rect 41509 32379 41567 32385
rect 42613 32385 42625 32419
rect 42659 32385 42671 32419
rect 42613 32379 42671 32385
rect 42797 32419 42855 32425
rect 42797 32385 42809 32419
rect 42843 32385 42855 32419
rect 42797 32379 42855 32385
rect 40586 32308 40592 32360
rect 40644 32308 40650 32360
rect 42058 32308 42064 32360
rect 42116 32348 42122 32360
rect 42628 32348 42656 32379
rect 42886 32376 42892 32428
rect 42944 32376 42950 32428
rect 43070 32376 43076 32428
rect 43128 32376 43134 32428
rect 44284 32425 44312 32456
rect 44542 32444 44548 32496
rect 44600 32444 44606 32496
rect 44652 32484 44680 32524
rect 44910 32512 44916 32564
rect 44968 32552 44974 32564
rect 44968 32524 45324 32552
rect 44968 32512 44974 32524
rect 45189 32487 45247 32493
rect 45189 32484 45201 32487
rect 44652 32456 45201 32484
rect 45189 32453 45201 32456
rect 45235 32453 45247 32487
rect 45189 32447 45247 32453
rect 43901 32419 43959 32425
rect 43901 32385 43913 32419
rect 43947 32385 43959 32419
rect 43901 32379 43959 32385
rect 44269 32419 44327 32425
rect 44269 32385 44281 32419
rect 44315 32385 44327 32419
rect 44821 32419 44879 32425
rect 44821 32416 44833 32419
rect 44269 32379 44327 32385
rect 44376 32414 44588 32416
rect 44652 32414 44833 32416
rect 44376 32388 44833 32414
rect 42116 32320 42656 32348
rect 43088 32348 43116 32376
rect 43622 32348 43628 32360
rect 43088 32320 43628 32348
rect 42116 32308 42122 32320
rect 43622 32308 43628 32320
rect 43680 32308 43686 32360
rect 43916 32348 43944 32379
rect 44174 32348 44180 32360
rect 43916 32320 44180 32348
rect 44174 32308 44180 32320
rect 44232 32348 44238 32360
rect 44376 32348 44404 32388
rect 44560 32386 44680 32388
rect 44821 32385 44833 32388
rect 44867 32416 44879 32419
rect 44910 32416 44916 32428
rect 44867 32388 44916 32416
rect 44867 32385 44879 32388
rect 44821 32379 44879 32385
rect 44910 32376 44916 32388
rect 44968 32376 44974 32428
rect 45296 32425 45324 32524
rect 45646 32512 45652 32564
rect 45704 32552 45710 32564
rect 52730 32552 52736 32564
rect 45704 32524 52736 32552
rect 45704 32512 45710 32524
rect 52730 32512 52736 32524
rect 52788 32512 52794 32564
rect 55122 32552 55128 32564
rect 52840 32524 55128 32552
rect 46658 32444 46664 32496
rect 46716 32444 46722 32496
rect 49878 32484 49884 32496
rect 48884 32456 49884 32484
rect 45097 32420 45155 32425
rect 45020 32419 45155 32420
rect 45020 32392 45109 32419
rect 44232 32320 44404 32348
rect 44637 32351 44695 32357
rect 44232 32308 44238 32320
rect 44637 32317 44649 32351
rect 44683 32348 44695 32351
rect 45020 32348 45048 32392
rect 45097 32385 45109 32392
rect 45143 32385 45155 32419
rect 45097 32379 45155 32385
rect 45281 32419 45339 32425
rect 45281 32385 45293 32419
rect 45327 32416 45339 32419
rect 45462 32416 45468 32428
rect 45327 32388 45468 32416
rect 45327 32385 45339 32388
rect 45281 32379 45339 32385
rect 45462 32376 45468 32388
rect 45520 32376 45526 32428
rect 47394 32376 47400 32428
rect 47452 32376 47458 32428
rect 47670 32376 47676 32428
rect 47728 32416 47734 32428
rect 48884 32425 48912 32456
rect 49878 32444 49884 32456
rect 49936 32444 49942 32496
rect 47857 32419 47915 32425
rect 47857 32416 47869 32419
rect 47728 32388 47869 32416
rect 47728 32376 47734 32388
rect 47857 32385 47869 32388
rect 47903 32385 47915 32419
rect 47857 32379 47915 32385
rect 48869 32419 48927 32425
rect 48869 32385 48881 32419
rect 48915 32385 48927 32419
rect 48869 32379 48927 32385
rect 49053 32419 49111 32425
rect 49053 32385 49065 32419
rect 49099 32416 49111 32419
rect 49234 32416 49240 32428
rect 49099 32388 49240 32416
rect 49099 32385 49111 32388
rect 49053 32379 49111 32385
rect 49234 32376 49240 32388
rect 49292 32376 49298 32428
rect 52840 32425 52868 32524
rect 55122 32512 55128 32524
rect 55180 32512 55186 32564
rect 53742 32444 53748 32496
rect 53800 32484 53806 32496
rect 58253 32487 58311 32493
rect 58253 32484 58265 32487
rect 53800 32456 58265 32484
rect 53800 32444 53806 32456
rect 58253 32453 58265 32456
rect 58299 32453 58311 32487
rect 58253 32447 58311 32453
rect 52825 32419 52883 32425
rect 52825 32385 52837 32419
rect 52871 32385 52883 32419
rect 52825 32379 52883 32385
rect 53009 32419 53067 32425
rect 53009 32385 53021 32419
rect 53055 32416 53067 32419
rect 53190 32416 53196 32428
rect 53055 32388 53196 32416
rect 53055 32385 53067 32388
rect 53009 32379 53067 32385
rect 53190 32376 53196 32388
rect 53248 32416 53254 32428
rect 53837 32419 53895 32425
rect 53837 32416 53849 32419
rect 53248 32388 53849 32416
rect 53248 32376 53254 32388
rect 53837 32385 53849 32388
rect 53883 32385 53895 32419
rect 53837 32379 53895 32385
rect 58345 32419 58403 32425
rect 58345 32385 58357 32419
rect 58391 32416 58403 32419
rect 58912 32416 58940 32728
rect 58391 32388 58940 32416
rect 58391 32385 58403 32388
rect 58345 32379 58403 32385
rect 44683 32320 45048 32348
rect 44683 32317 44695 32320
rect 44637 32311 44695 32317
rect 39316 32252 39436 32280
rect 39316 32224 39344 32252
rect 44450 32240 44456 32292
rect 44508 32240 44514 32292
rect 44652 32224 44680 32311
rect 45554 32308 45560 32360
rect 45612 32348 45618 32360
rect 46658 32348 46664 32360
rect 45612 32320 46664 32348
rect 45612 32308 45618 32320
rect 46658 32308 46664 32320
rect 46716 32308 46722 32360
rect 47026 32308 47032 32360
rect 47084 32308 47090 32360
rect 47581 32351 47639 32357
rect 47581 32317 47593 32351
rect 47627 32317 47639 32351
rect 47581 32311 47639 32317
rect 52917 32351 52975 32357
rect 52917 32317 52929 32351
rect 52963 32348 52975 32351
rect 53653 32351 53711 32357
rect 53653 32348 53665 32351
rect 52963 32320 53665 32348
rect 52963 32317 52975 32320
rect 52917 32311 52975 32317
rect 53653 32317 53665 32320
rect 53699 32317 53711 32351
rect 53653 32311 53711 32317
rect 46198 32280 46204 32292
rect 45020 32252 46204 32280
rect 8849 32215 8907 32221
rect 8849 32212 8861 32215
rect 8220 32184 8861 32212
rect 8849 32181 8861 32184
rect 8895 32181 8907 32215
rect 8849 32175 8907 32181
rect 10597 32215 10655 32221
rect 10597 32181 10609 32215
rect 10643 32212 10655 32215
rect 12342 32212 12348 32224
rect 10643 32184 12348 32212
rect 10643 32181 10655 32184
rect 10597 32175 10655 32181
rect 12342 32172 12348 32184
rect 12400 32172 12406 32224
rect 39117 32215 39175 32221
rect 39117 32181 39129 32215
rect 39163 32212 39175 32215
rect 39298 32212 39304 32224
rect 39163 32184 39304 32212
rect 39163 32181 39175 32184
rect 39117 32175 39175 32181
rect 39298 32172 39304 32184
rect 39356 32172 39362 32224
rect 39390 32172 39396 32224
rect 39448 32172 39454 32224
rect 41230 32172 41236 32224
rect 41288 32172 41294 32224
rect 44634 32172 44640 32224
rect 44692 32172 44698 32224
rect 44726 32172 44732 32224
rect 44784 32172 44790 32224
rect 45020 32221 45048 32252
rect 46198 32240 46204 32252
rect 46256 32240 46262 32292
rect 45005 32215 45063 32221
rect 45005 32181 45017 32215
rect 45051 32181 45063 32215
rect 45005 32175 45063 32181
rect 45554 32172 45560 32224
rect 45612 32221 45618 32224
rect 45612 32215 45661 32221
rect 45612 32181 45615 32215
rect 45649 32212 45661 32215
rect 47596 32212 47624 32311
rect 54386 32308 54392 32360
rect 54444 32308 54450 32360
rect 55582 32308 55588 32360
rect 55640 32308 55646 32360
rect 55490 32280 55496 32292
rect 51046 32252 55496 32280
rect 45649 32184 47624 32212
rect 48961 32215 49019 32221
rect 45649 32181 45661 32184
rect 45612 32175 45661 32181
rect 48961 32181 48973 32215
rect 49007 32212 49019 32215
rect 49050 32212 49056 32224
rect 49007 32184 49056 32212
rect 49007 32181 49019 32184
rect 48961 32175 49019 32181
rect 45612 32172 45618 32175
rect 49050 32172 49056 32184
rect 49108 32172 49114 32224
rect 49510 32172 49516 32224
rect 49568 32212 49574 32224
rect 51046 32212 51074 32252
rect 55490 32240 55496 32252
rect 55548 32240 55554 32292
rect 49568 32184 51074 32212
rect 49568 32172 49574 32184
rect 53098 32172 53104 32224
rect 53156 32172 53162 32224
rect 55030 32172 55036 32224
rect 55088 32172 55094 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 2148 31980 2820 32008
rect 2148 31813 2176 31980
rect 2317 31943 2375 31949
rect 2317 31909 2329 31943
rect 2363 31940 2375 31943
rect 2792 31940 2820 31980
rect 2866 31968 2872 32020
rect 2924 32008 2930 32020
rect 3329 32011 3387 32017
rect 3329 32008 3341 32011
rect 2924 31980 3341 32008
rect 2924 31968 2930 31980
rect 3329 31977 3341 31980
rect 3375 31977 3387 32011
rect 3329 31971 3387 31977
rect 3418 31968 3424 32020
rect 3476 31968 3482 32020
rect 3510 31968 3516 32020
rect 3568 31968 3574 32020
rect 4614 31968 4620 32020
rect 4672 31968 4678 32020
rect 4982 31968 4988 32020
rect 5040 31968 5046 32020
rect 6273 32011 6331 32017
rect 6273 31977 6285 32011
rect 6319 32008 6331 32011
rect 6362 32008 6368 32020
rect 6319 31980 6368 32008
rect 6319 31977 6331 31980
rect 6273 31971 6331 31977
rect 6362 31968 6368 31980
rect 6420 31968 6426 32020
rect 6457 32011 6515 32017
rect 6457 31977 6469 32011
rect 6503 32008 6515 32011
rect 6914 32008 6920 32020
rect 6503 31980 6920 32008
rect 6503 31977 6515 31980
rect 6457 31971 6515 31977
rect 6914 31968 6920 31980
rect 6972 31968 6978 32020
rect 7834 31968 7840 32020
rect 7892 32008 7898 32020
rect 8389 32011 8447 32017
rect 8389 32008 8401 32011
rect 7892 31980 8401 32008
rect 7892 31968 7898 31980
rect 8389 31977 8401 31980
rect 8435 32008 8447 32011
rect 10226 32008 10232 32020
rect 8435 31980 10232 32008
rect 8435 31977 8447 31980
rect 8389 31971 8447 31977
rect 3436 31940 3464 31968
rect 2363 31912 2728 31940
rect 2792 31912 3464 31940
rect 2363 31909 2375 31912
rect 2317 31903 2375 31909
rect 2409 31875 2467 31881
rect 2409 31841 2421 31875
rect 2455 31872 2467 31875
rect 2498 31872 2504 31884
rect 2455 31844 2504 31872
rect 2455 31841 2467 31844
rect 2409 31835 2467 31841
rect 2498 31832 2504 31844
rect 2556 31832 2562 31884
rect 2700 31881 2728 31912
rect 2685 31875 2743 31881
rect 2685 31841 2697 31875
rect 2731 31841 2743 31875
rect 2685 31835 2743 31841
rect 2133 31807 2191 31813
rect 2133 31773 2145 31807
rect 2179 31773 2191 31807
rect 2133 31767 2191 31773
rect 2225 31807 2283 31813
rect 2225 31773 2237 31807
rect 2271 31804 2283 31807
rect 3326 31804 3332 31816
rect 2271 31776 3332 31804
rect 2271 31773 2283 31776
rect 2225 31767 2283 31773
rect 3326 31764 3332 31776
rect 3384 31764 3390 31816
rect 3421 31807 3479 31813
rect 3421 31773 3433 31807
rect 3467 31804 3479 31807
rect 3528 31804 3556 31968
rect 3467 31776 3556 31804
rect 3605 31807 3663 31813
rect 3467 31773 3479 31776
rect 3421 31767 3479 31773
rect 3605 31773 3617 31807
rect 3651 31773 3663 31807
rect 4632 31804 4660 31968
rect 6641 31943 6699 31949
rect 6641 31940 6653 31943
rect 6288 31912 6653 31940
rect 4982 31832 4988 31884
rect 5040 31872 5046 31884
rect 5040 31844 5764 31872
rect 5040 31832 5046 31844
rect 4709 31807 4767 31813
rect 4709 31804 4721 31807
rect 4632 31776 4721 31804
rect 3605 31767 3663 31773
rect 4709 31773 4721 31776
rect 4755 31773 4767 31807
rect 4709 31767 4767 31773
rect 4801 31807 4859 31813
rect 4801 31773 4813 31807
rect 4847 31804 4859 31807
rect 4890 31804 4896 31816
rect 4847 31776 4896 31804
rect 4847 31773 4859 31776
rect 4801 31767 4859 31773
rect 3620 31736 3648 31767
rect 4890 31764 4896 31776
rect 4948 31804 4954 31816
rect 5258 31804 5264 31816
rect 4948 31776 5264 31804
rect 4948 31764 4954 31776
rect 5258 31764 5264 31776
rect 5316 31764 5322 31816
rect 5736 31804 5764 31844
rect 6288 31804 6316 31912
rect 6641 31909 6653 31912
rect 6687 31909 6699 31943
rect 6641 31903 6699 31909
rect 8021 31875 8079 31881
rect 8021 31841 8033 31875
rect 8067 31872 8079 31875
rect 8404 31872 8432 31971
rect 10226 31968 10232 31980
rect 10284 31968 10290 32020
rect 39390 32008 39396 32020
rect 39132 31980 39396 32008
rect 10321 31943 10379 31949
rect 10321 31909 10333 31943
rect 10367 31909 10379 31943
rect 10321 31903 10379 31909
rect 8067 31844 8432 31872
rect 10336 31872 10364 31903
rect 37734 31900 37740 31952
rect 37792 31940 37798 31952
rect 38289 31943 38347 31949
rect 38289 31940 38301 31943
rect 37792 31912 38301 31940
rect 37792 31900 37798 31912
rect 38289 31909 38301 31912
rect 38335 31909 38347 31943
rect 38289 31903 38347 31909
rect 10336 31844 10548 31872
rect 8067 31841 8079 31844
rect 8021 31835 8079 31841
rect 6355 31807 6413 31813
rect 6355 31804 6367 31807
rect 5736 31776 6367 31804
rect 6355 31773 6367 31776
rect 6401 31773 6413 31807
rect 6355 31767 6413 31773
rect 6454 31764 6460 31816
rect 6512 31804 6518 31816
rect 10520 31813 10548 31844
rect 38838 31832 38844 31884
rect 38896 31832 38902 31884
rect 6549 31807 6607 31813
rect 6549 31804 6561 31807
rect 6512 31776 6561 31804
rect 6512 31764 6518 31776
rect 6549 31773 6561 31776
rect 6595 31773 6607 31807
rect 6549 31767 6607 31773
rect 10045 31807 10103 31813
rect 10045 31773 10057 31807
rect 10091 31804 10103 31807
rect 10229 31807 10287 31813
rect 10229 31804 10241 31807
rect 10091 31776 10241 31804
rect 10091 31773 10103 31776
rect 10045 31767 10103 31773
rect 10229 31773 10241 31776
rect 10275 31804 10287 31807
rect 10505 31807 10563 31813
rect 10275 31776 10309 31804
rect 10275 31773 10287 31776
rect 10229 31767 10287 31773
rect 10505 31773 10517 31807
rect 10551 31773 10563 31807
rect 10505 31767 10563 31773
rect 4338 31736 4344 31748
rect 3620 31708 4344 31736
rect 4338 31696 4344 31708
rect 4396 31696 4402 31748
rect 4985 31739 5043 31745
rect 4985 31705 4997 31739
rect 5031 31736 5043 31739
rect 5350 31736 5356 31748
rect 5031 31708 5356 31736
rect 5031 31705 5043 31708
rect 4985 31699 5043 31705
rect 5350 31696 5356 31708
rect 5408 31736 5414 31748
rect 6270 31736 6276 31748
rect 5408 31708 6276 31736
rect 5408 31696 5414 31708
rect 6270 31696 6276 31708
rect 6328 31696 6334 31748
rect 7190 31696 7196 31748
rect 7248 31736 7254 31748
rect 7754 31739 7812 31745
rect 7754 31736 7766 31739
rect 7248 31708 7766 31736
rect 7248 31696 7254 31708
rect 7754 31705 7766 31708
rect 7800 31705 7812 31739
rect 10244 31736 10272 31767
rect 10594 31764 10600 31816
rect 10652 31804 10658 31816
rect 10761 31807 10819 31813
rect 10761 31804 10773 31807
rect 10652 31776 10773 31804
rect 10652 31764 10658 31776
rect 10761 31773 10773 31776
rect 10807 31773 10819 31807
rect 10761 31767 10819 31773
rect 36262 31764 36268 31816
rect 36320 31804 36326 31816
rect 36449 31807 36507 31813
rect 36449 31804 36461 31807
rect 36320 31776 36461 31804
rect 36320 31764 36326 31776
rect 36449 31773 36461 31776
rect 36495 31773 36507 31807
rect 38378 31804 38384 31816
rect 37858 31776 38384 31804
rect 36449 31767 36507 31773
rect 38378 31764 38384 31776
rect 38436 31764 38442 31816
rect 39132 31813 39160 31980
rect 39390 31968 39396 31980
rect 39448 31968 39454 32020
rect 39669 32011 39727 32017
rect 39669 31977 39681 32011
rect 39715 32008 39727 32011
rect 40586 32008 40592 32020
rect 39715 31980 40592 32008
rect 39715 31977 39727 31980
rect 39669 31971 39727 31977
rect 40586 31968 40592 31980
rect 40644 31968 40650 32020
rect 42058 31968 42064 32020
rect 42116 31968 42122 32020
rect 42429 32011 42487 32017
rect 42429 31977 42441 32011
rect 42475 32008 42487 32011
rect 43070 32008 43076 32020
rect 42475 31980 43076 32008
rect 42475 31977 42487 31980
rect 42429 31971 42487 31977
rect 43070 31968 43076 31980
rect 43128 31968 43134 32020
rect 44361 32011 44419 32017
rect 43732 31980 44312 32008
rect 43165 31943 43223 31949
rect 43165 31940 43177 31943
rect 42812 31912 43177 31940
rect 39853 31875 39911 31881
rect 39853 31841 39865 31875
rect 39899 31872 39911 31875
rect 40034 31872 40040 31884
rect 39899 31844 40040 31872
rect 39899 31841 39911 31844
rect 39853 31835 39911 31841
rect 40034 31832 40040 31844
rect 40092 31832 40098 31884
rect 41230 31832 41236 31884
rect 41288 31872 41294 31884
rect 41325 31875 41383 31881
rect 41325 31872 41337 31875
rect 41288 31844 41337 31872
rect 41288 31832 41294 31844
rect 41325 31841 41337 31844
rect 41371 31841 41383 31875
rect 41325 31835 41383 31841
rect 41598 31832 41604 31884
rect 41656 31832 41662 31884
rect 42812 31881 42840 31912
rect 43165 31909 43177 31912
rect 43211 31940 43223 31943
rect 43346 31940 43352 31952
rect 43211 31912 43352 31940
rect 43211 31909 43223 31912
rect 43165 31903 43223 31909
rect 43346 31900 43352 31912
rect 43404 31900 43410 31952
rect 42797 31875 42855 31881
rect 42797 31872 42809 31875
rect 42536 31844 42809 31872
rect 39117 31807 39175 31813
rect 38580 31776 39068 31804
rect 10410 31736 10416 31748
rect 10244 31708 10416 31736
rect 7754 31699 7812 31705
rect 10410 31696 10416 31708
rect 10468 31736 10474 31748
rect 13446 31736 13452 31748
rect 10468 31708 13452 31736
rect 10468 31696 10474 31708
rect 13446 31696 13452 31708
rect 13504 31696 13510 31748
rect 36722 31696 36728 31748
rect 36780 31696 36786 31748
rect 38580 31736 38608 31776
rect 38749 31739 38807 31745
rect 38749 31736 38761 31739
rect 38580 31708 38761 31736
rect 38749 31705 38761 31708
rect 38795 31705 38807 31739
rect 39040 31736 39068 31776
rect 39117 31773 39129 31807
rect 39163 31773 39175 31807
rect 39485 31807 39543 31813
rect 39485 31804 39497 31807
rect 39117 31767 39175 31773
rect 39230 31776 39497 31804
rect 39230 31736 39258 31776
rect 39485 31773 39497 31776
rect 39531 31804 39543 31807
rect 39942 31804 39948 31816
rect 39531 31776 39948 31804
rect 39531 31773 39543 31776
rect 39485 31767 39543 31773
rect 39942 31764 39948 31776
rect 40000 31764 40006 31816
rect 42536 31813 42564 31844
rect 42797 31841 42809 31844
rect 42843 31841 42855 31875
rect 42797 31835 42855 31841
rect 42981 31875 43039 31881
rect 42981 31841 42993 31875
rect 43027 31872 43039 31875
rect 43732 31872 43760 31980
rect 44174 31940 44180 31952
rect 43027 31844 43208 31872
rect 43027 31841 43039 31844
rect 42981 31835 43039 31841
rect 42521 31807 42579 31813
rect 42521 31773 42533 31807
rect 42567 31773 42579 31807
rect 42521 31767 42579 31773
rect 43072 31785 43130 31791
rect 43072 31751 43084 31785
rect 43118 31751 43130 31785
rect 39040 31708 39258 31736
rect 39301 31739 39359 31745
rect 38749 31699 38807 31705
rect 39301 31705 39313 31739
rect 39347 31705 39359 31739
rect 39301 31699 39359 31705
rect 3510 31628 3516 31680
rect 3568 31628 3574 31680
rect 4062 31628 4068 31680
rect 4120 31668 4126 31680
rect 10134 31668 10140 31680
rect 4120 31640 10140 31668
rect 4120 31628 4126 31640
rect 10134 31628 10140 31640
rect 10192 31628 10198 31680
rect 11698 31628 11704 31680
rect 11756 31668 11762 31680
rect 11885 31671 11943 31677
rect 11885 31668 11897 31671
rect 11756 31640 11897 31668
rect 11756 31628 11762 31640
rect 11885 31637 11897 31640
rect 11931 31637 11943 31671
rect 11885 31631 11943 31637
rect 38197 31671 38255 31677
rect 38197 31637 38209 31671
rect 38243 31668 38255 31671
rect 38470 31668 38476 31680
rect 38243 31640 38476 31668
rect 38243 31637 38255 31640
rect 38197 31631 38255 31637
rect 38470 31628 38476 31640
rect 38528 31628 38534 31680
rect 38654 31628 38660 31680
rect 38712 31668 38718 31680
rect 39316 31668 39344 31699
rect 39390 31696 39396 31748
rect 39448 31696 39454 31748
rect 41414 31736 41420 31748
rect 40894 31708 41420 31736
rect 41414 31696 41420 31708
rect 41472 31696 41478 31748
rect 43072 31745 43130 31751
rect 43180 31745 43208 31844
rect 43548 31844 43760 31872
rect 44008 31912 44180 31940
rect 43548 31813 43576 31844
rect 43533 31807 43591 31813
rect 43533 31773 43545 31807
rect 43579 31773 43591 31807
rect 43533 31767 43591 31773
rect 43622 31764 43628 31816
rect 43680 31764 43686 31816
rect 44008 31813 44036 31912
rect 44174 31900 44180 31912
rect 44232 31900 44238 31952
rect 44284 31940 44312 31980
rect 44361 31977 44373 32011
rect 44407 32008 44419 32011
rect 44634 32008 44640 32020
rect 44407 31980 44640 32008
rect 44407 31977 44419 31980
rect 44361 31971 44419 31977
rect 44634 31968 44640 31980
rect 44692 31968 44698 32020
rect 45741 32011 45799 32017
rect 45741 31977 45753 32011
rect 45787 32008 45799 32011
rect 46845 32011 46903 32017
rect 46845 32008 46857 32011
rect 45787 31980 46857 32008
rect 45787 31977 45799 31980
rect 45741 31971 45799 31977
rect 46845 31977 46857 31980
rect 46891 31977 46903 32011
rect 46845 31971 46903 31977
rect 47026 31968 47032 32020
rect 47084 31968 47090 32020
rect 47118 31968 47124 32020
rect 47176 31968 47182 32020
rect 48590 31968 48596 32020
rect 48648 32008 48654 32020
rect 50617 32011 50675 32017
rect 48648 31980 49280 32008
rect 48648 31968 48654 31980
rect 44542 31940 44548 31952
rect 44284 31912 44548 31940
rect 44542 31900 44548 31912
rect 44600 31900 44606 31952
rect 45833 31943 45891 31949
rect 45833 31909 45845 31943
rect 45879 31909 45891 31943
rect 45833 31903 45891 31909
rect 46661 31943 46719 31949
rect 46661 31909 46673 31943
rect 46707 31940 46719 31943
rect 47044 31940 47072 31968
rect 46707 31912 47072 31940
rect 47136 31940 47164 31968
rect 47136 31912 47532 31940
rect 46707 31909 46719 31912
rect 46661 31903 46719 31909
rect 43993 31807 44051 31813
rect 43993 31773 44005 31807
rect 44039 31773 44051 31807
rect 43993 31767 44051 31773
rect 44269 31807 44327 31813
rect 44269 31773 44281 31807
rect 44315 31804 44327 31807
rect 44634 31804 44640 31816
rect 44315 31776 44640 31804
rect 44315 31773 44327 31776
rect 44269 31767 44327 31773
rect 38712 31640 39344 31668
rect 42797 31671 42855 31677
rect 38712 31628 38718 31640
rect 42797 31637 42809 31671
rect 42843 31668 42855 31671
rect 42886 31668 42892 31680
rect 42843 31640 42892 31668
rect 42843 31637 42855 31640
rect 42797 31631 42855 31637
rect 42886 31628 42892 31640
rect 42944 31628 42950 31680
rect 43088 31668 43116 31745
rect 43165 31739 43223 31745
rect 43165 31705 43177 31739
rect 43211 31736 43223 31739
rect 44284 31736 44312 31767
rect 44634 31764 44640 31776
rect 44692 31764 44698 31816
rect 45557 31807 45615 31813
rect 45557 31773 45569 31807
rect 45603 31804 45615 31807
rect 45646 31804 45652 31816
rect 45603 31776 45652 31804
rect 45603 31773 45615 31776
rect 45557 31767 45615 31773
rect 45646 31764 45652 31776
rect 45704 31764 45710 31816
rect 45848 31804 45876 31903
rect 45925 31875 45983 31881
rect 45925 31841 45937 31875
rect 45971 31872 45983 31875
rect 47121 31875 47179 31881
rect 47121 31872 47133 31875
rect 45971 31844 47133 31872
rect 45971 31841 45983 31844
rect 45925 31835 45983 31841
rect 47121 31841 47133 31844
rect 47167 31841 47179 31875
rect 47121 31835 47179 31841
rect 46017 31807 46075 31813
rect 46017 31804 46029 31807
rect 45848 31776 46029 31804
rect 46017 31773 46029 31776
rect 46063 31773 46075 31807
rect 46017 31767 46075 31773
rect 46750 31764 46756 31816
rect 46808 31764 46814 31816
rect 47029 31807 47087 31813
rect 47029 31773 47041 31807
rect 47075 31804 47087 31807
rect 47213 31807 47271 31813
rect 47075 31776 47109 31804
rect 47075 31773 47087 31776
rect 47029 31767 47087 31773
rect 47213 31773 47225 31807
rect 47259 31804 47271 31807
rect 47302 31804 47308 31816
rect 47259 31776 47308 31804
rect 47259 31773 47271 31776
rect 47213 31767 47271 31773
rect 43211 31708 44312 31736
rect 43211 31705 43223 31708
rect 43165 31699 43223 31705
rect 44358 31696 44364 31748
rect 44416 31736 44422 31748
rect 45186 31736 45192 31748
rect 44416 31708 45192 31736
rect 44416 31696 44422 31708
rect 45186 31696 45192 31708
rect 45244 31696 45250 31748
rect 47044 31736 47072 31767
rect 47302 31764 47308 31776
rect 47360 31764 47366 31816
rect 47504 31813 47532 31912
rect 48314 31900 48320 31952
rect 48372 31900 48378 31952
rect 49050 31940 49056 31952
rect 48884 31912 49056 31940
rect 47489 31807 47547 31813
rect 47489 31773 47501 31807
rect 47535 31773 47547 31807
rect 48332 31804 48360 31900
rect 48884 31813 48912 31912
rect 49050 31900 49056 31912
rect 49108 31900 49114 31952
rect 48958 31832 48964 31884
rect 49016 31832 49022 31884
rect 49252 31881 49280 31980
rect 50617 31977 50629 32011
rect 50663 32008 50675 32011
rect 51074 32008 51080 32020
rect 50663 31980 51080 32008
rect 50663 31977 50675 31980
rect 50617 31971 50675 31977
rect 51074 31968 51080 31980
rect 51132 31968 51138 32020
rect 53929 32011 53987 32017
rect 53929 31977 53941 32011
rect 53975 32008 53987 32011
rect 54386 32008 54392 32020
rect 53975 31980 54392 32008
rect 53975 31977 53987 31980
rect 53929 31971 53987 31977
rect 54386 31968 54392 31980
rect 54444 31968 54450 32020
rect 55033 32011 55091 32017
rect 55033 31977 55045 32011
rect 55079 32008 55091 32011
rect 55582 32008 55588 32020
rect 55079 31980 55588 32008
rect 55079 31977 55091 31980
rect 55033 31971 55091 31977
rect 55582 31968 55588 31980
rect 55640 31968 55646 32020
rect 50890 31900 50896 31952
rect 50948 31900 50954 31952
rect 52181 31943 52239 31949
rect 52181 31909 52193 31943
rect 52227 31940 52239 31943
rect 52546 31940 52552 31952
rect 52227 31912 52552 31940
rect 52227 31909 52239 31912
rect 52181 31903 52239 31909
rect 52546 31900 52552 31912
rect 52604 31900 52610 31952
rect 54036 31912 55352 31940
rect 49237 31875 49295 31881
rect 49237 31841 49249 31875
rect 49283 31841 49295 31875
rect 49237 31835 49295 31841
rect 49421 31875 49479 31881
rect 49421 31841 49433 31875
rect 49467 31872 49479 31875
rect 49881 31875 49939 31881
rect 49881 31872 49893 31875
rect 49467 31844 49893 31872
rect 49467 31841 49479 31844
rect 49421 31835 49479 31841
rect 49881 31841 49893 31844
rect 49927 31841 49939 31875
rect 49881 31835 49939 31841
rect 48869 31807 48927 31813
rect 48332 31776 48820 31804
rect 47489 31767 47547 31773
rect 47670 31736 47676 31748
rect 47044 31708 47676 31736
rect 47044 31680 47072 31708
rect 47670 31696 47676 31708
rect 47728 31696 47734 31748
rect 48792 31736 48820 31776
rect 48869 31773 48881 31807
rect 48915 31773 48927 31807
rect 49053 31807 49111 31813
rect 49053 31804 49065 31807
rect 48869 31767 48927 31773
rect 48976 31776 49065 31804
rect 48976 31736 49004 31776
rect 49053 31773 49065 31776
rect 49099 31804 49111 31807
rect 49099 31776 49464 31804
rect 49099 31773 49111 31776
rect 49053 31767 49111 31773
rect 48792 31708 49004 31736
rect 49436 31736 49464 31776
rect 49510 31764 49516 31816
rect 49568 31764 49574 31816
rect 49786 31804 49792 31816
rect 49620 31776 49792 31804
rect 49620 31736 49648 31776
rect 49786 31764 49792 31776
rect 49844 31764 49850 31816
rect 49973 31807 50031 31813
rect 49973 31773 49985 31807
rect 50019 31804 50031 31807
rect 50908 31804 50936 31900
rect 52365 31875 52423 31881
rect 52012 31844 52316 31872
rect 50019 31776 50936 31804
rect 50019 31773 50031 31776
rect 49973 31767 50031 31773
rect 51442 31764 51448 31816
rect 51500 31804 51506 31816
rect 52012 31813 52040 31844
rect 51997 31807 52055 31813
rect 51997 31804 52009 31807
rect 51500 31776 52009 31804
rect 51500 31764 51506 31776
rect 51997 31773 52009 31776
rect 52043 31773 52055 31807
rect 51997 31767 52055 31773
rect 52086 31764 52092 31816
rect 52144 31764 52150 31816
rect 52288 31804 52316 31844
rect 52365 31841 52377 31875
rect 52411 31872 52423 31875
rect 52454 31872 52460 31884
rect 52411 31844 52460 31872
rect 52411 31841 52423 31844
rect 52365 31835 52423 31841
rect 52454 31832 52460 31844
rect 52512 31832 52518 31884
rect 52549 31807 52607 31813
rect 52549 31804 52561 31807
rect 52288 31776 52561 31804
rect 52549 31773 52561 31776
rect 52595 31804 52607 31807
rect 54036 31804 54064 31912
rect 55324 31881 55352 31912
rect 55309 31875 55367 31881
rect 55309 31841 55321 31875
rect 55355 31841 55367 31875
rect 55309 31835 55367 31841
rect 54941 31807 54999 31813
rect 54941 31804 54953 31807
rect 52595 31776 54064 31804
rect 54864 31776 54953 31804
rect 52595 31773 52607 31776
rect 52549 31767 52607 31773
rect 49436 31708 49648 31736
rect 51752 31739 51810 31745
rect 48976 31680 49004 31708
rect 51752 31705 51764 31739
rect 51798 31736 51810 31739
rect 52365 31739 52423 31745
rect 52365 31736 52377 31739
rect 51798 31708 52377 31736
rect 51798 31705 51810 31708
rect 51752 31699 51810 31705
rect 52365 31705 52377 31708
rect 52411 31705 52423 31739
rect 52365 31699 52423 31705
rect 52816 31739 52874 31745
rect 52816 31705 52828 31739
rect 52862 31736 52874 31739
rect 53006 31736 53012 31748
rect 52862 31708 53012 31736
rect 52862 31705 52874 31708
rect 52816 31699 52874 31705
rect 53006 31696 53012 31708
rect 53064 31696 53070 31748
rect 54864 31680 54892 31776
rect 54941 31773 54953 31776
rect 54987 31773 54999 31807
rect 54941 31767 54999 31773
rect 55122 31764 55128 31816
rect 55180 31764 55186 31816
rect 55324 31804 55352 31835
rect 56502 31804 56508 31816
rect 55324 31776 56508 31804
rect 56502 31764 56508 31776
rect 56560 31804 56566 31816
rect 56781 31807 56839 31813
rect 56781 31804 56793 31807
rect 56560 31776 56793 31804
rect 56560 31764 56566 31776
rect 56781 31773 56793 31776
rect 56827 31773 56839 31807
rect 56781 31767 56839 31773
rect 58529 31807 58587 31813
rect 58529 31773 58541 31807
rect 58575 31804 58587 31807
rect 58894 31804 58900 31816
rect 58575 31776 58900 31804
rect 58575 31773 58587 31776
rect 58529 31767 58587 31773
rect 58894 31764 58900 31776
rect 58952 31764 58958 31816
rect 55214 31696 55220 31748
rect 55272 31736 55278 31748
rect 55554 31739 55612 31745
rect 55554 31736 55566 31739
rect 55272 31708 55566 31736
rect 55272 31696 55278 31708
rect 55554 31705 55566 31708
rect 55600 31705 55612 31739
rect 55554 31699 55612 31705
rect 56870 31696 56876 31748
rect 56928 31736 56934 31748
rect 57026 31739 57084 31745
rect 57026 31736 57038 31739
rect 56928 31708 57038 31736
rect 56928 31696 56934 31708
rect 57026 31705 57038 31708
rect 57072 31705 57084 31739
rect 57026 31699 57084 31705
rect 46934 31668 46940 31680
rect 43088 31640 46940 31668
rect 46934 31628 46940 31640
rect 46992 31628 46998 31680
rect 47026 31628 47032 31680
rect 47084 31628 47090 31680
rect 47210 31628 47216 31680
rect 47268 31668 47274 31680
rect 47397 31671 47455 31677
rect 47397 31668 47409 31671
rect 47268 31640 47409 31668
rect 47268 31628 47274 31640
rect 47397 31637 47409 31640
rect 47443 31637 47455 31671
rect 47397 31631 47455 31637
rect 48958 31628 48964 31680
rect 49016 31628 49022 31680
rect 49234 31628 49240 31680
rect 49292 31628 49298 31680
rect 54846 31628 54852 31680
rect 54904 31628 54910 31680
rect 56686 31628 56692 31680
rect 56744 31628 56750 31680
rect 58158 31628 58164 31680
rect 58216 31628 58222 31680
rect 58342 31628 58348 31680
rect 58400 31628 58406 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 4890 31424 4896 31476
rect 4948 31424 4954 31476
rect 5626 31424 5632 31476
rect 5684 31464 5690 31476
rect 5997 31467 6055 31473
rect 5997 31464 6009 31467
rect 5684 31436 6009 31464
rect 5684 31424 5690 31436
rect 5997 31433 6009 31436
rect 6043 31433 6055 31467
rect 5997 31427 6055 31433
rect 8386 31424 8392 31476
rect 8444 31464 8450 31476
rect 8481 31467 8539 31473
rect 8481 31464 8493 31467
rect 8444 31436 8493 31464
rect 8444 31424 8450 31436
rect 8481 31433 8493 31436
rect 8527 31433 8539 31467
rect 8481 31427 8539 31433
rect 8588 31436 9674 31464
rect 4982 31396 4988 31408
rect 4080 31368 4988 31396
rect 2682 31288 2688 31340
rect 2740 31288 2746 31340
rect 3878 31288 3884 31340
rect 3936 31288 3942 31340
rect 4080 31337 4108 31368
rect 4982 31356 4988 31368
rect 5040 31356 5046 31408
rect 5077 31399 5135 31405
rect 5077 31365 5089 31399
rect 5123 31396 5135 31399
rect 8588 31396 8616 31436
rect 5123 31368 8616 31396
rect 8849 31399 8907 31405
rect 5123 31365 5135 31368
rect 5077 31359 5135 31365
rect 8849 31365 8861 31399
rect 8895 31396 8907 31399
rect 9030 31396 9036 31408
rect 8895 31368 9036 31396
rect 8895 31365 8907 31368
rect 8849 31359 8907 31365
rect 9030 31356 9036 31368
rect 9088 31356 9094 31408
rect 9646 31396 9674 31436
rect 36722 31424 36728 31476
rect 36780 31464 36786 31476
rect 36909 31467 36967 31473
rect 36909 31464 36921 31467
rect 36780 31436 36921 31464
rect 36780 31424 36786 31436
rect 36909 31433 36921 31436
rect 36955 31433 36967 31467
rect 36909 31427 36967 31433
rect 38289 31467 38347 31473
rect 38289 31433 38301 31467
rect 38335 31464 38347 31467
rect 38654 31464 38660 31476
rect 38335 31436 38660 31464
rect 38335 31433 38347 31436
rect 38289 31427 38347 31433
rect 38654 31424 38660 31436
rect 38712 31424 38718 31476
rect 38838 31424 38844 31476
rect 38896 31464 38902 31476
rect 39117 31467 39175 31473
rect 39117 31464 39129 31467
rect 38896 31436 39129 31464
rect 38896 31424 38902 31436
rect 39117 31433 39129 31436
rect 39163 31433 39175 31467
rect 39117 31427 39175 31433
rect 39482 31424 39488 31476
rect 39540 31464 39546 31476
rect 39577 31467 39635 31473
rect 39577 31464 39589 31467
rect 39540 31436 39589 31464
rect 39540 31424 39546 31436
rect 39577 31433 39589 31436
rect 39623 31433 39635 31467
rect 45554 31464 45560 31476
rect 39577 31427 39635 31433
rect 43456 31436 45560 31464
rect 10042 31396 10048 31408
rect 9646 31368 10048 31396
rect 10042 31356 10048 31368
rect 10100 31356 10106 31408
rect 4065 31331 4123 31337
rect 4065 31297 4077 31331
rect 4111 31297 4123 31331
rect 4065 31291 4123 31297
rect 4154 31288 4160 31340
rect 4212 31288 4218 31340
rect 4338 31288 4344 31340
rect 4396 31328 4402 31340
rect 5166 31328 5172 31340
rect 4396 31300 5172 31328
rect 4396 31288 4402 31300
rect 5166 31288 5172 31300
rect 5224 31288 5230 31340
rect 5261 31331 5319 31337
rect 5261 31297 5273 31331
rect 5307 31328 5319 31331
rect 5997 31331 6055 31337
rect 5997 31328 6009 31331
rect 5307 31300 5672 31328
rect 5307 31297 5319 31300
rect 5261 31291 5319 31297
rect 934 31220 940 31272
rect 992 31260 998 31272
rect 1581 31263 1639 31269
rect 1581 31260 1593 31263
rect 992 31232 1593 31260
rect 992 31220 998 31232
rect 1581 31229 1593 31232
rect 1627 31229 1639 31263
rect 1581 31223 1639 31229
rect 3694 31220 3700 31272
rect 3752 31220 3758 31272
rect 3786 31220 3792 31272
rect 3844 31260 3850 31272
rect 4356 31260 4384 31288
rect 3844 31232 4384 31260
rect 3844 31220 3850 31232
rect 5644 31201 5672 31300
rect 5828 31300 6009 31328
rect 5828 31272 5856 31300
rect 5997 31297 6009 31300
rect 6043 31297 6055 31331
rect 5997 31291 6055 31297
rect 6086 31288 6092 31340
rect 6144 31328 6150 31340
rect 6181 31331 6239 31337
rect 6181 31328 6193 31331
rect 6144 31300 6193 31328
rect 6144 31288 6150 31300
rect 6181 31297 6193 31300
rect 6227 31297 6239 31331
rect 6181 31291 6239 31297
rect 6270 31288 6276 31340
rect 6328 31328 6334 31340
rect 6328 31300 6776 31328
rect 6328 31288 6334 31300
rect 5810 31220 5816 31272
rect 5868 31260 5874 31272
rect 6549 31263 6607 31269
rect 6549 31260 6561 31263
rect 5868 31232 6561 31260
rect 5868 31220 5874 31232
rect 6549 31229 6561 31232
rect 6595 31229 6607 31263
rect 6748 31260 6776 31300
rect 6914 31288 6920 31340
rect 6972 31288 6978 31340
rect 7009 31331 7067 31337
rect 7009 31297 7021 31331
rect 7055 31328 7067 31331
rect 7098 31328 7104 31340
rect 7055 31300 7104 31328
rect 7055 31297 7067 31300
rect 7009 31291 7067 31297
rect 7098 31288 7104 31300
rect 7156 31288 7162 31340
rect 7193 31331 7251 31337
rect 7193 31297 7205 31331
rect 7239 31297 7251 31331
rect 7193 31291 7251 31297
rect 7208 31260 7236 31291
rect 8478 31288 8484 31340
rect 8536 31288 8542 31340
rect 8665 31331 8723 31337
rect 8665 31318 8677 31331
rect 8588 31297 8677 31318
rect 8711 31297 8723 31331
rect 8588 31291 8723 31297
rect 8588 31290 8708 31291
rect 6748 31232 7236 31260
rect 8588 31260 8616 31290
rect 8754 31288 8760 31340
rect 8812 31288 8818 31340
rect 8941 31331 8999 31337
rect 8941 31297 8953 31331
rect 8987 31328 8999 31331
rect 10962 31328 10968 31340
rect 8987 31300 10968 31328
rect 8987 31297 8999 31300
rect 8941 31291 8999 31297
rect 10962 31288 10968 31300
rect 11020 31288 11026 31340
rect 11514 31288 11520 31340
rect 11572 31328 11578 31340
rect 12526 31328 12532 31340
rect 11572 31300 12532 31328
rect 11572 31288 11578 31300
rect 12526 31288 12532 31300
rect 12584 31328 12590 31340
rect 12621 31331 12679 31337
rect 12621 31328 12633 31331
rect 12584 31300 12633 31328
rect 12584 31288 12590 31300
rect 12621 31297 12633 31300
rect 12667 31297 12679 31331
rect 12621 31291 12679 31297
rect 37093 31331 37151 31337
rect 37093 31297 37105 31331
rect 37139 31328 37151 31331
rect 37734 31328 37740 31340
rect 37139 31300 37740 31328
rect 37139 31297 37151 31300
rect 37093 31291 37151 31297
rect 37734 31288 37740 31300
rect 37792 31288 37798 31340
rect 38194 31288 38200 31340
rect 38252 31288 38258 31340
rect 38470 31288 38476 31340
rect 38528 31288 38534 31340
rect 38654 31288 38660 31340
rect 38712 31328 38718 31340
rect 39022 31328 39028 31340
rect 38712 31300 39028 31328
rect 38712 31288 38718 31300
rect 39022 31288 39028 31300
rect 39080 31328 39086 31340
rect 39209 31331 39267 31337
rect 39209 31328 39221 31331
rect 39080 31300 39221 31328
rect 39080 31288 39086 31300
rect 39209 31297 39221 31300
rect 39255 31297 39267 31331
rect 39209 31291 39267 31297
rect 39390 31288 39396 31340
rect 39448 31288 39454 31340
rect 40218 31288 40224 31340
rect 40276 31288 40282 31340
rect 41233 31331 41291 31337
rect 41233 31297 41245 31331
rect 41279 31328 41291 31331
rect 41693 31331 41751 31337
rect 41279 31300 41414 31328
rect 41279 31297 41291 31300
rect 41233 31291 41291 31297
rect 8588 31232 9720 31260
rect 6549 31223 6607 31229
rect 5629 31195 5687 31201
rect 5629 31161 5641 31195
rect 5675 31192 5687 31195
rect 5902 31192 5908 31204
rect 5675 31164 5908 31192
rect 5675 31161 5687 31164
rect 5629 31155 5687 31161
rect 5902 31152 5908 31164
rect 5960 31192 5966 31204
rect 6362 31192 6368 31204
rect 5960 31164 6368 31192
rect 5960 31152 5966 31164
rect 6362 31152 6368 31164
rect 6420 31152 6426 31204
rect 7208 31192 7236 31232
rect 8846 31192 8852 31204
rect 7208 31164 8852 31192
rect 8846 31152 8852 31164
rect 8904 31152 8910 31204
rect 9692 31136 9720 31232
rect 13446 31220 13452 31272
rect 13504 31220 13510 31272
rect 15838 31220 15844 31272
rect 15896 31260 15902 31272
rect 40957 31263 41015 31269
rect 40957 31260 40969 31263
rect 15896 31232 40969 31260
rect 15896 31220 15902 31232
rect 40957 31229 40969 31232
rect 41003 31229 41015 31263
rect 40957 31223 41015 31229
rect 39114 31152 39120 31204
rect 39172 31192 39178 31204
rect 39390 31192 39396 31204
rect 39172 31164 39396 31192
rect 39172 31152 39178 31164
rect 39390 31152 39396 31164
rect 39448 31192 39454 31204
rect 39669 31195 39727 31201
rect 39669 31192 39681 31195
rect 39448 31164 39681 31192
rect 39448 31152 39454 31164
rect 39669 31161 39681 31164
rect 39715 31161 39727 31195
rect 41386 31192 41414 31300
rect 41693 31297 41705 31331
rect 41739 31328 41751 31331
rect 43456 31328 43484 31436
rect 45554 31424 45560 31436
rect 45612 31424 45618 31476
rect 47026 31464 47032 31476
rect 45664 31436 47032 31464
rect 41739 31300 43484 31328
rect 41739 31297 41751 31300
rect 41693 31291 41751 31297
rect 45186 31288 45192 31340
rect 45244 31288 45250 31340
rect 41598 31220 41604 31272
rect 41656 31260 41662 31272
rect 42518 31260 42524 31272
rect 41656 31232 42524 31260
rect 41656 31220 41662 31232
rect 42518 31220 42524 31232
rect 42576 31260 42582 31272
rect 43809 31263 43867 31269
rect 43809 31260 43821 31263
rect 42576 31232 43821 31260
rect 42576 31220 42582 31232
rect 43809 31229 43821 31232
rect 43855 31229 43867 31263
rect 43809 31223 43867 31229
rect 44082 31220 44088 31272
rect 44140 31220 44146 31272
rect 43162 31192 43168 31204
rect 41386 31164 43168 31192
rect 39669 31155 39727 31161
rect 43162 31152 43168 31164
rect 43220 31152 43226 31204
rect 3142 31084 3148 31136
rect 3200 31084 3206 31136
rect 3418 31084 3424 31136
rect 3476 31124 3482 31136
rect 3973 31127 4031 31133
rect 3973 31124 3985 31127
rect 3476 31096 3985 31124
rect 3476 31084 3482 31096
rect 3973 31093 3985 31096
rect 4019 31093 4031 31127
rect 3973 31087 4031 31093
rect 4249 31127 4307 31133
rect 4249 31093 4261 31127
rect 4295 31124 4307 31127
rect 4614 31124 4620 31136
rect 4295 31096 4620 31124
rect 4295 31093 4307 31096
rect 4249 31087 4307 31093
rect 4614 31084 4620 31096
rect 4672 31084 4678 31136
rect 7190 31084 7196 31136
rect 7248 31084 7254 31136
rect 8478 31084 8484 31136
rect 8536 31124 8542 31136
rect 8754 31124 8760 31136
rect 8536 31096 8760 31124
rect 8536 31084 8542 31096
rect 8754 31084 8760 31096
rect 8812 31124 8818 31136
rect 8938 31124 8944 31136
rect 8812 31096 8944 31124
rect 8812 31084 8818 31096
rect 8938 31084 8944 31096
rect 8996 31124 9002 31136
rect 9217 31127 9275 31133
rect 9217 31124 9229 31127
rect 8996 31096 9229 31124
rect 8996 31084 9002 31096
rect 9217 31093 9229 31096
rect 9263 31124 9275 31127
rect 9585 31127 9643 31133
rect 9585 31124 9597 31127
rect 9263 31096 9597 31124
rect 9263 31093 9275 31096
rect 9217 31087 9275 31093
rect 9585 31093 9597 31096
rect 9631 31093 9643 31127
rect 9585 31087 9643 31093
rect 9674 31084 9680 31136
rect 9732 31084 9738 31136
rect 40126 31084 40132 31136
rect 40184 31124 40190 31136
rect 45664 31124 45692 31436
rect 47026 31424 47032 31436
rect 47084 31424 47090 31476
rect 47118 31424 47124 31476
rect 47176 31464 47182 31476
rect 47305 31467 47363 31473
rect 47305 31464 47317 31467
rect 47176 31436 47317 31464
rect 47176 31424 47182 31436
rect 47305 31433 47317 31436
rect 47351 31433 47363 31467
rect 47305 31427 47363 31433
rect 49234 31424 49240 31476
rect 49292 31424 49298 31476
rect 52454 31424 52460 31476
rect 52512 31424 52518 31476
rect 53006 31424 53012 31476
rect 53064 31464 53070 31476
rect 53101 31467 53159 31473
rect 53101 31464 53113 31467
rect 53064 31436 53113 31464
rect 53064 31424 53070 31436
rect 53101 31433 53113 31436
rect 53147 31433 53159 31467
rect 53101 31427 53159 31433
rect 54941 31467 54999 31473
rect 54941 31433 54953 31467
rect 54987 31464 54999 31467
rect 55214 31464 55220 31476
rect 54987 31436 55220 31464
rect 54987 31433 54999 31436
rect 54941 31427 54999 31433
rect 55214 31424 55220 31436
rect 55272 31424 55278 31476
rect 56781 31467 56839 31473
rect 56781 31433 56793 31467
rect 56827 31464 56839 31467
rect 56870 31464 56876 31476
rect 56827 31436 56876 31464
rect 56827 31433 56839 31436
rect 56781 31427 56839 31433
rect 56870 31424 56876 31436
rect 56928 31424 56934 31476
rect 46077 31399 46135 31405
rect 46077 31396 46089 31399
rect 45756 31368 46089 31396
rect 45756 31136 45784 31368
rect 46077 31365 46089 31368
rect 46123 31365 46135 31399
rect 46077 31359 46135 31365
rect 46198 31356 46204 31408
rect 46256 31396 46262 31408
rect 46293 31399 46351 31405
rect 46293 31396 46305 31399
rect 46256 31368 46305 31396
rect 46256 31356 46262 31368
rect 46293 31365 46305 31368
rect 46339 31365 46351 31399
rect 46293 31359 46351 31365
rect 47044 31328 47072 31424
rect 48225 31399 48283 31405
rect 48225 31365 48237 31399
rect 48271 31396 48283 31399
rect 48271 31368 48636 31396
rect 48271 31365 48283 31368
rect 48225 31359 48283 31365
rect 47213 31331 47271 31337
rect 47213 31328 47225 31331
rect 47044 31300 47225 31328
rect 47213 31297 47225 31300
rect 47259 31297 47271 31331
rect 47213 31291 47271 31297
rect 48041 31331 48099 31337
rect 48041 31297 48053 31331
rect 48087 31297 48099 31331
rect 48041 31291 48099 31297
rect 45830 31220 45836 31272
rect 45888 31260 45894 31272
rect 46750 31260 46756 31272
rect 45888 31232 46756 31260
rect 45888 31220 45894 31232
rect 46750 31220 46756 31232
rect 46808 31220 46814 31272
rect 48056 31260 48084 31291
rect 48314 31288 48320 31340
rect 48372 31288 48378 31340
rect 48608 31337 48636 31368
rect 48593 31331 48651 31337
rect 48593 31297 48605 31331
rect 48639 31297 48651 31331
rect 48593 31291 48651 31297
rect 49145 31331 49203 31337
rect 49145 31297 49157 31331
rect 49191 31328 49203 31331
rect 49252 31328 49280 31424
rect 52914 31396 52920 31408
rect 52840 31368 52920 31396
rect 49191 31300 49280 31328
rect 49191 31297 49203 31300
rect 49145 31291 49203 31297
rect 48056 31232 48544 31260
rect 48516 31136 48544 31232
rect 48608 31192 48636 31291
rect 51074 31288 51080 31340
rect 51132 31288 51138 31340
rect 52840 31337 52868 31368
rect 52914 31356 52920 31368
rect 52972 31396 52978 31408
rect 53742 31396 53748 31408
rect 52972 31368 53748 31396
rect 52972 31356 52978 31368
rect 53742 31356 53748 31368
rect 53800 31356 53806 31408
rect 54846 31396 54852 31408
rect 54588 31368 54852 31396
rect 54588 31337 54616 31368
rect 54846 31356 54852 31368
rect 54904 31396 54910 31408
rect 56962 31396 56968 31408
rect 54904 31368 55260 31396
rect 54904 31356 54910 31368
rect 52825 31331 52883 31337
rect 52825 31297 52837 31331
rect 52871 31297 52883 31331
rect 52825 31291 52883 31297
rect 54573 31331 54631 31337
rect 54573 31297 54585 31331
rect 54619 31297 54631 31331
rect 54573 31291 54631 31297
rect 54665 31331 54723 31337
rect 54665 31297 54677 31331
rect 54711 31328 54723 31331
rect 54711 31300 54892 31328
rect 54711 31297 54723 31300
rect 54665 31291 54723 31297
rect 48866 31220 48872 31272
rect 48924 31220 48930 31272
rect 51810 31220 51816 31272
rect 51868 31220 51874 31272
rect 53098 31220 53104 31272
rect 53156 31220 53162 31272
rect 54864 31204 54892 31300
rect 55122 31288 55128 31340
rect 55180 31288 55186 31340
rect 55232 31337 55260 31368
rect 56428 31368 56968 31396
rect 56428 31337 56456 31368
rect 56962 31356 56968 31368
rect 57020 31396 57026 31408
rect 57885 31399 57943 31405
rect 57885 31396 57897 31399
rect 57020 31368 57897 31396
rect 57020 31356 57026 31368
rect 57885 31365 57897 31368
rect 57931 31365 57943 31399
rect 57885 31359 57943 31365
rect 55217 31331 55275 31337
rect 55217 31297 55229 31331
rect 55263 31297 55275 31331
rect 56229 31331 56287 31337
rect 56229 31328 56241 31331
rect 55217 31291 55275 31297
rect 55324 31300 56241 31328
rect 54938 31220 54944 31272
rect 54996 31220 55002 31272
rect 55140 31260 55168 31288
rect 55324 31260 55352 31300
rect 56229 31297 56241 31300
rect 56275 31297 56287 31331
rect 56229 31291 56287 31297
rect 56413 31331 56471 31337
rect 56413 31297 56425 31331
rect 56459 31297 56471 31331
rect 56413 31291 56471 31297
rect 56505 31331 56563 31337
rect 56505 31297 56517 31331
rect 56551 31328 56563 31331
rect 57330 31328 57336 31340
rect 56551 31300 57336 31328
rect 56551 31297 56563 31300
rect 56505 31291 56563 31297
rect 57330 31288 57336 31300
rect 57388 31288 57394 31340
rect 58158 31288 58164 31340
rect 58216 31328 58222 31340
rect 58437 31331 58495 31337
rect 58437 31328 58449 31331
rect 58216 31300 58449 31328
rect 58216 31288 58222 31300
rect 58437 31297 58449 31300
rect 58483 31297 58495 31331
rect 58437 31291 58495 31297
rect 55140 31232 55352 31260
rect 55861 31263 55919 31269
rect 55861 31229 55873 31263
rect 55907 31260 55919 31263
rect 56686 31260 56692 31272
rect 55907 31232 56692 31260
rect 55907 31229 55919 31232
rect 55861 31223 55919 31229
rect 56686 31220 56692 31232
rect 56744 31220 56750 31272
rect 56781 31263 56839 31269
rect 56781 31229 56793 31263
rect 56827 31260 56839 31263
rect 56873 31263 56931 31269
rect 56873 31260 56885 31263
rect 56827 31232 56885 31260
rect 56827 31229 56839 31232
rect 56781 31223 56839 31229
rect 56873 31229 56885 31232
rect 56919 31229 56931 31263
rect 56873 31223 56931 31229
rect 57425 31263 57483 31269
rect 57425 31229 57437 31263
rect 57471 31229 57483 31263
rect 57425 31223 57483 31229
rect 48608 31164 51396 31192
rect 51368 31136 51396 31164
rect 52932 31164 54616 31192
rect 40184 31096 45692 31124
rect 40184 31084 40190 31096
rect 45738 31084 45744 31136
rect 45796 31084 45802 31136
rect 45922 31084 45928 31136
rect 45980 31084 45986 31136
rect 46109 31127 46167 31133
rect 46109 31093 46121 31127
rect 46155 31124 46167 31127
rect 47118 31124 47124 31136
rect 46155 31096 47124 31124
rect 46155 31093 46167 31096
rect 46109 31087 46167 31093
rect 47118 31084 47124 31096
rect 47176 31084 47182 31136
rect 47857 31127 47915 31133
rect 47857 31093 47869 31127
rect 47903 31124 47915 31127
rect 48406 31124 48412 31136
rect 47903 31096 48412 31124
rect 47903 31093 47915 31096
rect 47857 31087 47915 31093
rect 48406 31084 48412 31096
rect 48464 31084 48470 31136
rect 48498 31084 48504 31136
rect 48556 31084 48562 31136
rect 48682 31084 48688 31136
rect 48740 31084 48746 31136
rect 48774 31084 48780 31136
rect 48832 31084 48838 31136
rect 49053 31127 49111 31133
rect 49053 31093 49065 31127
rect 49099 31124 49111 31127
rect 49510 31124 49516 31136
rect 49099 31096 49516 31124
rect 49099 31093 49111 31096
rect 49053 31087 49111 31093
rect 49510 31084 49516 31096
rect 49568 31084 49574 31136
rect 51350 31084 51356 31136
rect 51408 31084 51414 31136
rect 51718 31084 51724 31136
rect 51776 31084 51782 31136
rect 52546 31084 52552 31136
rect 52604 31124 52610 31136
rect 52932 31133 52960 31164
rect 52917 31127 52975 31133
rect 52917 31124 52929 31127
rect 52604 31096 52929 31124
rect 52604 31084 52610 31096
rect 52917 31093 52929 31096
rect 52963 31093 52975 31127
rect 52917 31087 52975 31093
rect 54478 31084 54484 31136
rect 54536 31084 54542 31136
rect 54588 31124 54616 31164
rect 54846 31152 54852 31204
rect 54904 31152 54910 31204
rect 56321 31195 56379 31201
rect 56321 31161 56333 31195
rect 56367 31192 56379 31195
rect 57440 31192 57468 31223
rect 56367 31164 57468 31192
rect 56367 31161 56379 31164
rect 56321 31155 56379 31161
rect 54757 31127 54815 31133
rect 54757 31124 54769 31127
rect 54588 31096 54769 31124
rect 54757 31093 54769 31096
rect 54803 31124 54815 31127
rect 56134 31124 56140 31136
rect 54803 31096 56140 31124
rect 54803 31093 54815 31096
rect 54757 31087 54815 31093
rect 56134 31084 56140 31096
rect 56192 31124 56198 31136
rect 56597 31127 56655 31133
rect 56597 31124 56609 31127
rect 56192 31096 56609 31124
rect 56192 31084 56198 31096
rect 56597 31093 56609 31096
rect 56643 31093 56655 31127
rect 56597 31087 56655 31093
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 3142 30920 3148 30932
rect 3068 30892 3148 30920
rect 2869 30787 2927 30793
rect 2869 30753 2881 30787
rect 2915 30784 2927 30787
rect 3068 30784 3096 30892
rect 3142 30880 3148 30892
rect 3200 30880 3206 30932
rect 3421 30923 3479 30929
rect 3421 30889 3433 30923
rect 3467 30920 3479 30923
rect 3694 30920 3700 30932
rect 3467 30892 3700 30920
rect 3467 30889 3479 30892
rect 3421 30883 3479 30889
rect 3694 30880 3700 30892
rect 3752 30880 3758 30932
rect 7006 30880 7012 30932
rect 7064 30920 7070 30932
rect 7101 30923 7159 30929
rect 7101 30920 7113 30923
rect 7064 30892 7113 30920
rect 7064 30880 7070 30892
rect 7101 30889 7113 30892
rect 7147 30889 7159 30923
rect 7101 30883 7159 30889
rect 8294 30880 8300 30932
rect 8352 30920 8358 30932
rect 9033 30923 9091 30929
rect 9033 30920 9045 30923
rect 8352 30892 9045 30920
rect 8352 30880 8358 30892
rect 9033 30889 9045 30892
rect 9079 30889 9091 30923
rect 9033 30883 9091 30889
rect 9214 30880 9220 30932
rect 9272 30920 9278 30932
rect 9309 30923 9367 30929
rect 9309 30920 9321 30923
rect 9272 30892 9321 30920
rect 9272 30880 9278 30892
rect 9309 30889 9321 30892
rect 9355 30889 9367 30923
rect 9309 30883 9367 30889
rect 10134 30880 10140 30932
rect 10192 30920 10198 30932
rect 10689 30923 10747 30929
rect 10689 30920 10701 30923
rect 10192 30892 10701 30920
rect 10192 30880 10198 30892
rect 10689 30889 10701 30892
rect 10735 30889 10747 30923
rect 10689 30883 10747 30889
rect 38105 30923 38163 30929
rect 38105 30889 38117 30923
rect 38151 30920 38163 30923
rect 38194 30920 38200 30932
rect 38151 30892 38200 30920
rect 38151 30889 38163 30892
rect 38105 30883 38163 30889
rect 38194 30880 38200 30892
rect 38252 30880 38258 30932
rect 38654 30880 38660 30932
rect 38712 30880 38718 30932
rect 39942 30880 39948 30932
rect 40000 30880 40006 30932
rect 44082 30880 44088 30932
rect 44140 30920 44146 30932
rect 44637 30923 44695 30929
rect 44637 30920 44649 30923
rect 44140 30892 44649 30920
rect 44140 30880 44146 30892
rect 44637 30889 44649 30892
rect 44683 30889 44695 30923
rect 45922 30920 45928 30932
rect 44637 30883 44695 30889
rect 44928 30892 45928 30920
rect 3160 30824 8248 30852
rect 3160 30796 3188 30824
rect 8220 30796 8248 30824
rect 9674 30812 9680 30864
rect 9732 30852 9738 30864
rect 11698 30852 11704 30864
rect 9732 30824 11704 30852
rect 9732 30812 9738 30824
rect 11698 30812 11704 30824
rect 11756 30812 11762 30864
rect 39960 30852 39988 30880
rect 38488 30824 39988 30852
rect 42245 30855 42303 30861
rect 2915 30756 3096 30784
rect 2915 30753 2927 30756
rect 2869 30747 2927 30753
rect 3142 30744 3148 30796
rect 3200 30744 3206 30796
rect 3418 30784 3424 30796
rect 3252 30756 3424 30784
rect 3252 30725 3280 30756
rect 3418 30744 3424 30756
rect 3476 30744 3482 30796
rect 3513 30787 3571 30793
rect 3513 30753 3525 30787
rect 3559 30784 3571 30787
rect 3789 30787 3847 30793
rect 3789 30784 3801 30787
rect 3559 30756 3801 30784
rect 3559 30753 3571 30756
rect 3513 30747 3571 30753
rect 3789 30753 3801 30756
rect 3835 30753 3847 30787
rect 3789 30747 3847 30753
rect 4433 30787 4491 30793
rect 4433 30753 4445 30787
rect 4479 30784 4491 30787
rect 4614 30784 4620 30796
rect 4479 30756 4620 30784
rect 4479 30753 4491 30756
rect 4433 30747 4491 30753
rect 4614 30744 4620 30756
rect 4672 30744 4678 30796
rect 8202 30744 8208 30796
rect 8260 30744 8266 30796
rect 9140 30756 9628 30784
rect 3237 30719 3295 30725
rect 3237 30685 3249 30719
rect 3283 30685 3295 30719
rect 3237 30679 3295 30685
rect 3326 30676 3332 30728
rect 3384 30676 3390 30728
rect 3878 30676 3884 30728
rect 3936 30676 3942 30728
rect 4525 30719 4583 30725
rect 4525 30685 4537 30719
rect 4571 30716 4583 30719
rect 5810 30716 5816 30728
rect 4571 30688 5816 30716
rect 4571 30685 4583 30688
rect 4525 30679 4583 30685
rect 2406 30608 2412 30660
rect 2464 30608 2470 30660
rect 3896 30648 3924 30676
rect 4801 30651 4859 30657
rect 4801 30648 4813 30651
rect 3896 30620 4813 30648
rect 4801 30617 4813 30620
rect 4847 30648 4859 30651
rect 5074 30648 5080 30660
rect 4847 30620 5080 30648
rect 4847 30617 4859 30620
rect 4801 30611 4859 30617
rect 5074 30608 5080 30620
rect 5132 30608 5138 30660
rect 1397 30583 1455 30589
rect 1397 30549 1409 30583
rect 1443 30580 1455 30583
rect 2682 30580 2688 30592
rect 1443 30552 2688 30580
rect 1443 30549 1455 30552
rect 1397 30543 1455 30549
rect 2682 30540 2688 30552
rect 2740 30540 2746 30592
rect 5368 30589 5396 30688
rect 5810 30676 5816 30688
rect 5868 30676 5874 30728
rect 6089 30719 6147 30725
rect 6089 30685 6101 30719
rect 6135 30716 6147 30719
rect 6362 30716 6368 30728
rect 6135 30688 6368 30716
rect 6135 30685 6147 30688
rect 6089 30679 6147 30685
rect 6362 30676 6368 30688
rect 6420 30676 6426 30728
rect 7009 30719 7067 30725
rect 7009 30685 7021 30719
rect 7055 30685 7067 30719
rect 7009 30679 7067 30685
rect 7193 30719 7251 30725
rect 7193 30685 7205 30719
rect 7239 30716 7251 30719
rect 7466 30716 7472 30728
rect 7239 30688 7472 30716
rect 7239 30685 7251 30688
rect 7193 30679 7251 30685
rect 5828 30648 5856 30676
rect 7024 30648 7052 30679
rect 7466 30676 7472 30688
rect 7524 30676 7530 30728
rect 8938 30676 8944 30728
rect 8996 30676 9002 30728
rect 9140 30725 9168 30756
rect 9125 30719 9183 30725
rect 9125 30685 9137 30719
rect 9171 30685 9183 30719
rect 9125 30679 9183 30685
rect 9217 30719 9275 30725
rect 9217 30685 9229 30719
rect 9263 30685 9275 30719
rect 9401 30719 9459 30725
rect 9401 30716 9413 30719
rect 9217 30679 9275 30685
rect 9324 30688 9413 30716
rect 7561 30651 7619 30657
rect 7561 30648 7573 30651
rect 5828 30620 7573 30648
rect 7561 30617 7573 30620
rect 7607 30648 7619 30651
rect 8665 30651 8723 30657
rect 8665 30648 8677 30651
rect 7607 30620 8677 30648
rect 7607 30617 7619 30620
rect 7561 30611 7619 30617
rect 8665 30617 8677 30620
rect 8711 30648 8723 30651
rect 8956 30648 8984 30676
rect 9232 30648 9260 30679
rect 8711 30620 9260 30648
rect 8711 30617 8723 30620
rect 8665 30611 8723 30617
rect 9324 30592 9352 30688
rect 9401 30685 9413 30688
rect 9447 30685 9459 30719
rect 9401 30679 9459 30685
rect 9600 30648 9628 30756
rect 9692 30725 9720 30812
rect 38488 30725 38516 30824
rect 42245 30821 42257 30855
rect 42291 30821 42303 30855
rect 42245 30815 42303 30821
rect 39574 30744 39580 30796
rect 39632 30784 39638 30796
rect 39853 30787 39911 30793
rect 39853 30784 39865 30787
rect 39632 30756 39865 30784
rect 39632 30744 39638 30756
rect 39853 30753 39865 30756
rect 39899 30753 39911 30787
rect 39853 30747 39911 30753
rect 41322 30744 41328 30796
rect 41380 30744 41386 30796
rect 41966 30744 41972 30796
rect 42024 30784 42030 30796
rect 42024 30756 42104 30784
rect 42024 30744 42030 30756
rect 9677 30719 9735 30725
rect 9677 30685 9689 30719
rect 9723 30685 9735 30719
rect 9677 30679 9735 30685
rect 9861 30719 9919 30725
rect 9861 30685 9873 30719
rect 9907 30716 9919 30719
rect 9953 30719 10011 30725
rect 9953 30716 9965 30719
rect 9907 30688 9965 30716
rect 9907 30685 9919 30688
rect 9861 30679 9919 30685
rect 9953 30685 9965 30688
rect 9999 30685 10011 30719
rect 9953 30679 10011 30685
rect 38473 30719 38531 30725
rect 38473 30685 38485 30719
rect 38519 30685 38531 30719
rect 38473 30679 38531 30685
rect 38749 30719 38807 30725
rect 38749 30685 38761 30719
rect 38795 30716 38807 30719
rect 38838 30716 38844 30728
rect 38795 30688 38844 30716
rect 38795 30685 38807 30688
rect 38749 30679 38807 30685
rect 9766 30648 9772 30660
rect 9600 30620 9772 30648
rect 9766 30608 9772 30620
rect 9824 30608 9830 30660
rect 9968 30592 9996 30679
rect 38838 30676 38844 30688
rect 38896 30676 38902 30728
rect 40034 30676 40040 30728
rect 40092 30676 40098 30728
rect 40126 30676 40132 30728
rect 40184 30676 40190 30728
rect 42076 30725 42104 30756
rect 42061 30719 42119 30725
rect 42061 30685 42073 30719
rect 42107 30685 42119 30719
rect 42260 30716 42288 30815
rect 43809 30787 43867 30793
rect 43809 30753 43821 30787
rect 43855 30784 43867 30787
rect 43993 30787 44051 30793
rect 43993 30784 44005 30787
rect 43855 30756 44005 30784
rect 43855 30753 43867 30756
rect 43809 30747 43867 30753
rect 43993 30753 44005 30756
rect 44039 30753 44051 30787
rect 43993 30747 44051 30753
rect 42978 30716 42984 30728
rect 42260 30688 42984 30716
rect 42061 30679 42119 30685
rect 42978 30676 42984 30688
rect 43036 30676 43042 30728
rect 43162 30676 43168 30728
rect 43220 30676 43226 30728
rect 43714 30676 43720 30728
rect 43772 30676 43778 30728
rect 43901 30719 43959 30725
rect 43901 30685 43913 30719
rect 43947 30716 43959 30719
rect 44928 30716 44956 30892
rect 45922 30880 45928 30892
rect 45980 30880 45986 30932
rect 48498 30880 48504 30932
rect 48556 30880 48562 30932
rect 48774 30880 48780 30932
rect 48832 30920 48838 30932
rect 51445 30923 51503 30929
rect 48832 30892 49280 30920
rect 48832 30880 48838 30892
rect 45738 30812 45744 30864
rect 45796 30812 45802 30864
rect 45830 30784 45836 30796
rect 43947 30688 44956 30716
rect 45388 30756 45836 30784
rect 45388 30716 45416 30756
rect 45830 30744 45836 30756
rect 45888 30744 45894 30796
rect 47394 30784 47400 30796
rect 46676 30756 47400 30784
rect 45465 30719 45523 30725
rect 45465 30716 45477 30719
rect 45388 30688 45477 30716
rect 43947 30685 43959 30688
rect 43901 30679 43959 30685
rect 45465 30685 45477 30688
rect 45511 30685 45523 30719
rect 45465 30679 45523 30685
rect 10042 30608 10048 30660
rect 10100 30648 10106 30660
rect 10137 30651 10195 30657
rect 10137 30648 10149 30651
rect 10100 30620 10149 30648
rect 10100 30608 10106 30620
rect 10137 30617 10149 30620
rect 10183 30617 10195 30651
rect 10137 30611 10195 30617
rect 12161 30651 12219 30657
rect 12161 30617 12173 30651
rect 12207 30648 12219 30651
rect 12529 30651 12587 30657
rect 12529 30648 12541 30651
rect 12207 30620 12541 30648
rect 12207 30617 12219 30620
rect 12161 30611 12219 30617
rect 12529 30617 12541 30620
rect 12575 30648 12587 30651
rect 13722 30648 13728 30660
rect 12575 30620 13728 30648
rect 12575 30617 12587 30620
rect 12529 30611 12587 30617
rect 13722 30608 13728 30620
rect 13780 30648 13786 30660
rect 15657 30651 15715 30657
rect 15657 30648 15669 30651
rect 13780 30620 15669 30648
rect 13780 30608 13786 30620
rect 15657 30617 15669 30620
rect 15703 30617 15715 30651
rect 15657 30611 15715 30617
rect 5353 30583 5411 30589
rect 5353 30549 5365 30583
rect 5399 30580 5411 30583
rect 5442 30580 5448 30592
rect 5399 30552 5448 30580
rect 5399 30549 5411 30552
rect 5353 30543 5411 30549
rect 5442 30540 5448 30552
rect 5500 30540 5506 30592
rect 6178 30540 6184 30592
rect 6236 30540 6242 30592
rect 6362 30540 6368 30592
rect 6420 30580 6426 30592
rect 6549 30583 6607 30589
rect 6549 30580 6561 30583
rect 6420 30552 6561 30580
rect 6420 30540 6426 30552
rect 6549 30549 6561 30552
rect 6595 30580 6607 30583
rect 6730 30580 6736 30592
rect 6595 30552 6736 30580
rect 6595 30549 6607 30552
rect 6549 30543 6607 30549
rect 6730 30540 6736 30552
rect 6788 30540 6794 30592
rect 9306 30540 9312 30592
rect 9364 30540 9370 30592
rect 9858 30540 9864 30592
rect 9916 30540 9922 30592
rect 9950 30540 9956 30592
rect 10008 30540 10014 30592
rect 10318 30540 10324 30592
rect 10376 30540 10382 30592
rect 10594 30540 10600 30592
rect 10652 30580 10658 30592
rect 12894 30580 12900 30592
rect 10652 30552 12900 30580
rect 10652 30540 10658 30552
rect 12894 30540 12900 30552
rect 12952 30540 12958 30592
rect 15672 30580 15700 30611
rect 17126 30608 17132 30660
rect 17184 30648 17190 30660
rect 17405 30651 17463 30657
rect 17405 30648 17417 30651
rect 17184 30620 17417 30648
rect 17184 30608 17190 30620
rect 17405 30617 17417 30620
rect 17451 30648 17463 30651
rect 17451 30620 22094 30648
rect 17451 30617 17463 30620
rect 17405 30611 17463 30617
rect 17681 30583 17739 30589
rect 17681 30580 17693 30583
rect 15672 30552 17693 30580
rect 17681 30549 17693 30552
rect 17727 30549 17739 30583
rect 22066 30580 22094 30620
rect 38286 30608 38292 30660
rect 38344 30608 38350 30660
rect 41969 30651 42027 30657
rect 41969 30617 41981 30651
rect 42015 30648 42027 30651
rect 42794 30648 42800 30660
rect 42015 30620 42800 30648
rect 42015 30617 42027 30620
rect 41969 30611 42027 30617
rect 42794 30608 42800 30620
rect 42852 30608 42858 30660
rect 43180 30648 43208 30676
rect 45480 30648 45508 30679
rect 45554 30676 45560 30728
rect 45612 30676 45618 30728
rect 45646 30676 45652 30728
rect 45704 30716 45710 30728
rect 46676 30725 46704 30756
rect 47394 30744 47400 30756
rect 47452 30744 47458 30796
rect 49252 30793 49280 30892
rect 51445 30889 51457 30923
rect 51491 30920 51503 30923
rect 51810 30920 51816 30932
rect 51491 30892 51816 30920
rect 51491 30889 51503 30892
rect 51445 30883 51503 30889
rect 51810 30880 51816 30892
rect 51868 30880 51874 30932
rect 54478 30880 54484 30932
rect 54536 30880 54542 30932
rect 56962 30880 56968 30932
rect 57020 30880 57026 30932
rect 57330 30880 57336 30932
rect 57388 30880 57394 30932
rect 48409 30787 48467 30793
rect 48409 30753 48421 30787
rect 48455 30784 48467 30787
rect 49053 30787 49111 30793
rect 49053 30784 49065 30787
rect 48455 30756 49065 30784
rect 48455 30753 48467 30756
rect 48409 30747 48467 30753
rect 49053 30753 49065 30756
rect 49099 30753 49111 30787
rect 49053 30747 49111 30753
rect 49237 30787 49295 30793
rect 49237 30753 49249 30787
rect 49283 30753 49295 30787
rect 51718 30784 51724 30796
rect 49237 30747 49295 30753
rect 51368 30756 51724 30784
rect 51368 30725 51396 30756
rect 51718 30744 51724 30756
rect 51776 30744 51782 30796
rect 54496 30784 54524 30880
rect 53024 30756 53328 30784
rect 46661 30719 46719 30725
rect 46661 30716 46673 30719
rect 45704 30688 46673 30716
rect 45704 30676 45710 30688
rect 46661 30685 46673 30688
rect 46707 30685 46719 30719
rect 46661 30679 46719 30685
rect 51353 30719 51411 30725
rect 51353 30685 51365 30719
rect 51399 30685 51411 30719
rect 51537 30719 51595 30725
rect 51537 30716 51549 30719
rect 51353 30679 51411 30685
rect 51442 30688 51549 30716
rect 43180 30620 45508 30648
rect 36262 30580 36268 30592
rect 22066 30552 36268 30580
rect 17681 30543 17739 30549
rect 36262 30540 36268 30552
rect 36320 30540 36326 30592
rect 43070 30540 43076 30592
rect 43128 30540 43134 30592
rect 45572 30580 45600 30676
rect 45738 30608 45744 30660
rect 45796 30608 45802 30660
rect 46937 30651 46995 30657
rect 46937 30617 46949 30651
rect 46983 30648 46995 30651
rect 47210 30648 47216 30660
rect 46983 30620 47216 30648
rect 46983 30617 46995 30620
rect 46937 30611 46995 30617
rect 47210 30608 47216 30620
rect 47268 30608 47274 30660
rect 47320 30620 47426 30648
rect 47320 30592 47348 30620
rect 51166 30608 51172 30660
rect 51224 30648 51230 30660
rect 51442 30648 51470 30688
rect 51537 30685 51549 30688
rect 51583 30685 51595 30719
rect 53024 30716 53052 30756
rect 51537 30679 51595 30685
rect 51644 30688 53052 30716
rect 51224 30620 51470 30648
rect 51224 30608 51230 30620
rect 51644 30592 51672 30688
rect 53098 30676 53104 30728
rect 53156 30676 53162 30728
rect 53300 30725 53328 30756
rect 54312 30756 54524 30784
rect 54312 30725 54340 30756
rect 56980 30725 57008 30880
rect 57348 30852 57376 30880
rect 58253 30855 58311 30861
rect 58253 30852 58265 30855
rect 57348 30824 58265 30852
rect 57241 30787 57299 30793
rect 57241 30753 57253 30787
rect 57287 30784 57299 30787
rect 57425 30787 57483 30793
rect 57425 30784 57437 30787
rect 57287 30756 57437 30784
rect 57287 30753 57299 30756
rect 57241 30747 57299 30753
rect 57425 30753 57437 30756
rect 57471 30753 57483 30787
rect 57425 30747 57483 30753
rect 57532 30725 57560 30824
rect 58253 30821 58265 30824
rect 58299 30821 58311 30855
rect 58253 30815 58311 30821
rect 58618 30784 58624 30796
rect 57900 30756 58624 30784
rect 57900 30725 57928 30756
rect 58618 30744 58624 30756
rect 58676 30744 58682 30796
rect 53193 30719 53251 30725
rect 53193 30685 53205 30719
rect 53239 30685 53251 30719
rect 53193 30679 53251 30685
rect 53285 30719 53343 30725
rect 53285 30685 53297 30719
rect 53331 30716 53343 30719
rect 54297 30719 54355 30725
rect 53331 30688 54248 30716
rect 53331 30685 53343 30688
rect 53285 30679 53343 30685
rect 51810 30608 51816 30660
rect 51868 30648 51874 30660
rect 53208 30648 53236 30679
rect 54113 30651 54171 30657
rect 54113 30648 54125 30651
rect 51868 30620 54125 30648
rect 51868 30608 51874 30620
rect 54113 30617 54125 30620
rect 54159 30617 54171 30651
rect 54220 30648 54248 30688
rect 54297 30685 54309 30719
rect 54343 30685 54355 30719
rect 54297 30679 54355 30685
rect 54389 30719 54447 30725
rect 54389 30685 54401 30719
rect 54435 30685 54447 30719
rect 54389 30679 54447 30685
rect 56965 30719 57023 30725
rect 56965 30685 56977 30719
rect 57011 30685 57023 30719
rect 56965 30679 57023 30685
rect 57057 30719 57115 30725
rect 57057 30685 57069 30719
rect 57103 30716 57115 30719
rect 57333 30719 57391 30725
rect 57333 30716 57345 30719
rect 57103 30688 57345 30716
rect 57103 30685 57115 30688
rect 57057 30679 57115 30685
rect 57333 30685 57345 30688
rect 57379 30685 57391 30719
rect 57333 30679 57391 30685
rect 57517 30719 57575 30725
rect 57517 30685 57529 30719
rect 57563 30685 57575 30719
rect 57517 30679 57575 30685
rect 57885 30719 57943 30725
rect 57885 30685 57897 30719
rect 57931 30685 57943 30719
rect 57885 30679 57943 30685
rect 54404 30648 54432 30679
rect 54220 30620 54432 30648
rect 57348 30648 57376 30679
rect 58342 30676 58348 30728
rect 58400 30676 58406 30728
rect 57348 30620 57652 30648
rect 54113 30611 54171 30617
rect 57624 30592 57652 30620
rect 46017 30583 46075 30589
rect 46017 30580 46029 30583
rect 45572 30552 46029 30580
rect 46017 30549 46029 30552
rect 46063 30549 46075 30583
rect 46017 30543 46075 30549
rect 46658 30540 46664 30592
rect 46716 30580 46722 30592
rect 47302 30580 47308 30592
rect 46716 30552 47308 30580
rect 46716 30540 46722 30552
rect 47302 30540 47308 30552
rect 47360 30540 47366 30592
rect 49881 30583 49939 30589
rect 49881 30549 49893 30583
rect 49927 30580 49939 30583
rect 50154 30580 50160 30592
rect 49927 30552 50160 30580
rect 49927 30549 49939 30552
rect 49881 30543 49939 30549
rect 50154 30540 50160 30552
rect 50212 30540 50218 30592
rect 51626 30540 51632 30592
rect 51684 30540 51690 30592
rect 53466 30540 53472 30592
rect 53524 30540 53530 30592
rect 54294 30540 54300 30592
rect 54352 30540 54358 30592
rect 57238 30540 57244 30592
rect 57296 30540 57302 30592
rect 57606 30540 57612 30592
rect 57664 30540 57670 30592
rect 58066 30540 58072 30592
rect 58124 30540 58130 30592
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 3329 30379 3387 30385
rect 3329 30345 3341 30379
rect 3375 30376 3387 30379
rect 4062 30376 4068 30388
rect 3375 30348 4068 30376
rect 3375 30345 3387 30348
rect 3329 30339 3387 30345
rect 4062 30336 4068 30348
rect 4120 30336 4126 30388
rect 5451 30379 5509 30385
rect 5451 30345 5463 30379
rect 5497 30345 5509 30379
rect 5451 30339 5509 30345
rect 2593 30311 2651 30317
rect 2593 30277 2605 30311
rect 2639 30308 2651 30311
rect 3142 30308 3148 30320
rect 2639 30280 3148 30308
rect 2639 30277 2651 30280
rect 2593 30271 2651 30277
rect 3142 30268 3148 30280
rect 3200 30268 3206 30320
rect 5016 30311 5074 30317
rect 5016 30277 5028 30311
rect 5062 30308 5074 30311
rect 5460 30308 5488 30339
rect 5902 30336 5908 30388
rect 5960 30336 5966 30388
rect 9858 30336 9864 30388
rect 9916 30336 9922 30388
rect 10229 30379 10287 30385
rect 10229 30345 10241 30379
rect 10275 30376 10287 30379
rect 10318 30376 10324 30388
rect 10275 30348 10324 30376
rect 10275 30345 10287 30348
rect 10229 30339 10287 30345
rect 10318 30336 10324 30348
rect 10376 30376 10382 30388
rect 10689 30379 10747 30385
rect 10689 30376 10701 30379
rect 10376 30348 10701 30376
rect 10376 30336 10382 30348
rect 10689 30345 10701 30348
rect 10735 30345 10747 30379
rect 11054 30376 11060 30388
rect 10689 30339 10747 30345
rect 10796 30348 11060 30376
rect 5813 30311 5871 30317
rect 5813 30308 5825 30311
rect 5062 30280 5488 30308
rect 5644 30280 5825 30308
rect 5062 30277 5074 30280
rect 5016 30271 5074 30277
rect 2682 30200 2688 30252
rect 2740 30200 2746 30252
rect 3421 30243 3479 30249
rect 3421 30209 3433 30243
rect 3467 30240 3479 30243
rect 4062 30240 4068 30252
rect 3467 30212 4068 30240
rect 3467 30209 3479 30212
rect 3421 30203 3479 30209
rect 4062 30200 4068 30212
rect 4120 30200 4126 30252
rect 5166 30240 5172 30252
rect 4264 30212 5172 30240
rect 3694 30132 3700 30184
rect 3752 30132 3758 30184
rect 3326 30064 3332 30116
rect 3384 30104 3390 30116
rect 3513 30107 3571 30113
rect 3513 30104 3525 30107
rect 3384 30076 3525 30104
rect 3384 30064 3390 30076
rect 3513 30073 3525 30076
rect 3559 30104 3571 30107
rect 4264 30104 4292 30212
rect 5166 30200 5172 30212
rect 5224 30200 5230 30252
rect 5350 30200 5356 30252
rect 5408 30200 5414 30252
rect 5534 30200 5540 30252
rect 5592 30200 5598 30252
rect 5644 30249 5672 30280
rect 5813 30277 5825 30280
rect 5859 30277 5871 30311
rect 5813 30271 5871 30277
rect 5920 30249 5948 30336
rect 6822 30268 6828 30320
rect 6880 30268 6886 30320
rect 5629 30243 5687 30249
rect 5629 30209 5641 30243
rect 5675 30209 5687 30243
rect 5629 30203 5687 30209
rect 5721 30243 5779 30249
rect 5721 30209 5733 30243
rect 5767 30209 5779 30243
rect 5721 30203 5779 30209
rect 5905 30243 5963 30249
rect 5905 30209 5917 30243
rect 5951 30209 5963 30243
rect 5905 30203 5963 30209
rect 5261 30175 5319 30181
rect 5261 30141 5273 30175
rect 5307 30141 5319 30175
rect 5261 30135 5319 30141
rect 3559 30076 4292 30104
rect 5276 30104 5304 30135
rect 5626 30104 5632 30116
rect 5276 30076 5632 30104
rect 3559 30073 3571 30076
rect 3513 30067 3571 30073
rect 5626 30064 5632 30076
rect 5684 30064 5690 30116
rect 3602 29996 3608 30048
rect 3660 29996 3666 30048
rect 3881 30039 3939 30045
rect 3881 30005 3893 30039
rect 3927 30036 3939 30039
rect 4890 30036 4896 30048
rect 3927 30008 4896 30036
rect 3927 30005 3939 30008
rect 3881 29999 3939 30005
rect 4890 29996 4896 30008
rect 4948 30036 4954 30048
rect 5736 30036 5764 30203
rect 6178 30200 6184 30252
rect 6236 30240 6242 30252
rect 6638 30249 6644 30252
rect 6365 30243 6423 30249
rect 6365 30240 6377 30243
rect 6236 30212 6377 30240
rect 6236 30200 6242 30212
rect 6365 30209 6377 30212
rect 6411 30209 6423 30243
rect 6632 30240 6644 30249
rect 6599 30212 6644 30240
rect 6365 30203 6423 30209
rect 6632 30203 6644 30212
rect 6638 30200 6644 30203
rect 6696 30200 6702 30252
rect 6840 30240 6868 30268
rect 9876 30240 9904 30336
rect 10413 30311 10471 30317
rect 10413 30277 10425 30311
rect 10459 30308 10471 30311
rect 10594 30308 10600 30320
rect 10459 30280 10600 30308
rect 10459 30277 10471 30280
rect 10413 30271 10471 30277
rect 10137 30243 10195 30249
rect 10137 30240 10149 30243
rect 6840 30212 9674 30240
rect 9876 30212 10149 30240
rect 9646 30172 9674 30212
rect 10137 30209 10149 30212
rect 10183 30209 10195 30243
rect 10137 30203 10195 30209
rect 10428 30172 10456 30271
rect 10594 30268 10600 30280
rect 10652 30268 10658 30320
rect 10502 30243 10560 30249
rect 10502 30209 10514 30243
rect 10548 30240 10560 30243
rect 10686 30240 10692 30252
rect 10548 30212 10692 30240
rect 10548 30209 10560 30212
rect 10502 30203 10560 30209
rect 10686 30200 10692 30212
rect 10744 30200 10750 30252
rect 10796 30249 10824 30348
rect 11054 30336 11060 30348
rect 11112 30336 11118 30388
rect 12897 30379 12955 30385
rect 12897 30345 12909 30379
rect 12943 30345 12955 30379
rect 12897 30339 12955 30345
rect 39945 30379 40003 30385
rect 39945 30345 39957 30379
rect 39991 30376 40003 30379
rect 40034 30376 40040 30388
rect 39991 30348 40040 30376
rect 39991 30345 40003 30348
rect 39945 30339 40003 30345
rect 10962 30268 10968 30320
rect 11020 30308 11026 30320
rect 12618 30308 12624 30320
rect 11020 30280 12624 30308
rect 11020 30268 11026 30280
rect 12618 30268 12624 30280
rect 12676 30308 12682 30320
rect 12912 30308 12940 30339
rect 39960 30308 39988 30339
rect 40034 30336 40040 30348
rect 40092 30336 40098 30388
rect 43070 30336 43076 30388
rect 43128 30336 43134 30388
rect 43714 30336 43720 30388
rect 43772 30336 43778 30388
rect 45738 30336 45744 30388
rect 45796 30376 45802 30388
rect 46477 30379 46535 30385
rect 46477 30376 46489 30379
rect 45796 30348 46489 30376
rect 45796 30336 45802 30348
rect 46477 30345 46489 30348
rect 46523 30376 46535 30379
rect 46566 30376 46572 30388
rect 46523 30348 46572 30376
rect 46523 30345 46535 30348
rect 46477 30339 46535 30345
rect 46566 30336 46572 30348
rect 46624 30336 46630 30388
rect 49602 30376 49608 30388
rect 49344 30348 49608 30376
rect 12676 30280 12940 30308
rect 38856 30280 39988 30308
rect 12676 30268 12682 30280
rect 10781 30243 10839 30249
rect 10781 30209 10793 30243
rect 10827 30209 10839 30243
rect 10781 30203 10839 30209
rect 10870 30190 10876 30242
rect 10928 30190 10934 30242
rect 10980 30240 11008 30268
rect 38856 30249 38884 30280
rect 41414 30268 41420 30320
rect 41472 30268 41478 30320
rect 41969 30311 42027 30317
rect 41969 30277 41981 30311
rect 42015 30308 42027 30311
rect 42429 30311 42487 30317
rect 42429 30308 42441 30311
rect 42015 30280 42441 30308
rect 42015 30277 42027 30280
rect 41969 30271 42027 30277
rect 42429 30277 42441 30280
rect 42475 30277 42487 30311
rect 43088 30308 43116 30336
rect 43088 30280 43668 30308
rect 42429 30271 42487 30277
rect 11057 30243 11115 30249
rect 11057 30240 11069 30243
rect 10980 30212 11069 30240
rect 11057 30209 11069 30212
rect 11103 30209 11115 30243
rect 11773 30243 11831 30249
rect 11773 30240 11785 30243
rect 11057 30203 11115 30209
rect 11164 30212 11785 30240
rect 9646 30144 10456 30172
rect 10410 30064 10416 30116
rect 10468 30064 10474 30116
rect 11164 30104 11192 30212
rect 11773 30209 11785 30212
rect 11819 30209 11831 30243
rect 11773 30203 11831 30209
rect 38841 30243 38899 30249
rect 38841 30209 38853 30243
rect 38887 30209 38899 30243
rect 38841 30203 38899 30209
rect 39206 30200 39212 30252
rect 39264 30200 39270 30252
rect 39390 30200 39396 30252
rect 39448 30200 39454 30252
rect 39482 30200 39488 30252
rect 39540 30240 39546 30252
rect 40129 30243 40187 30249
rect 40129 30240 40141 30243
rect 39540 30212 40141 30240
rect 39540 30200 39546 30212
rect 40129 30209 40141 30212
rect 40175 30240 40187 30243
rect 40402 30240 40408 30252
rect 40175 30212 40408 30240
rect 40175 30209 40187 30212
rect 40129 30203 40187 30209
rect 40402 30200 40408 30212
rect 40460 30200 40466 30252
rect 42794 30200 42800 30252
rect 42852 30240 42858 30252
rect 43257 30243 43315 30249
rect 43257 30240 43269 30243
rect 42852 30212 43269 30240
rect 42852 30200 42858 30212
rect 43257 30209 43269 30212
rect 43303 30209 43315 30243
rect 43257 30203 43315 30209
rect 43346 30200 43352 30252
rect 43404 30200 43410 30252
rect 43640 30249 43668 30280
rect 47302 30268 47308 30320
rect 47360 30308 47366 30320
rect 48685 30311 48743 30317
rect 47360 30280 48544 30308
rect 47360 30268 47366 30280
rect 43625 30243 43683 30249
rect 43625 30209 43637 30243
rect 43671 30240 43683 30243
rect 43901 30243 43959 30249
rect 43901 30240 43913 30243
rect 43671 30212 43913 30240
rect 43671 30209 43683 30212
rect 43625 30203 43683 30209
rect 43901 30209 43913 30212
rect 43947 30209 43959 30243
rect 43901 30203 43959 30209
rect 44085 30243 44143 30249
rect 44085 30209 44097 30243
rect 44131 30209 44143 30243
rect 44085 30203 44143 30209
rect 11514 30132 11520 30184
rect 11572 30132 11578 30184
rect 15378 30132 15384 30184
rect 15436 30172 15442 30184
rect 40497 30175 40555 30181
rect 15436 30144 40080 30172
rect 15436 30132 15442 30144
rect 10612 30076 11192 30104
rect 4948 30008 5764 30036
rect 4948 29996 4954 30008
rect 7466 29996 7472 30048
rect 7524 30036 7530 30048
rect 7745 30039 7803 30045
rect 7745 30036 7757 30039
rect 7524 30008 7757 30036
rect 7524 29996 7530 30008
rect 7745 30005 7757 30008
rect 7791 30005 7803 30039
rect 7745 29999 7803 30005
rect 9214 29996 9220 30048
rect 9272 30036 9278 30048
rect 9493 30039 9551 30045
rect 9493 30036 9505 30039
rect 9272 30008 9505 30036
rect 9272 29996 9278 30008
rect 9493 30005 9505 30008
rect 9539 30005 9551 30039
rect 9493 29999 9551 30005
rect 10505 30039 10563 30045
rect 10505 30005 10517 30039
rect 10551 30036 10563 30039
rect 10612 30036 10640 30076
rect 31018 30064 31024 30116
rect 31076 30104 31082 30116
rect 31076 30076 31754 30104
rect 31076 30064 31082 30076
rect 10551 30008 10640 30036
rect 10965 30039 11023 30045
rect 10551 30005 10563 30008
rect 10505 29999 10563 30005
rect 10965 30005 10977 30039
rect 11011 30036 11023 30039
rect 11054 30036 11060 30048
rect 11011 30008 11060 30036
rect 11011 30005 11023 30008
rect 10965 29999 11023 30005
rect 11054 29996 11060 30008
rect 11112 29996 11118 30048
rect 31726 30036 31754 30076
rect 37366 30064 37372 30116
rect 37424 30104 37430 30116
rect 38286 30104 38292 30116
rect 37424 30076 38292 30104
rect 37424 30064 37430 30076
rect 38286 30064 38292 30076
rect 38344 30104 38350 30116
rect 38749 30107 38807 30113
rect 38749 30104 38761 30107
rect 38344 30076 38761 30104
rect 38344 30064 38350 30076
rect 38749 30073 38761 30076
rect 38795 30073 38807 30107
rect 38749 30067 38807 30073
rect 38654 30036 38660 30048
rect 31726 30008 38660 30036
rect 38654 29996 38660 30008
rect 38712 29996 38718 30048
rect 38930 29996 38936 30048
rect 38988 30036 38994 30048
rect 39393 30039 39451 30045
rect 39393 30036 39405 30039
rect 38988 30008 39405 30036
rect 38988 29996 38994 30008
rect 39393 30005 39405 30008
rect 39439 30036 39451 30039
rect 39758 30036 39764 30048
rect 39439 30008 39764 30036
rect 39439 30005 39451 30008
rect 39393 29999 39451 30005
rect 39758 29996 39764 30008
rect 39816 29996 39822 30048
rect 40052 30036 40080 30144
rect 40497 30141 40509 30175
rect 40543 30172 40555 30175
rect 41966 30172 41972 30184
rect 40543 30144 41972 30172
rect 40543 30141 40555 30144
rect 40497 30135 40555 30141
rect 41966 30132 41972 30144
rect 42024 30132 42030 30184
rect 42245 30175 42303 30181
rect 42245 30141 42257 30175
rect 42291 30172 42303 30175
rect 42518 30172 42524 30184
rect 42291 30144 42524 30172
rect 42291 30141 42303 30144
rect 42245 30135 42303 30141
rect 42518 30132 42524 30144
rect 42576 30132 42582 30184
rect 43073 30175 43131 30181
rect 43073 30141 43085 30175
rect 43119 30172 43131 30175
rect 43119 30144 43208 30172
rect 43119 30141 43131 30144
rect 43073 30135 43131 30141
rect 43180 30113 43208 30144
rect 43990 30132 43996 30184
rect 44048 30172 44054 30184
rect 44100 30172 44128 30203
rect 44174 30200 44180 30252
rect 44232 30200 44238 30252
rect 45649 30243 45707 30249
rect 45649 30240 45661 30243
rect 45388 30212 45661 30240
rect 44048 30144 45324 30172
rect 44048 30132 44054 30144
rect 45296 30113 45324 30144
rect 43165 30107 43223 30113
rect 43165 30073 43177 30107
rect 43211 30073 43223 30107
rect 43165 30067 43223 30073
rect 45281 30107 45339 30113
rect 45281 30073 45293 30107
rect 45327 30073 45339 30107
rect 45281 30067 45339 30073
rect 43438 30036 43444 30048
rect 40052 30008 43444 30036
rect 43438 29996 43444 30008
rect 43496 29996 43502 30048
rect 43530 29996 43536 30048
rect 43588 29996 43594 30048
rect 45094 29996 45100 30048
rect 45152 30036 45158 30048
rect 45388 30036 45416 30212
rect 45649 30209 45661 30212
rect 45695 30209 45707 30243
rect 45649 30203 45707 30209
rect 48406 30200 48412 30252
rect 48464 30200 48470 30252
rect 48516 30240 48544 30280
rect 48685 30277 48697 30311
rect 48731 30308 48743 30311
rect 48958 30308 48964 30320
rect 48731 30280 48964 30308
rect 48731 30277 48743 30280
rect 48685 30271 48743 30277
rect 48958 30268 48964 30280
rect 49016 30268 49022 30320
rect 49344 30240 49372 30348
rect 49602 30336 49608 30348
rect 49660 30336 49666 30388
rect 51718 30376 51724 30388
rect 51460 30348 51724 30376
rect 50154 30268 50160 30320
rect 50212 30308 50218 30320
rect 50433 30311 50491 30317
rect 50433 30308 50445 30311
rect 50212 30280 50445 30308
rect 50212 30268 50218 30280
rect 50433 30277 50445 30280
rect 50479 30277 50491 30311
rect 50433 30271 50491 30277
rect 51460 30249 51488 30348
rect 51718 30336 51724 30348
rect 51776 30336 51782 30388
rect 53466 30336 53472 30388
rect 53524 30336 53530 30388
rect 57790 30376 57796 30388
rect 54772 30348 57796 30376
rect 51813 30311 51871 30317
rect 51813 30277 51825 30311
rect 51859 30308 51871 30311
rect 53009 30311 53067 30317
rect 51859 30280 52224 30308
rect 51859 30277 51871 30280
rect 51813 30271 51871 30277
rect 51629 30252 51687 30255
rect 48516 30226 49372 30240
rect 51445 30243 51503 30249
rect 48516 30212 49358 30226
rect 51445 30209 51457 30243
rect 51491 30209 51503 30243
rect 51445 30203 51503 30209
rect 51537 30243 51595 30249
rect 51537 30209 51549 30243
rect 51583 30209 51595 30243
rect 51537 30203 51595 30209
rect 45557 30175 45615 30181
rect 45557 30141 45569 30175
rect 45603 30172 45615 30175
rect 45738 30172 45744 30184
rect 45603 30144 45744 30172
rect 45603 30141 45615 30144
rect 45557 30135 45615 30141
rect 45738 30132 45744 30144
rect 45796 30132 45802 30184
rect 47026 30132 47032 30184
rect 47084 30132 47090 30184
rect 50709 30175 50767 30181
rect 50709 30141 50721 30175
rect 50755 30172 50767 30175
rect 50755 30144 51074 30172
rect 50755 30141 50767 30144
rect 50709 30135 50767 30141
rect 46014 30104 46020 30116
rect 45664 30076 46020 30104
rect 45664 30045 45692 30076
rect 46014 30064 46020 30076
rect 46072 30104 46078 30116
rect 46293 30107 46351 30113
rect 46293 30104 46305 30107
rect 46072 30076 46305 30104
rect 46072 30064 46078 30076
rect 46293 30073 46305 30076
rect 46339 30073 46351 30107
rect 46293 30067 46351 30073
rect 45152 30008 45416 30036
rect 45649 30039 45707 30045
rect 45152 29996 45158 30008
rect 45649 30005 45661 30039
rect 45695 30005 45707 30039
rect 45649 29999 45707 30005
rect 45738 29996 45744 30048
rect 45796 30036 45802 30048
rect 45925 30039 45983 30045
rect 45925 30036 45937 30039
rect 45796 30008 45937 30036
rect 45796 29996 45802 30008
rect 45925 30005 45937 30008
rect 45971 30005 45983 30039
rect 45925 29999 45983 30005
rect 47854 29996 47860 30048
rect 47912 29996 47918 30048
rect 51046 30036 51074 30144
rect 51542 30104 51570 30203
rect 51626 30200 51632 30252
rect 51684 30246 51690 30252
rect 51684 30218 51723 30246
rect 51905 30243 51963 30249
rect 51684 30200 51690 30218
rect 51905 30209 51917 30243
rect 51951 30209 51963 30243
rect 51905 30203 51963 30209
rect 51810 30132 51816 30184
rect 51868 30132 51874 30184
rect 51828 30104 51856 30132
rect 51542 30076 51856 30104
rect 51920 30104 51948 30203
rect 52086 30200 52092 30252
rect 52144 30200 52150 30252
rect 52196 30249 52224 30280
rect 53009 30277 53021 30311
rect 53055 30308 53067 30311
rect 53055 30280 53420 30308
rect 53055 30277 53067 30280
rect 53009 30271 53067 30277
rect 52181 30243 52239 30249
rect 52181 30209 52193 30243
rect 52227 30209 52239 30243
rect 52181 30203 52239 30209
rect 52365 30243 52423 30249
rect 52365 30209 52377 30243
rect 52411 30209 52423 30243
rect 52365 30203 52423 30209
rect 51997 30175 52055 30181
rect 51997 30141 52009 30175
rect 52043 30172 52055 30175
rect 52380 30172 52408 30203
rect 52914 30200 52920 30252
rect 52972 30200 52978 30252
rect 53101 30243 53159 30249
rect 53101 30209 53113 30243
rect 53147 30240 53159 30243
rect 53190 30240 53196 30252
rect 53147 30212 53196 30240
rect 53147 30209 53159 30212
rect 53101 30203 53159 30209
rect 53190 30200 53196 30212
rect 53248 30200 53254 30252
rect 53285 30243 53343 30249
rect 53285 30209 53297 30243
rect 53331 30238 53343 30243
rect 53392 30238 53420 30280
rect 53484 30249 53512 30336
rect 53558 30268 53564 30320
rect 53616 30308 53622 30320
rect 54772 30308 54800 30348
rect 57790 30336 57796 30348
rect 57848 30336 57854 30388
rect 53616 30280 54800 30308
rect 53616 30268 53622 30280
rect 53331 30210 53420 30238
rect 53469 30243 53527 30249
rect 53331 30209 53343 30210
rect 53285 30203 53343 30209
rect 53469 30209 53481 30243
rect 53515 30209 53527 30243
rect 53469 30203 53527 30209
rect 54294 30200 54300 30252
rect 54352 30200 54358 30252
rect 54481 30243 54539 30249
rect 54481 30209 54493 30243
rect 54527 30240 54539 30243
rect 54662 30240 54668 30252
rect 54527 30212 54668 30240
rect 54527 30209 54539 30212
rect 54481 30203 54539 30209
rect 54662 30200 54668 30212
rect 54720 30200 54726 30252
rect 54772 30249 54800 30280
rect 54846 30268 54852 30320
rect 54904 30308 54910 30320
rect 57609 30311 57667 30317
rect 57609 30308 57621 30311
rect 54904 30280 55352 30308
rect 54904 30268 54910 30280
rect 54956 30249 54984 30280
rect 55324 30264 55352 30280
rect 55784 30280 57621 30308
rect 54757 30243 54815 30249
rect 54757 30209 54769 30243
rect 54803 30209 54815 30243
rect 54757 30203 54815 30209
rect 54941 30243 54999 30249
rect 54941 30209 54953 30243
rect 54987 30209 54999 30243
rect 54941 30203 54999 30209
rect 55214 30200 55220 30252
rect 55272 30200 55278 30252
rect 55324 30240 55444 30264
rect 55784 30240 55812 30280
rect 57609 30277 57621 30280
rect 57655 30277 57667 30311
rect 57609 30271 57667 30277
rect 57716 30280 58572 30308
rect 55324 30236 55812 30240
rect 55416 30212 55812 30236
rect 57514 30200 57520 30252
rect 57572 30200 57578 30252
rect 52043 30144 52408 30172
rect 52043 30141 52055 30144
rect 51997 30135 52055 30141
rect 54570 30132 54576 30184
rect 54628 30172 54634 30184
rect 57716 30172 57744 30280
rect 58544 30252 58572 30280
rect 57885 30243 57943 30249
rect 57885 30209 57897 30243
rect 57931 30209 57943 30243
rect 57885 30203 57943 30209
rect 54628 30144 57744 30172
rect 57900 30172 57928 30203
rect 58066 30200 58072 30252
rect 58124 30240 58130 30252
rect 58161 30243 58219 30249
rect 58161 30240 58173 30243
rect 58124 30212 58173 30240
rect 58124 30200 58130 30212
rect 58161 30209 58173 30212
rect 58207 30209 58219 30243
rect 58161 30203 58219 30209
rect 58526 30200 58532 30252
rect 58584 30200 58590 30252
rect 57900 30144 58664 30172
rect 54628 30132 54634 30144
rect 58636 30116 58664 30144
rect 51920 30076 52040 30104
rect 52012 30048 52040 30076
rect 52086 30064 52092 30116
rect 52144 30104 52150 30116
rect 58253 30107 58311 30113
rect 58253 30104 58265 30107
rect 52144 30076 58265 30104
rect 52144 30064 52150 30076
rect 58253 30073 58265 30076
rect 58299 30073 58311 30107
rect 58253 30067 58311 30073
rect 58618 30064 58624 30116
rect 58676 30064 58682 30116
rect 51902 30036 51908 30048
rect 51046 30008 51908 30036
rect 51902 29996 51908 30008
rect 51960 29996 51966 30048
rect 51994 29996 52000 30048
rect 52052 29996 52058 30048
rect 52178 29996 52184 30048
rect 52236 30036 52242 30048
rect 52273 30039 52331 30045
rect 52273 30036 52285 30039
rect 52236 30008 52285 30036
rect 52236 29996 52242 30008
rect 52273 30005 52285 30008
rect 52319 30005 52331 30039
rect 52273 29999 52331 30005
rect 53374 29996 53380 30048
rect 53432 29996 53438 30048
rect 54386 29996 54392 30048
rect 54444 29996 54450 30048
rect 54662 29996 54668 30048
rect 54720 30036 54726 30048
rect 54849 30039 54907 30045
rect 54849 30036 54861 30039
rect 54720 30008 54861 30036
rect 54720 29996 54726 30008
rect 54849 30005 54861 30008
rect 54895 30005 54907 30039
rect 54849 29999 54907 30005
rect 55858 29996 55864 30048
rect 55916 29996 55922 30048
rect 58066 29996 58072 30048
rect 58124 29996 58130 30048
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 3602 29792 3608 29844
rect 3660 29792 3666 29844
rect 3694 29792 3700 29844
rect 3752 29832 3758 29844
rect 3789 29835 3847 29841
rect 3789 29832 3801 29835
rect 3752 29804 3801 29832
rect 3752 29792 3758 29804
rect 3789 29801 3801 29804
rect 3835 29801 3847 29835
rect 3789 29795 3847 29801
rect 4062 29792 4068 29844
rect 4120 29832 4126 29844
rect 4617 29835 4675 29841
rect 4617 29832 4629 29835
rect 4120 29804 4629 29832
rect 4120 29792 4126 29804
rect 4617 29801 4629 29804
rect 4663 29801 4675 29835
rect 5074 29832 5080 29844
rect 4617 29795 4675 29801
rect 4715 29804 5080 29832
rect 3620 29705 3648 29792
rect 3605 29699 3663 29705
rect 3605 29665 3617 29699
rect 3651 29665 3663 29699
rect 4715 29696 4743 29804
rect 5074 29792 5080 29804
rect 5132 29792 5138 29844
rect 5902 29792 5908 29844
rect 5960 29832 5966 29844
rect 5997 29835 6055 29841
rect 5997 29832 6009 29835
rect 5960 29804 6009 29832
rect 5960 29792 5966 29804
rect 5997 29801 6009 29804
rect 6043 29801 6055 29835
rect 5997 29795 6055 29801
rect 6549 29835 6607 29841
rect 6549 29801 6561 29835
rect 6595 29832 6607 29835
rect 6638 29832 6644 29844
rect 6595 29804 6644 29832
rect 6595 29801 6607 29804
rect 6549 29795 6607 29801
rect 6638 29792 6644 29804
rect 6696 29792 6702 29844
rect 6730 29792 6736 29844
rect 6788 29832 6794 29844
rect 6788 29804 15056 29832
rect 6788 29792 6794 29804
rect 15028 29776 15056 29804
rect 15838 29792 15844 29844
rect 15896 29792 15902 29844
rect 31018 29832 31024 29844
rect 26206 29804 31024 29832
rect 5166 29724 5172 29776
rect 5224 29764 5230 29776
rect 9769 29767 9827 29773
rect 9769 29764 9781 29767
rect 5224 29736 8156 29764
rect 5224 29724 5230 29736
rect 4890 29696 4896 29708
rect 3605 29659 3663 29665
rect 4540 29668 4743 29696
rect 4816 29668 4896 29696
rect 4540 29637 4568 29668
rect 2593 29631 2651 29637
rect 2593 29628 2605 29631
rect 2424 29600 2605 29628
rect 934 29520 940 29572
rect 992 29560 998 29572
rect 1581 29563 1639 29569
rect 1581 29560 1593 29563
rect 992 29532 1593 29560
rect 992 29520 998 29532
rect 1581 29529 1593 29532
rect 1627 29529 1639 29563
rect 1581 29523 1639 29529
rect 1394 29452 1400 29504
rect 1452 29492 1458 29504
rect 2424 29492 2452 29600
rect 2593 29597 2605 29600
rect 2639 29597 2651 29631
rect 2593 29591 2651 29597
rect 4433 29631 4491 29637
rect 4433 29597 4445 29631
rect 4479 29597 4491 29631
rect 4433 29591 4491 29597
rect 4525 29631 4583 29637
rect 4525 29597 4537 29631
rect 4571 29597 4583 29631
rect 4525 29591 4583 29597
rect 4709 29631 4767 29637
rect 4709 29597 4721 29631
rect 4755 29628 4767 29631
rect 4816 29628 4844 29668
rect 4890 29656 4896 29668
rect 4948 29656 4954 29708
rect 6730 29656 6736 29708
rect 6788 29656 6794 29708
rect 8128 29705 8156 29736
rect 9646 29736 9781 29764
rect 7009 29699 7067 29705
rect 7009 29696 7021 29699
rect 6840 29668 7021 29696
rect 6748 29628 6776 29656
rect 6840 29637 6868 29668
rect 7009 29665 7021 29668
rect 7055 29665 7067 29699
rect 7009 29659 7067 29665
rect 8113 29699 8171 29705
rect 8113 29665 8125 29699
rect 8159 29665 8171 29699
rect 8113 29659 8171 29665
rect 9122 29656 9128 29708
rect 9180 29656 9186 29708
rect 4755 29600 4844 29628
rect 4908 29600 6776 29628
rect 6825 29631 6883 29637
rect 4755 29597 4767 29600
rect 4709 29591 4767 29597
rect 4448 29560 4476 29591
rect 4798 29560 4804 29572
rect 4448 29532 4804 29560
rect 4798 29520 4804 29532
rect 4856 29520 4862 29572
rect 1452 29464 2452 29492
rect 1452 29452 1458 29464
rect 2958 29452 2964 29504
rect 3016 29452 3022 29504
rect 3142 29452 3148 29504
rect 3200 29492 3206 29504
rect 4908 29492 4936 29600
rect 6825 29597 6837 29631
rect 6871 29597 6883 29631
rect 6825 29591 6883 29597
rect 6917 29631 6975 29637
rect 6917 29597 6929 29631
rect 6963 29597 6975 29631
rect 6917 29591 6975 29597
rect 7101 29631 7159 29637
rect 7101 29597 7113 29631
rect 7147 29628 7159 29631
rect 8665 29631 8723 29637
rect 7147 29600 7512 29628
rect 7147 29597 7159 29600
rect 7101 29591 7159 29597
rect 5810 29520 5816 29572
rect 5868 29560 5874 29572
rect 6546 29560 6552 29572
rect 5868 29532 6552 29560
rect 5868 29520 5874 29532
rect 6546 29520 6552 29532
rect 6604 29520 6610 29572
rect 6932 29504 6960 29591
rect 7484 29504 7512 29600
rect 8665 29597 8677 29631
rect 8711 29628 8723 29631
rect 8938 29628 8944 29640
rect 8711 29600 8944 29628
rect 8711 29597 8723 29600
rect 8665 29591 8723 29597
rect 8938 29588 8944 29600
rect 8996 29628 9002 29640
rect 9401 29631 9459 29637
rect 9401 29628 9413 29631
rect 8996 29600 9413 29628
rect 8996 29588 9002 29600
rect 9401 29597 9413 29600
rect 9447 29628 9459 29631
rect 9646 29628 9674 29736
rect 9769 29733 9781 29736
rect 9815 29764 9827 29767
rect 10226 29764 10232 29776
rect 9815 29736 10232 29764
rect 9815 29733 9827 29736
rect 9769 29727 9827 29733
rect 10226 29724 10232 29736
rect 10284 29764 10290 29776
rect 10284 29736 12480 29764
rect 10284 29724 10290 29736
rect 12452 29696 12480 29736
rect 15010 29724 15016 29776
rect 15068 29724 15074 29776
rect 26206 29764 26234 29804
rect 31018 29792 31024 29804
rect 31076 29792 31082 29844
rect 39942 29832 39948 29844
rect 37384 29804 39948 29832
rect 37384 29764 37412 29804
rect 39942 29792 39948 29804
rect 40000 29792 40006 29844
rect 40037 29835 40095 29841
rect 40037 29801 40049 29835
rect 40083 29832 40095 29835
rect 41322 29832 41328 29844
rect 40083 29804 41328 29832
rect 40083 29801 40095 29804
rect 40037 29795 40095 29801
rect 41322 29792 41328 29804
rect 41380 29792 41386 29844
rect 43257 29835 43315 29841
rect 43257 29801 43269 29835
rect 43303 29832 43315 29835
rect 43530 29832 43536 29844
rect 43303 29804 43536 29832
rect 43303 29801 43315 29804
rect 43257 29795 43315 29801
rect 15120 29736 26234 29764
rect 31726 29736 37412 29764
rect 15120 29696 15148 29736
rect 10612 29668 11652 29696
rect 12452 29668 15148 29696
rect 9447 29600 9674 29628
rect 9447 29597 9459 29600
rect 9401 29591 9459 29597
rect 9766 29588 9772 29640
rect 9824 29628 9830 29640
rect 10612 29637 10640 29668
rect 10597 29631 10655 29637
rect 10597 29628 10609 29631
rect 9824 29600 10609 29628
rect 9824 29588 9830 29600
rect 10597 29597 10609 29600
rect 10643 29597 10655 29631
rect 10597 29591 10655 29597
rect 10781 29631 10839 29637
rect 10781 29597 10793 29631
rect 10827 29628 10839 29631
rect 10870 29628 10876 29640
rect 10827 29600 10876 29628
rect 10827 29597 10839 29600
rect 10781 29591 10839 29597
rect 9950 29520 9956 29572
rect 10008 29560 10014 29572
rect 10796 29560 10824 29591
rect 10870 29588 10876 29600
rect 10928 29588 10934 29640
rect 11624 29572 11652 29668
rect 15838 29656 15844 29708
rect 15896 29656 15902 29708
rect 31726 29696 31754 29736
rect 38654 29724 38660 29776
rect 38712 29764 38718 29776
rect 41785 29767 41843 29773
rect 41785 29764 41797 29767
rect 38712 29736 41797 29764
rect 38712 29724 38718 29736
rect 41785 29733 41797 29736
rect 41831 29733 41843 29767
rect 43272 29764 43300 29795
rect 43530 29792 43536 29804
rect 43588 29792 43594 29844
rect 43717 29835 43775 29841
rect 43717 29801 43729 29835
rect 43763 29832 43775 29835
rect 44174 29832 44180 29844
rect 43763 29804 44180 29832
rect 43763 29801 43775 29804
rect 43717 29795 43775 29801
rect 44174 29792 44180 29804
rect 44232 29792 44238 29844
rect 46753 29835 46811 29841
rect 45112 29804 46704 29832
rect 41785 29727 41843 29733
rect 42444 29736 43300 29764
rect 22066 29668 31754 29696
rect 11882 29588 11888 29640
rect 11940 29588 11946 29640
rect 15473 29631 15531 29637
rect 15473 29597 15485 29631
rect 15519 29628 15531 29631
rect 15856 29628 15884 29656
rect 15519 29600 15884 29628
rect 15519 29597 15531 29600
rect 15473 29591 15531 29597
rect 10008 29532 10824 29560
rect 10008 29520 10014 29532
rect 11606 29520 11612 29572
rect 11664 29520 11670 29572
rect 12434 29520 12440 29572
rect 12492 29560 12498 29572
rect 22066 29560 22094 29668
rect 36262 29656 36268 29708
rect 36320 29696 36326 29708
rect 37182 29696 37188 29708
rect 36320 29668 37188 29696
rect 36320 29656 36326 29668
rect 37182 29656 37188 29668
rect 37240 29696 37246 29708
rect 37277 29699 37335 29705
rect 37277 29696 37289 29699
rect 37240 29668 37289 29696
rect 37240 29656 37246 29668
rect 37277 29665 37289 29668
rect 37323 29696 37335 29699
rect 37369 29699 37427 29705
rect 37369 29696 37381 29699
rect 37323 29668 37381 29696
rect 37323 29665 37335 29668
rect 37277 29659 37335 29665
rect 37369 29665 37381 29668
rect 37415 29665 37427 29699
rect 37369 29659 37427 29665
rect 39390 29656 39396 29708
rect 39448 29696 39454 29708
rect 39448 29668 39528 29696
rect 39448 29656 39454 29668
rect 39500 29637 39528 29668
rect 39574 29656 39580 29708
rect 39632 29656 39638 29708
rect 40034 29696 40040 29708
rect 39684 29668 40040 29696
rect 39684 29637 39712 29668
rect 40034 29656 40040 29668
rect 40092 29656 40098 29708
rect 39485 29631 39543 29637
rect 39485 29597 39497 29631
rect 39531 29597 39543 29631
rect 39485 29591 39543 29597
rect 39669 29631 39727 29637
rect 39669 29597 39681 29631
rect 39715 29597 39727 29631
rect 39669 29591 39727 29597
rect 39758 29588 39764 29640
rect 39816 29628 39822 29640
rect 39945 29631 40003 29637
rect 39945 29628 39957 29631
rect 39816 29600 39957 29628
rect 39816 29588 39822 29600
rect 39945 29597 39957 29600
rect 39991 29597 40003 29631
rect 40052 29628 40080 29656
rect 40129 29631 40187 29637
rect 40129 29628 40141 29631
rect 40052 29600 40141 29628
rect 39945 29591 40003 29597
rect 40129 29597 40141 29600
rect 40175 29597 40187 29631
rect 40129 29591 40187 29597
rect 41966 29588 41972 29640
rect 42024 29588 42030 29640
rect 42444 29637 42472 29736
rect 43438 29724 43444 29776
rect 43496 29764 43502 29776
rect 45112 29764 45140 29804
rect 43496 29736 45140 29764
rect 46676 29764 46704 29804
rect 46753 29801 46765 29835
rect 46799 29832 46811 29835
rect 47026 29832 47032 29844
rect 46799 29804 47032 29832
rect 46799 29801 46811 29804
rect 46753 29795 46811 29801
rect 47026 29792 47032 29804
rect 47084 29792 47090 29844
rect 47118 29792 47124 29844
rect 47176 29832 47182 29844
rect 50893 29835 50951 29841
rect 50893 29832 50905 29835
rect 47176 29804 50905 29832
rect 47176 29792 47182 29804
rect 50893 29801 50905 29804
rect 50939 29801 50951 29835
rect 50893 29795 50951 29801
rect 51353 29835 51411 29841
rect 51353 29801 51365 29835
rect 51399 29832 51411 29835
rect 51810 29832 51816 29844
rect 51399 29804 51816 29832
rect 51399 29801 51411 29804
rect 51353 29795 51411 29801
rect 51810 29792 51816 29804
rect 51868 29792 51874 29844
rect 52086 29792 52092 29844
rect 52144 29832 52150 29844
rect 53190 29832 53196 29844
rect 52144 29804 53196 29832
rect 52144 29792 52150 29804
rect 53190 29792 53196 29804
rect 53248 29792 53254 29844
rect 53374 29792 53380 29844
rect 53432 29792 53438 29844
rect 55033 29835 55091 29841
rect 55033 29801 55045 29835
rect 55079 29832 55091 29835
rect 55214 29832 55220 29844
rect 55079 29804 55220 29832
rect 55079 29801 55091 29804
rect 55033 29795 55091 29801
rect 55214 29792 55220 29804
rect 55272 29792 55278 29844
rect 56502 29792 56508 29844
rect 56560 29832 56566 29844
rect 56560 29804 56732 29832
rect 56560 29792 56566 29804
rect 47305 29767 47363 29773
rect 47305 29764 47317 29767
rect 46676 29736 47317 29764
rect 43496 29724 43502 29736
rect 45005 29699 45063 29705
rect 45005 29696 45017 29699
rect 42536 29668 45017 29696
rect 42536 29640 42564 29668
rect 45005 29665 45017 29668
rect 45051 29696 45063 29699
rect 45646 29696 45652 29708
rect 45051 29668 45652 29696
rect 45051 29665 45063 29668
rect 45005 29659 45063 29665
rect 45646 29656 45652 29668
rect 45704 29656 45710 29708
rect 42429 29631 42487 29637
rect 42429 29597 42441 29631
rect 42475 29597 42487 29631
rect 42429 29591 42487 29597
rect 42518 29588 42524 29640
rect 42576 29588 42582 29640
rect 42981 29631 43039 29637
rect 42981 29597 42993 29631
rect 43027 29597 43039 29631
rect 42981 29591 43039 29597
rect 43165 29631 43223 29637
rect 43165 29597 43177 29631
rect 43211 29597 43223 29631
rect 43165 29591 43223 29597
rect 43349 29631 43407 29637
rect 43349 29597 43361 29631
rect 43395 29628 43407 29631
rect 43990 29628 43996 29640
rect 43395 29600 43996 29628
rect 43395 29597 43407 29600
rect 43349 29591 43407 29597
rect 12492 29532 22094 29560
rect 12492 29520 12498 29532
rect 37642 29520 37648 29572
rect 37700 29520 37706 29572
rect 40954 29560 40960 29572
rect 38870 29532 40960 29560
rect 40954 29520 40960 29532
rect 41012 29560 41018 29572
rect 41414 29560 41420 29572
rect 41012 29532 41420 29560
rect 41012 29520 41018 29532
rect 41414 29520 41420 29532
rect 41472 29520 41478 29572
rect 3200 29464 4936 29492
rect 3200 29452 3206 29464
rect 6730 29452 6736 29504
rect 6788 29452 6794 29504
rect 6914 29452 6920 29504
rect 6972 29452 6978 29504
rect 7466 29452 7472 29504
rect 7524 29452 7530 29504
rect 10781 29495 10839 29501
rect 10781 29461 10793 29495
rect 10827 29492 10839 29495
rect 11146 29492 11152 29504
rect 10827 29464 11152 29492
rect 10827 29461 10839 29464
rect 10781 29455 10839 29461
rect 11146 29452 11152 29464
rect 11204 29452 11210 29504
rect 15378 29452 15384 29504
rect 15436 29452 15442 29504
rect 37458 29452 37464 29504
rect 37516 29492 37522 29504
rect 38930 29492 38936 29504
rect 37516 29464 38936 29492
rect 37516 29452 37522 29464
rect 38930 29452 38936 29464
rect 38988 29452 38994 29504
rect 39117 29495 39175 29501
rect 39117 29461 39129 29495
rect 39163 29492 39175 29495
rect 39482 29492 39488 29504
rect 39163 29464 39488 29492
rect 39163 29461 39175 29464
rect 39117 29455 39175 29461
rect 39482 29452 39488 29464
rect 39540 29452 39546 29504
rect 39574 29452 39580 29504
rect 39632 29492 39638 29504
rect 40034 29492 40040 29504
rect 39632 29464 40040 29492
rect 39632 29452 39638 29464
rect 40034 29452 40040 29464
rect 40092 29452 40098 29504
rect 42996 29492 43024 29591
rect 43180 29560 43208 29591
rect 43990 29588 43996 29600
rect 44048 29588 44054 29640
rect 44085 29631 44143 29637
rect 44085 29597 44097 29631
rect 44131 29628 44143 29631
rect 44818 29628 44824 29640
rect 44131 29600 44824 29628
rect 44131 29597 44143 29600
rect 44085 29591 44143 29597
rect 44818 29588 44824 29600
rect 44876 29588 44882 29640
rect 43622 29560 43628 29572
rect 43180 29532 43628 29560
rect 43622 29520 43628 29532
rect 43680 29560 43686 29572
rect 43901 29563 43959 29569
rect 43901 29560 43913 29563
rect 43680 29532 43913 29560
rect 43680 29520 43686 29532
rect 43901 29529 43913 29532
rect 43947 29529 43959 29563
rect 43901 29523 43959 29529
rect 44542 29520 44548 29572
rect 44600 29560 44606 29572
rect 45281 29563 45339 29569
rect 45281 29560 45293 29563
rect 44600 29532 45293 29560
rect 44600 29520 44606 29532
rect 45281 29529 45293 29532
rect 45327 29529 45339 29563
rect 45281 29523 45339 29529
rect 43530 29492 43536 29504
rect 42996 29464 43536 29492
rect 43530 29452 43536 29464
rect 43588 29452 43594 29504
rect 46400 29492 46428 29614
rect 46566 29588 46572 29640
rect 46624 29588 46630 29640
rect 46676 29628 46704 29736
rect 47305 29733 47317 29736
rect 47351 29733 47363 29767
rect 47305 29727 47363 29733
rect 50154 29724 50160 29776
rect 50212 29724 50218 29776
rect 51994 29724 52000 29776
rect 52052 29724 52058 29776
rect 52104 29736 53052 29764
rect 47394 29656 47400 29708
rect 47452 29696 47458 29708
rect 47489 29699 47547 29705
rect 47489 29696 47501 29699
rect 47452 29668 47501 29696
rect 47452 29656 47458 29668
rect 47489 29665 47501 29668
rect 47535 29665 47547 29699
rect 47489 29659 47547 29665
rect 47765 29699 47823 29705
rect 47765 29665 47777 29699
rect 47811 29696 47823 29699
rect 47854 29696 47860 29708
rect 47811 29668 47860 29696
rect 47811 29665 47823 29668
rect 47765 29659 47823 29665
rect 47854 29656 47860 29668
rect 47912 29656 47918 29708
rect 48958 29656 48964 29708
rect 49016 29696 49022 29708
rect 50614 29696 50620 29708
rect 49016 29668 50620 29696
rect 49016 29656 49022 29668
rect 50614 29656 50620 29668
rect 50672 29696 50678 29708
rect 50709 29699 50767 29705
rect 50709 29696 50721 29699
rect 50672 29668 50721 29696
rect 50672 29656 50678 29668
rect 50709 29665 50721 29668
rect 50755 29665 50767 29699
rect 51169 29699 51227 29705
rect 51169 29696 51181 29699
rect 50709 29659 50767 29665
rect 50816 29668 51181 29696
rect 46845 29631 46903 29637
rect 46845 29628 46857 29631
rect 46676 29600 46857 29628
rect 46845 29597 46857 29600
rect 46891 29597 46903 29631
rect 46845 29591 46903 29597
rect 47029 29631 47087 29637
rect 47029 29597 47041 29631
rect 47075 29597 47087 29631
rect 47029 29591 47087 29597
rect 46584 29560 46612 29588
rect 47044 29560 47072 29591
rect 47302 29588 47308 29640
rect 47360 29588 47366 29640
rect 49970 29588 49976 29640
rect 50028 29628 50034 29640
rect 50816 29628 50844 29668
rect 51169 29665 51181 29668
rect 51215 29665 51227 29699
rect 52012 29696 52040 29724
rect 51169 29659 51227 29665
rect 51368 29668 52040 29696
rect 50028 29600 50844 29628
rect 50028 29588 50034 29600
rect 51074 29588 51080 29640
rect 51132 29628 51138 29640
rect 51368 29628 51396 29668
rect 51132 29600 51396 29628
rect 51132 29588 51138 29600
rect 51442 29588 51448 29640
rect 51500 29588 51506 29640
rect 51721 29631 51779 29637
rect 51721 29597 51733 29631
rect 51767 29628 51779 29631
rect 51810 29628 51816 29640
rect 51767 29600 51816 29628
rect 51767 29597 51779 29600
rect 51721 29591 51779 29597
rect 51810 29588 51816 29600
rect 51868 29588 51874 29640
rect 51997 29631 52055 29637
rect 51997 29597 52009 29631
rect 52043 29628 52055 29631
rect 52104 29628 52132 29736
rect 52043 29600 52132 29628
rect 52043 29597 52055 29600
rect 51997 29591 52055 29597
rect 46584 29532 47072 29560
rect 47320 29560 47348 29588
rect 47320 29532 48254 29560
rect 51350 29520 51356 29572
rect 51408 29560 51414 29572
rect 51534 29560 51540 29572
rect 51408 29532 51540 29560
rect 51408 29520 51414 29532
rect 51534 29520 51540 29532
rect 51592 29520 51598 29572
rect 46566 29492 46572 29504
rect 46400 29464 46572 29492
rect 46566 29452 46572 29464
rect 46624 29452 46630 29504
rect 46842 29452 46848 29504
rect 46900 29492 46906 29504
rect 46937 29495 46995 29501
rect 46937 29492 46949 29495
rect 46900 29464 46949 29492
rect 46900 29452 46906 29464
rect 46937 29461 46949 29464
rect 46983 29461 46995 29495
rect 46937 29455 46995 29461
rect 49234 29452 49240 29504
rect 49292 29452 49298 29504
rect 49418 29452 49424 29504
rect 49476 29492 49482 29504
rect 52012 29492 52040 29591
rect 52178 29588 52184 29640
rect 52236 29588 52242 29640
rect 52281 29631 52339 29637
rect 52281 29597 52293 29631
rect 52327 29597 52339 29631
rect 52281 29591 52339 29597
rect 52089 29563 52147 29569
rect 52089 29529 52101 29563
rect 52135 29560 52147 29563
rect 52288 29560 52316 29591
rect 52454 29588 52460 29640
rect 52512 29588 52518 29640
rect 53024 29637 53052 29736
rect 53392 29696 53420 29792
rect 54021 29699 54079 29705
rect 54021 29696 54033 29699
rect 53208 29668 53420 29696
rect 53576 29668 54033 29696
rect 53208 29637 53236 29668
rect 53576 29640 53604 29668
rect 54021 29665 54033 29668
rect 54067 29665 54079 29699
rect 54021 29659 54079 29665
rect 54386 29656 54392 29708
rect 54444 29656 54450 29708
rect 55030 29656 55036 29708
rect 55088 29656 55094 29708
rect 56704 29705 56732 29804
rect 57514 29792 57520 29844
rect 57572 29792 57578 29844
rect 58710 29724 58716 29776
rect 58768 29724 58774 29776
rect 56689 29699 56747 29705
rect 56689 29665 56701 29699
rect 56735 29665 56747 29699
rect 58728 29696 58756 29724
rect 56689 29659 56747 29665
rect 57072 29668 58756 29696
rect 53009 29631 53067 29637
rect 53009 29597 53021 29631
rect 53055 29597 53067 29631
rect 53009 29591 53067 29597
rect 53193 29631 53251 29637
rect 53193 29597 53205 29631
rect 53239 29597 53251 29631
rect 53193 29591 53251 29597
rect 53285 29631 53343 29637
rect 53285 29597 53297 29631
rect 53331 29597 53343 29631
rect 53285 29591 53343 29597
rect 53469 29631 53527 29637
rect 53469 29597 53481 29631
rect 53515 29597 53527 29631
rect 53469 29591 53527 29597
rect 52135 29532 52316 29560
rect 52135 29529 52147 29532
rect 52089 29523 52147 29529
rect 53024 29504 53052 29591
rect 53101 29563 53159 29569
rect 53101 29529 53113 29563
rect 53147 29560 53159 29563
rect 53300 29560 53328 29591
rect 53147 29532 53328 29560
rect 53484 29560 53512 29591
rect 53558 29588 53564 29640
rect 53616 29588 53622 29640
rect 53745 29631 53803 29637
rect 53745 29597 53757 29631
rect 53791 29628 53803 29631
rect 54404 29628 54432 29656
rect 53791 29600 54432 29628
rect 54941 29631 54999 29637
rect 53791 29597 53803 29600
rect 53745 29591 53803 29597
rect 54941 29597 54953 29631
rect 54987 29628 54999 29631
rect 55048 29628 55076 29656
rect 54987 29600 55076 29628
rect 54987 29597 54999 29600
rect 54941 29591 54999 29597
rect 55122 29588 55128 29640
rect 55180 29588 55186 29640
rect 56962 29628 56968 29640
rect 55232 29600 56968 29628
rect 53653 29563 53711 29569
rect 53653 29560 53665 29563
rect 53484 29532 53665 29560
rect 53147 29529 53159 29532
rect 53101 29523 53159 29529
rect 53653 29529 53665 29532
rect 53699 29529 53711 29563
rect 53653 29523 53711 29529
rect 53834 29520 53840 29572
rect 53892 29560 53898 29572
rect 55232 29560 55260 29600
rect 56962 29588 56968 29600
rect 57020 29588 57026 29640
rect 53892 29532 55260 29560
rect 53892 29520 53898 29532
rect 56042 29520 56048 29572
rect 56100 29560 56106 29572
rect 56422 29563 56480 29569
rect 56422 29560 56434 29563
rect 56100 29532 56434 29560
rect 56100 29520 56106 29532
rect 56422 29529 56434 29532
rect 56468 29529 56480 29563
rect 57072 29560 57100 29668
rect 57149 29631 57207 29637
rect 57149 29597 57161 29631
rect 57195 29628 57207 29631
rect 57238 29628 57244 29640
rect 57195 29600 57244 29628
rect 57195 29597 57207 29600
rect 57149 29591 57207 29597
rect 57238 29588 57244 29600
rect 57296 29588 57302 29640
rect 57701 29631 57759 29637
rect 57701 29628 57713 29631
rect 57532 29600 57713 29628
rect 56422 29523 56480 29529
rect 56520 29532 57100 29560
rect 49476 29464 52040 29492
rect 49476 29452 49482 29464
rect 52270 29452 52276 29504
rect 52328 29452 52334 29504
rect 52825 29495 52883 29501
rect 52825 29461 52837 29495
rect 52871 29492 52883 29495
rect 53006 29492 53012 29504
rect 52871 29464 53012 29492
rect 52871 29461 52883 29464
rect 52825 29455 52883 29461
rect 53006 29452 53012 29464
rect 53064 29452 53070 29504
rect 53377 29495 53435 29501
rect 53377 29461 53389 29495
rect 53423 29492 53435 29495
rect 53558 29492 53564 29504
rect 53423 29464 53564 29492
rect 53423 29461 53435 29464
rect 53377 29455 53435 29461
rect 53558 29452 53564 29464
rect 53616 29452 53622 29504
rect 55306 29452 55312 29504
rect 55364 29452 55370 29504
rect 55398 29452 55404 29504
rect 55456 29492 55462 29504
rect 56520 29492 56548 29532
rect 55456 29464 56548 29492
rect 55456 29452 55462 29464
rect 57054 29452 57060 29504
rect 57112 29452 57118 29504
rect 57532 29492 57560 29600
rect 57701 29597 57713 29600
rect 57747 29597 57759 29631
rect 57701 29591 57759 29597
rect 57790 29588 57796 29640
rect 57848 29628 57854 29640
rect 57885 29631 57943 29637
rect 57885 29628 57897 29631
rect 57848 29600 57897 29628
rect 57848 29588 57854 29600
rect 57885 29597 57897 29600
rect 57931 29597 57943 29631
rect 57885 29591 57943 29597
rect 57606 29520 57612 29572
rect 57664 29560 57670 29572
rect 58253 29563 58311 29569
rect 58253 29560 58265 29563
rect 57664 29532 58265 29560
rect 57664 29520 57670 29532
rect 58253 29529 58265 29532
rect 58299 29529 58311 29563
rect 58253 29523 58311 29529
rect 58526 29492 58532 29504
rect 57532 29464 58532 29492
rect 58526 29452 58532 29464
rect 58584 29452 58590 29504
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 1394 29248 1400 29300
rect 1452 29288 1458 29300
rect 5442 29288 5448 29300
rect 1452 29260 3372 29288
rect 1452 29248 1458 29260
rect 2406 29180 2412 29232
rect 2464 29180 2470 29232
rect 2869 29223 2927 29229
rect 2869 29189 2881 29223
rect 2915 29220 2927 29223
rect 2958 29220 2964 29232
rect 2915 29192 2964 29220
rect 2915 29189 2927 29192
rect 2869 29183 2927 29189
rect 2958 29180 2964 29192
rect 3016 29180 3022 29232
rect 3145 29155 3203 29161
rect 3145 29121 3157 29155
rect 3191 29152 3203 29155
rect 3234 29152 3240 29164
rect 3191 29124 3240 29152
rect 3191 29121 3203 29124
rect 3145 29115 3203 29121
rect 3234 29112 3240 29124
rect 3292 29112 3298 29164
rect 3344 29161 3372 29260
rect 4172 29260 5448 29288
rect 4172 29161 4200 29260
rect 5442 29248 5448 29260
rect 5500 29288 5506 29300
rect 5813 29291 5871 29297
rect 5813 29288 5825 29291
rect 5500 29260 5825 29288
rect 5500 29248 5506 29260
rect 5813 29257 5825 29260
rect 5859 29288 5871 29291
rect 6454 29288 6460 29300
rect 5859 29260 6460 29288
rect 5859 29257 5871 29260
rect 5813 29251 5871 29257
rect 6454 29248 6460 29260
rect 6512 29248 6518 29300
rect 6549 29291 6607 29297
rect 6549 29257 6561 29291
rect 6595 29288 6607 29291
rect 6730 29288 6736 29300
rect 6595 29260 6736 29288
rect 6595 29257 6607 29260
rect 6549 29251 6607 29257
rect 6730 29248 6736 29260
rect 6788 29248 6794 29300
rect 8938 29248 8944 29300
rect 8996 29248 9002 29300
rect 10682 29291 10740 29297
rect 10682 29288 10694 29291
rect 10520 29260 10694 29288
rect 4706 29229 4712 29232
rect 4700 29183 4712 29229
rect 4764 29220 4770 29232
rect 4764 29192 4800 29220
rect 4706 29180 4712 29183
rect 4764 29180 4770 29192
rect 6270 29180 6276 29232
rect 6328 29220 6334 29232
rect 6328 29192 6776 29220
rect 6328 29180 6334 29192
rect 3329 29155 3387 29161
rect 3329 29121 3341 29155
rect 3375 29121 3387 29155
rect 3329 29115 3387 29121
rect 4157 29155 4215 29161
rect 4157 29121 4169 29155
rect 4203 29121 4215 29155
rect 4157 29115 4215 29121
rect 4341 29155 4399 29161
rect 4341 29121 4353 29155
rect 4387 29152 4399 29155
rect 4982 29152 4988 29164
rect 4387 29124 4988 29152
rect 4387 29121 4399 29124
rect 4341 29115 4399 29121
rect 4982 29112 4988 29124
rect 5040 29112 5046 29164
rect 5902 29112 5908 29164
rect 5960 29152 5966 29164
rect 6748 29161 6776 29192
rect 6914 29180 6920 29232
rect 6972 29220 6978 29232
rect 9950 29220 9956 29232
rect 6972 29192 9956 29220
rect 6972 29180 6978 29192
rect 9950 29180 9956 29192
rect 10008 29180 10014 29232
rect 10168 29223 10226 29229
rect 10168 29189 10180 29223
rect 10214 29220 10226 29223
rect 10520 29220 10548 29260
rect 10682 29257 10694 29260
rect 10728 29257 10740 29291
rect 10682 29251 10740 29257
rect 11072 29260 11192 29288
rect 11072 29232 11100 29260
rect 10214 29192 10548 29220
rect 10214 29189 10226 29192
rect 10168 29183 10226 29189
rect 10962 29180 10968 29232
rect 11020 29180 11026 29232
rect 11054 29180 11060 29232
rect 11112 29180 11118 29232
rect 11164 29229 11192 29260
rect 11606 29248 11612 29300
rect 11664 29248 11670 29300
rect 15010 29248 15016 29300
rect 15068 29288 15074 29300
rect 15068 29260 26234 29288
rect 15068 29248 15074 29260
rect 11149 29223 11207 29229
rect 11149 29189 11161 29223
rect 11195 29220 11207 29223
rect 11422 29220 11428 29232
rect 11195 29192 11428 29220
rect 11195 29189 11207 29192
rect 11149 29183 11207 29189
rect 11422 29180 11428 29192
rect 11480 29180 11486 29232
rect 6457 29155 6515 29161
rect 6457 29152 6469 29155
rect 5960 29124 6469 29152
rect 5960 29112 5966 29124
rect 6457 29121 6469 29124
rect 6503 29121 6515 29155
rect 6457 29115 6515 29121
rect 6733 29155 6791 29161
rect 6733 29121 6745 29155
rect 6779 29121 6791 29155
rect 6733 29115 6791 29121
rect 10502 29112 10508 29164
rect 10560 29112 10566 29164
rect 10594 29112 10600 29164
rect 10652 29112 10658 29164
rect 10686 29112 10692 29164
rect 10744 29158 10750 29164
rect 10781 29158 10839 29161
rect 10744 29155 10839 29158
rect 10744 29130 10793 29155
rect 10744 29112 10750 29130
rect 10781 29121 10793 29130
rect 10827 29121 10839 29155
rect 10781 29115 10839 29121
rect 10873 29155 10931 29161
rect 10873 29121 10885 29155
rect 10919 29121 10931 29155
rect 12722 29155 12780 29161
rect 12722 29152 12734 29155
rect 10873 29115 10931 29121
rect 11532 29124 12734 29152
rect 10888 29114 10919 29115
rect 4246 29044 4252 29096
rect 4304 29084 4310 29096
rect 4433 29087 4491 29093
rect 4433 29084 4445 29087
rect 4304 29056 4445 29084
rect 4304 29044 4310 29056
rect 4433 29053 4445 29056
rect 4479 29053 4491 29087
rect 4433 29047 4491 29053
rect 5626 29044 5632 29096
rect 5684 29084 5690 29096
rect 6822 29084 6828 29096
rect 5684 29056 6828 29084
rect 5684 29044 5690 29056
rect 6822 29044 6828 29056
rect 6880 29044 6886 29096
rect 10413 29087 10471 29093
rect 10413 29053 10425 29087
rect 10459 29053 10471 29087
rect 10891 29084 10919 29114
rect 11054 29084 11060 29096
rect 10891 29056 11060 29084
rect 10413 29047 10471 29053
rect 6733 29019 6791 29025
rect 6733 28985 6745 29019
rect 6779 29016 6791 29019
rect 7190 29016 7196 29028
rect 6779 28988 7196 29016
rect 6779 28985 6791 28988
rect 6733 28979 6791 28985
rect 7190 28976 7196 28988
rect 7248 28976 7254 29028
rect 9033 29019 9091 29025
rect 9033 28985 9045 29019
rect 9079 28985 9091 29019
rect 10428 29016 10456 29047
rect 11054 29044 11060 29056
rect 11112 29044 11118 29096
rect 11532 29084 11560 29124
rect 12722 29121 12734 29124
rect 12768 29121 12780 29155
rect 12722 29115 12780 29121
rect 11164 29056 11560 29084
rect 12989 29087 13047 29093
rect 11164 29025 11192 29056
rect 12989 29053 13001 29087
rect 13035 29084 13047 29087
rect 26206 29084 26234 29260
rect 37182 29248 37188 29300
rect 37240 29288 37246 29300
rect 40037 29291 40095 29297
rect 40037 29288 40049 29291
rect 37240 29260 40049 29288
rect 37240 29248 37246 29260
rect 40037 29257 40049 29260
rect 40083 29257 40095 29291
rect 40037 29251 40095 29257
rect 37642 29180 37648 29232
rect 37700 29220 37706 29232
rect 37737 29223 37795 29229
rect 37737 29220 37749 29223
rect 37700 29192 37749 29220
rect 37700 29180 37706 29192
rect 37737 29189 37749 29192
rect 37783 29189 37795 29223
rect 37737 29183 37795 29189
rect 37844 29192 39620 29220
rect 37366 29112 37372 29164
rect 37424 29112 37430 29164
rect 37844 29152 37872 29192
rect 37476 29124 37872 29152
rect 37476 29084 37504 29124
rect 39206 29112 39212 29164
rect 39264 29112 39270 29164
rect 39393 29155 39451 29161
rect 39393 29152 39405 29155
rect 39316 29124 39405 29152
rect 13035 29056 13400 29084
rect 26206 29056 37504 29084
rect 37645 29087 37703 29093
rect 13035 29053 13047 29056
rect 12989 29047 13047 29053
rect 11149 29019 11207 29025
rect 10428 28988 11100 29016
rect 9033 28979 9091 28985
rect 3602 28908 3608 28960
rect 3660 28948 3666 28960
rect 3881 28951 3939 28957
rect 3881 28948 3893 28951
rect 3660 28920 3893 28948
rect 3660 28908 3666 28920
rect 3881 28917 3893 28920
rect 3927 28917 3939 28951
rect 3881 28911 3939 28917
rect 4249 28951 4307 28957
rect 4249 28917 4261 28951
rect 4295 28948 4307 28951
rect 4614 28948 4620 28960
rect 4295 28920 4620 28948
rect 4295 28917 4307 28920
rect 4249 28911 4307 28917
rect 4614 28908 4620 28920
rect 4672 28908 4678 28960
rect 9048 28948 9076 28979
rect 9306 28948 9312 28960
rect 9048 28920 9312 28948
rect 9306 28908 9312 28920
rect 9364 28908 9370 28960
rect 11072 28948 11100 28988
rect 11149 28985 11161 29019
rect 11195 28985 11207 29019
rect 11514 29016 11520 29028
rect 11149 28979 11207 28985
rect 11256 28988 11520 29016
rect 11256 28948 11284 28988
rect 11514 28976 11520 28988
rect 11572 28976 11578 29028
rect 13372 28960 13400 29056
rect 37645 29053 37657 29087
rect 37691 29084 37703 29087
rect 37826 29084 37832 29096
rect 37691 29056 37832 29084
rect 37691 29053 37703 29056
rect 37645 29047 37703 29053
rect 37826 29044 37832 29056
rect 37884 29044 37890 29096
rect 38289 29087 38347 29093
rect 38289 29053 38301 29087
rect 38335 29053 38347 29087
rect 38289 29047 38347 29053
rect 37458 28976 37464 29028
rect 37516 28976 37522 29028
rect 37553 29019 37611 29025
rect 37553 28985 37565 29019
rect 37599 29016 37611 29019
rect 38304 29016 38332 29047
rect 39022 29044 39028 29096
rect 39080 29044 39086 29096
rect 37599 28988 38332 29016
rect 37599 28985 37611 28988
rect 37553 28979 37611 28985
rect 38654 28976 38660 29028
rect 38712 29016 38718 29028
rect 39316 29016 39344 29124
rect 39393 29121 39405 29124
rect 39439 29121 39451 29155
rect 39393 29115 39451 29121
rect 39485 29155 39543 29161
rect 39485 29121 39497 29155
rect 39531 29121 39543 29155
rect 39485 29115 39543 29121
rect 39500 29084 39528 29115
rect 39408 29056 39528 29084
rect 39592 29084 39620 29192
rect 40052 29152 40080 29251
rect 40126 29248 40132 29300
rect 40184 29288 40190 29300
rect 45094 29288 45100 29300
rect 40184 29260 45100 29288
rect 40184 29248 40190 29260
rect 45094 29248 45100 29260
rect 45152 29248 45158 29300
rect 45465 29291 45523 29297
rect 45465 29257 45477 29291
rect 45511 29288 45523 29291
rect 45646 29288 45652 29300
rect 45511 29260 45652 29288
rect 45511 29257 45523 29260
rect 45465 29251 45523 29257
rect 45646 29248 45652 29260
rect 45704 29248 45710 29300
rect 46842 29248 46848 29300
rect 46900 29248 46906 29300
rect 48593 29291 48651 29297
rect 48593 29257 48605 29291
rect 48639 29288 48651 29291
rect 48682 29288 48688 29300
rect 48639 29260 48688 29288
rect 48639 29257 48651 29260
rect 48593 29251 48651 29257
rect 48682 29248 48688 29260
rect 48740 29248 48746 29300
rect 49234 29248 49240 29300
rect 49292 29248 49298 29300
rect 51445 29291 51503 29297
rect 51445 29257 51457 29291
rect 51491 29288 51503 29291
rect 52454 29288 52460 29300
rect 51491 29260 52460 29288
rect 51491 29257 51503 29260
rect 51445 29251 51503 29257
rect 52454 29248 52460 29260
rect 52512 29248 52518 29300
rect 52546 29248 52552 29300
rect 52604 29248 52610 29300
rect 53006 29248 53012 29300
rect 53064 29288 53070 29300
rect 53469 29291 53527 29297
rect 53469 29288 53481 29291
rect 53064 29260 53481 29288
rect 53064 29248 53070 29260
rect 53469 29257 53481 29260
rect 53515 29288 53527 29291
rect 53834 29288 53840 29300
rect 53515 29260 53840 29288
rect 53515 29257 53527 29260
rect 53469 29251 53527 29257
rect 40954 29180 40960 29232
rect 41012 29180 41018 29232
rect 43530 29180 43536 29232
rect 43588 29220 43594 29232
rect 43588 29192 44772 29220
rect 43588 29180 43594 29192
rect 40221 29155 40279 29161
rect 40221 29152 40233 29155
rect 40052 29124 40233 29152
rect 40221 29121 40233 29124
rect 40267 29121 40279 29155
rect 40221 29115 40279 29121
rect 44177 29155 44235 29161
rect 44177 29121 44189 29155
rect 44223 29121 44235 29155
rect 44177 29115 44235 29121
rect 42245 29087 42303 29093
rect 42245 29084 42257 29087
rect 39592 29056 42257 29084
rect 39408 29025 39436 29056
rect 42245 29053 42257 29056
rect 42291 29084 42303 29087
rect 42794 29084 42800 29096
rect 42291 29056 42800 29084
rect 42291 29053 42303 29056
rect 42245 29047 42303 29053
rect 42794 29044 42800 29056
rect 42852 29084 42858 29096
rect 42981 29087 43039 29093
rect 42981 29084 42993 29087
rect 42852 29056 42993 29084
rect 42852 29044 42858 29056
rect 42981 29053 42993 29056
rect 43027 29053 43039 29087
rect 42981 29047 43039 29053
rect 38712 28988 39344 29016
rect 39393 29019 39451 29025
rect 38712 28976 38718 28988
rect 39393 28985 39405 29019
rect 39439 28985 39451 29019
rect 39393 28979 39451 28985
rect 39482 28976 39488 29028
rect 39540 29016 39546 29028
rect 39577 29019 39635 29025
rect 39577 29016 39589 29019
rect 39540 28988 39589 29016
rect 39540 28976 39546 28988
rect 39577 28985 39589 28988
rect 39623 28985 39635 29019
rect 39577 28979 39635 28985
rect 44082 28976 44088 29028
rect 44140 29016 44146 29028
rect 44192 29016 44220 29115
rect 44744 29096 44772 29192
rect 46661 29155 46719 29161
rect 46661 29121 46673 29155
rect 46707 29152 46719 29155
rect 46860 29152 46888 29248
rect 46707 29124 46888 29152
rect 46707 29121 46719 29124
rect 46661 29115 46719 29121
rect 49142 29112 49148 29164
rect 49200 29112 49206 29164
rect 49252 29152 49280 29248
rect 51350 29180 51356 29232
rect 51408 29220 51414 29232
rect 52564 29220 52592 29248
rect 51408 29192 52592 29220
rect 51408 29180 51414 29192
rect 49881 29155 49939 29161
rect 49881 29152 49893 29155
rect 49252 29124 49893 29152
rect 49881 29121 49893 29124
rect 49927 29121 49939 29155
rect 51261 29155 51319 29161
rect 51261 29152 51273 29155
rect 49881 29115 49939 29121
rect 51184 29124 51273 29152
rect 44726 29044 44732 29096
rect 44784 29044 44790 29096
rect 46106 29044 46112 29096
rect 46164 29084 46170 29096
rect 46753 29087 46811 29093
rect 46753 29084 46765 29087
rect 46164 29056 46765 29084
rect 46164 29044 46170 29056
rect 46753 29053 46765 29056
rect 46799 29053 46811 29087
rect 46753 29047 46811 29053
rect 48133 29087 48191 29093
rect 48133 29053 48145 29087
rect 48179 29084 48191 29087
rect 48222 29084 48228 29096
rect 48179 29056 48228 29084
rect 48179 29053 48191 29056
rect 48133 29047 48191 29053
rect 48222 29044 48228 29056
rect 48280 29044 48286 29096
rect 48409 29087 48467 29093
rect 48409 29053 48421 29087
rect 48455 29084 48467 29087
rect 49329 29087 49387 29093
rect 49329 29084 49341 29087
rect 48455 29056 49341 29084
rect 48455 29053 48467 29056
rect 48409 29047 48467 29053
rect 49329 29053 49341 29056
rect 49375 29053 49387 29087
rect 49329 29047 49387 29053
rect 49786 29016 49792 29028
rect 44140 28988 49792 29016
rect 44140 28976 44146 28988
rect 49786 28976 49792 28988
rect 49844 28976 49850 29028
rect 11072 28920 11284 28948
rect 13354 28908 13360 28960
rect 13412 28908 13418 28960
rect 38010 28908 38016 28960
rect 38068 28948 38074 28960
rect 38473 28951 38531 28957
rect 38473 28948 38485 28951
rect 38068 28920 38485 28948
rect 38068 28908 38074 28920
rect 38473 28917 38485 28920
rect 38519 28917 38531 28951
rect 38473 28911 38531 28917
rect 40484 28951 40542 28957
rect 40484 28917 40496 28951
rect 40530 28948 40542 28951
rect 40678 28948 40684 28960
rect 40530 28920 40684 28948
rect 40530 28917 40542 28920
rect 40484 28911 40542 28917
rect 40678 28908 40684 28920
rect 40736 28908 40742 28960
rect 42242 28908 42248 28960
rect 42300 28948 42306 28960
rect 42429 28951 42487 28957
rect 42429 28948 42441 28951
rect 42300 28920 42441 28948
rect 42300 28908 42306 28920
rect 42429 28917 42441 28920
rect 42475 28917 42487 28951
rect 42429 28911 42487 28917
rect 45554 28908 45560 28960
rect 45612 28948 45618 28960
rect 46017 28951 46075 28957
rect 46017 28948 46029 28951
rect 45612 28920 46029 28948
rect 45612 28908 45618 28920
rect 46017 28917 46029 28920
rect 46063 28917 46075 28951
rect 46017 28911 46075 28917
rect 47118 28908 47124 28960
rect 47176 28948 47182 28960
rect 51184 28957 51212 29124
rect 51261 29121 51273 29124
rect 51307 29121 51319 29155
rect 51261 29115 51319 29121
rect 51445 29155 51503 29161
rect 51445 29121 51457 29155
rect 51491 29121 51503 29155
rect 51445 29115 51503 29121
rect 51460 29084 51488 29115
rect 51534 29112 51540 29164
rect 51592 29152 51598 29164
rect 51629 29155 51687 29161
rect 51629 29152 51641 29155
rect 51592 29124 51641 29152
rect 51592 29112 51598 29124
rect 51629 29121 51641 29124
rect 51675 29121 51687 29155
rect 51629 29115 51687 29121
rect 51810 29112 51816 29164
rect 51868 29112 51874 29164
rect 52638 29152 52644 29164
rect 51920 29124 52644 29152
rect 51721 29087 51779 29093
rect 51721 29084 51733 29087
rect 51460 29056 51733 29084
rect 51721 29053 51733 29056
rect 51767 29053 51779 29087
rect 51920 29084 51948 29124
rect 52638 29112 52644 29124
rect 52696 29152 52702 29164
rect 53098 29152 53104 29164
rect 52696 29124 53104 29152
rect 52696 29112 52702 29124
rect 53098 29112 53104 29124
rect 53156 29152 53162 29164
rect 53466 29152 53472 29164
rect 53156 29124 53472 29152
rect 53156 29112 53162 29124
rect 53466 29112 53472 29124
rect 53524 29112 53530 29164
rect 53576 29161 53604 29260
rect 53834 29248 53840 29260
rect 53892 29248 53898 29300
rect 55122 29248 55128 29300
rect 55180 29288 55186 29300
rect 55217 29291 55275 29297
rect 55217 29288 55229 29291
rect 55180 29260 55229 29288
rect 55180 29248 55186 29260
rect 55217 29257 55229 29260
rect 55263 29257 55275 29291
rect 55217 29251 55275 29257
rect 55306 29248 55312 29300
rect 55364 29248 55370 29300
rect 55858 29248 55864 29300
rect 55916 29248 55922 29300
rect 55953 29291 56011 29297
rect 55953 29257 55965 29291
rect 55999 29288 56011 29291
rect 56042 29288 56048 29300
rect 55999 29260 56048 29288
rect 55999 29257 56011 29260
rect 55953 29251 56011 29257
rect 56042 29248 56048 29260
rect 56100 29248 56106 29300
rect 56873 29291 56931 29297
rect 56873 29257 56885 29291
rect 56919 29288 56931 29291
rect 56962 29288 56968 29300
rect 56919 29260 56968 29288
rect 56919 29257 56931 29260
rect 56873 29251 56931 29257
rect 56962 29248 56968 29260
rect 57020 29248 57026 29300
rect 57054 29248 57060 29300
rect 57112 29248 57118 29300
rect 58066 29248 58072 29300
rect 58124 29248 58130 29300
rect 54849 29223 54907 29229
rect 54849 29220 54861 29223
rect 53760 29192 54861 29220
rect 53760 29161 53788 29192
rect 54849 29189 54861 29192
rect 54895 29189 54907 29223
rect 54849 29183 54907 29189
rect 55140 29161 55168 29248
rect 53561 29155 53619 29161
rect 53561 29121 53573 29155
rect 53607 29121 53619 29155
rect 53561 29115 53619 29121
rect 53745 29155 53803 29161
rect 53745 29121 53757 29155
rect 53791 29121 53803 29155
rect 55125 29155 55183 29161
rect 53745 29115 53803 29121
rect 53852 29124 54984 29152
rect 51721 29047 51779 29053
rect 51828 29056 51948 29084
rect 47397 28951 47455 28957
rect 47397 28948 47409 28951
rect 47176 28920 47409 28948
rect 47176 28908 47182 28920
rect 47397 28917 47409 28920
rect 47443 28917 47455 28951
rect 47397 28911 47455 28917
rect 51169 28951 51227 28957
rect 51169 28917 51181 28951
rect 51215 28948 51227 28951
rect 51828 28948 51856 29056
rect 51994 29044 52000 29096
rect 52052 29084 52058 29096
rect 52181 29087 52239 29093
rect 52181 29084 52193 29087
rect 52052 29056 52193 29084
rect 52052 29044 52058 29056
rect 52181 29053 52193 29056
rect 52227 29084 52239 29087
rect 53852 29084 53880 29124
rect 52227 29056 53880 29084
rect 52227 29053 52239 29056
rect 52181 29047 52239 29053
rect 54570 29044 54576 29096
rect 54628 29044 54634 29096
rect 54849 29087 54907 29093
rect 54849 29053 54861 29087
rect 54895 29053 54907 29087
rect 54956 29084 54984 29124
rect 55125 29121 55137 29155
rect 55171 29121 55183 29155
rect 55324 29152 55352 29248
rect 55769 29155 55827 29161
rect 55769 29152 55781 29155
rect 55324 29124 55781 29152
rect 55125 29115 55183 29121
rect 55769 29121 55781 29124
rect 55815 29121 55827 29155
rect 55769 29115 55827 29121
rect 55398 29084 55404 29096
rect 54956 29056 55404 29084
rect 54849 29047 54907 29053
rect 52546 28976 52552 29028
rect 52604 29016 52610 29028
rect 54588 29016 54616 29044
rect 52604 28988 54616 29016
rect 54864 29016 54892 29047
rect 55398 29044 55404 29056
rect 55456 29044 55462 29096
rect 55876 29084 55904 29248
rect 56134 29112 56140 29164
rect 56192 29112 56198 29164
rect 56229 29155 56287 29161
rect 56229 29121 56241 29155
rect 56275 29121 56287 29155
rect 56229 29115 56287 29121
rect 56321 29155 56379 29161
rect 56321 29121 56333 29155
rect 56367 29152 56379 29155
rect 56410 29152 56416 29164
rect 56367 29124 56416 29152
rect 56367 29121 56379 29124
rect 56321 29115 56379 29121
rect 55953 29087 56011 29093
rect 55953 29084 55965 29087
rect 55876 29056 55965 29084
rect 55953 29053 55965 29056
rect 55999 29053 56011 29087
rect 56244 29084 56272 29115
rect 56410 29112 56416 29124
rect 56468 29112 56474 29164
rect 56505 29155 56563 29161
rect 56505 29121 56517 29155
rect 56551 29121 56563 29155
rect 56505 29115 56563 29121
rect 56965 29155 57023 29161
rect 56965 29121 56977 29155
rect 57011 29152 57023 29155
rect 57072 29152 57100 29248
rect 57333 29223 57391 29229
rect 57333 29220 57345 29223
rect 57164 29192 57345 29220
rect 57164 29161 57192 29192
rect 57333 29189 57345 29192
rect 57379 29189 57391 29223
rect 57333 29183 57391 29189
rect 57011 29124 57100 29152
rect 57149 29155 57207 29161
rect 57011 29121 57023 29124
rect 56965 29115 57023 29121
rect 57149 29121 57161 29155
rect 57195 29121 57207 29155
rect 57149 29115 57207 29121
rect 56520 29084 56548 29115
rect 57238 29112 57244 29164
rect 57296 29112 57302 29164
rect 57422 29112 57428 29164
rect 57480 29112 57486 29164
rect 58084 29152 58112 29248
rect 58161 29155 58219 29161
rect 58161 29152 58173 29155
rect 58084 29124 58173 29152
rect 58161 29121 58173 29124
rect 58207 29121 58219 29155
rect 58161 29115 58219 29121
rect 58253 29087 58311 29093
rect 58253 29084 58265 29087
rect 56244 29056 58265 29084
rect 55953 29047 56011 29053
rect 58253 29053 58265 29056
rect 58299 29053 58311 29087
rect 58253 29047 58311 29053
rect 56413 29019 56471 29025
rect 56413 29016 56425 29019
rect 54864 28988 56425 29016
rect 52604 28976 52610 28988
rect 56413 28985 56425 28988
rect 56459 28985 56471 29019
rect 56413 28979 56471 28985
rect 56686 28976 56692 29028
rect 56744 29016 56750 29028
rect 57057 29019 57115 29025
rect 57057 29016 57069 29019
rect 56744 28988 57069 29016
rect 56744 28976 56750 28988
rect 57057 28985 57069 28988
rect 57103 28985 57115 29019
rect 57057 28979 57115 28985
rect 51215 28920 51856 28948
rect 51215 28917 51227 28920
rect 51169 28911 51227 28917
rect 53650 28908 53656 28960
rect 53708 28908 53714 28960
rect 55033 28951 55091 28957
rect 55033 28917 55045 28951
rect 55079 28948 55091 28951
rect 55858 28948 55864 28960
rect 55079 28920 55864 28948
rect 55079 28917 55091 28920
rect 55033 28911 55091 28917
rect 55858 28908 55864 28920
rect 55916 28908 55922 28960
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 2038 28704 2044 28756
rect 2096 28704 2102 28756
rect 3973 28747 4031 28753
rect 3973 28713 3985 28747
rect 4019 28744 4031 28747
rect 4062 28744 4068 28756
rect 4019 28716 4068 28744
rect 4019 28713 4031 28716
rect 3973 28707 4031 28713
rect 4062 28704 4068 28716
rect 4120 28704 4126 28756
rect 4706 28704 4712 28756
rect 4764 28744 4770 28756
rect 4801 28747 4859 28753
rect 4801 28744 4813 28747
rect 4764 28716 4813 28744
rect 4764 28704 4770 28716
rect 4801 28713 4813 28716
rect 4847 28713 4859 28747
rect 4801 28707 4859 28713
rect 4890 28704 4896 28756
rect 4948 28744 4954 28756
rect 5810 28744 5816 28756
rect 4948 28716 5816 28744
rect 4948 28704 4954 28716
rect 5810 28704 5816 28716
rect 5868 28704 5874 28756
rect 5902 28704 5908 28756
rect 5960 28704 5966 28756
rect 6086 28704 6092 28756
rect 6144 28704 6150 28756
rect 6457 28747 6515 28753
rect 6457 28713 6469 28747
rect 6503 28744 6515 28747
rect 6730 28744 6736 28756
rect 6503 28716 6736 28744
rect 6503 28713 6515 28716
rect 6457 28707 6515 28713
rect 6730 28704 6736 28716
rect 6788 28704 6794 28756
rect 6822 28704 6828 28756
rect 6880 28744 6886 28756
rect 7282 28744 7288 28756
rect 6880 28716 7288 28744
rect 6880 28704 6886 28716
rect 7282 28704 7288 28716
rect 7340 28744 7346 28756
rect 9953 28747 10011 28753
rect 7340 28716 7972 28744
rect 7340 28704 7346 28716
rect 2056 28676 2084 28704
rect 4249 28679 4307 28685
rect 4249 28676 4261 28679
rect 2056 28648 4261 28676
rect 4249 28645 4261 28648
rect 4295 28645 4307 28679
rect 4249 28639 4307 28645
rect 6104 28676 6132 28704
rect 6546 28676 6552 28688
rect 6104 28648 6552 28676
rect 3329 28611 3387 28617
rect 3329 28577 3341 28611
rect 3375 28608 3387 28611
rect 4798 28608 4804 28620
rect 3375 28580 4804 28608
rect 3375 28577 3387 28580
rect 3329 28571 3387 28577
rect 4798 28568 4804 28580
rect 4856 28568 4862 28620
rect 5442 28568 5448 28620
rect 5500 28568 5506 28620
rect 3237 28543 3295 28549
rect 3237 28509 3249 28543
rect 3283 28509 3295 28543
rect 3237 28503 3295 28509
rect 3421 28543 3479 28549
rect 3421 28509 3433 28543
rect 3467 28540 3479 28543
rect 3602 28540 3608 28552
rect 3467 28512 3608 28540
rect 3467 28509 3479 28512
rect 3421 28503 3479 28509
rect 3252 28472 3280 28503
rect 3602 28500 3608 28512
rect 3660 28500 3666 28552
rect 3694 28500 3700 28552
rect 3752 28540 3758 28552
rect 3881 28543 3939 28549
rect 3881 28540 3893 28543
rect 3752 28512 3893 28540
rect 3752 28500 3758 28512
rect 3881 28509 3893 28512
rect 3927 28540 3939 28543
rect 4062 28540 4068 28552
rect 3927 28512 4068 28540
rect 3927 28509 3939 28512
rect 3881 28503 3939 28509
rect 4062 28500 4068 28512
rect 4120 28500 4126 28552
rect 4154 28500 4160 28552
rect 4212 28500 4218 28552
rect 4341 28543 4399 28549
rect 4341 28509 4353 28543
rect 4387 28509 4399 28543
rect 4341 28503 4399 28509
rect 4525 28543 4583 28549
rect 4525 28509 4537 28543
rect 4571 28540 4583 28543
rect 4614 28540 4620 28552
rect 4571 28512 4620 28540
rect 4571 28509 4583 28512
rect 4525 28503 4583 28509
rect 3786 28472 3792 28484
rect 3252 28444 3792 28472
rect 3786 28432 3792 28444
rect 3844 28432 3850 28484
rect 4356 28472 4384 28503
rect 4614 28500 4620 28512
rect 4672 28500 4678 28552
rect 5460 28540 5488 28568
rect 4724 28512 5488 28540
rect 5813 28543 5871 28549
rect 4724 28472 4752 28512
rect 5813 28509 5825 28543
rect 5859 28509 5871 28543
rect 5813 28503 5871 28509
rect 5997 28543 6055 28549
rect 5997 28509 6009 28543
rect 6043 28540 6055 28543
rect 6104 28540 6132 28648
rect 6546 28636 6552 28648
rect 6604 28636 6610 28688
rect 7944 28617 7972 28716
rect 9953 28713 9965 28747
rect 9999 28744 10011 28747
rect 10502 28744 10508 28756
rect 9999 28716 10508 28744
rect 9999 28713 10011 28716
rect 9953 28707 10011 28713
rect 10502 28704 10508 28716
rect 10560 28704 10566 28756
rect 10594 28704 10600 28756
rect 10652 28704 10658 28756
rect 11238 28704 11244 28756
rect 11296 28704 11302 28756
rect 11609 28747 11667 28753
rect 11609 28713 11621 28747
rect 11655 28744 11667 28747
rect 11882 28744 11888 28756
rect 11655 28716 11888 28744
rect 11655 28713 11667 28716
rect 11609 28707 11667 28713
rect 11882 28704 11888 28716
rect 11940 28704 11946 28756
rect 36262 28704 36268 28756
rect 36320 28744 36326 28756
rect 36541 28747 36599 28753
rect 36541 28744 36553 28747
rect 36320 28716 36553 28744
rect 36320 28704 36326 28716
rect 36541 28713 36553 28716
rect 36587 28713 36599 28747
rect 36541 28707 36599 28713
rect 9858 28636 9864 28688
rect 9916 28636 9922 28688
rect 7929 28611 7987 28617
rect 7929 28577 7941 28611
rect 7975 28577 7987 28611
rect 9876 28608 9904 28636
rect 9876 28580 10456 28608
rect 7929 28571 7987 28577
rect 6914 28540 6920 28552
rect 6043 28512 6132 28540
rect 6196 28512 6920 28540
rect 6043 28509 6055 28512
rect 5997 28503 6055 28509
rect 4356 28444 4752 28472
rect 4801 28475 4859 28481
rect 4801 28441 4813 28475
rect 4847 28472 4859 28475
rect 4890 28472 4896 28484
rect 4847 28444 4896 28472
rect 4847 28441 4859 28444
rect 4801 28435 4859 28441
rect 4890 28432 4896 28444
rect 4948 28432 4954 28484
rect 4982 28432 4988 28484
rect 5040 28472 5046 28484
rect 5828 28472 5856 28503
rect 6089 28475 6147 28481
rect 6089 28472 6101 28475
rect 5040 28444 6101 28472
rect 5040 28432 5046 28444
rect 6089 28441 6101 28444
rect 6135 28472 6147 28475
rect 6196 28472 6224 28512
rect 6914 28500 6920 28512
rect 6972 28500 6978 28552
rect 7190 28500 7196 28552
rect 7248 28540 7254 28552
rect 7662 28543 7720 28549
rect 7662 28540 7674 28543
rect 7248 28512 7674 28540
rect 7248 28500 7254 28512
rect 7662 28509 7674 28512
rect 7708 28509 7720 28543
rect 9861 28543 9919 28549
rect 9861 28540 9873 28543
rect 7662 28503 7720 28509
rect 9324 28512 9873 28540
rect 6135 28444 6224 28472
rect 6273 28475 6331 28481
rect 6135 28441 6147 28444
rect 6089 28435 6147 28441
rect 6273 28441 6285 28475
rect 6319 28472 6331 28475
rect 8386 28472 8392 28484
rect 6319 28444 8392 28472
rect 6319 28441 6331 28444
rect 6273 28435 6331 28441
rect 8386 28432 8392 28444
rect 8444 28432 8450 28484
rect 9324 28416 9352 28512
rect 9861 28509 9873 28512
rect 9907 28509 9919 28543
rect 9861 28503 9919 28509
rect 9950 28500 9956 28552
rect 10008 28540 10014 28552
rect 10428 28549 10456 28580
rect 12526 28568 12532 28620
rect 12584 28608 12590 28620
rect 36556 28608 36584 28707
rect 37458 28704 37464 28756
rect 37516 28744 37522 28756
rect 38378 28744 38384 28756
rect 37516 28716 38384 28744
rect 37516 28704 37522 28716
rect 38378 28704 38384 28716
rect 38436 28704 38442 28756
rect 38657 28747 38715 28753
rect 38657 28713 38669 28747
rect 38703 28744 38715 28747
rect 39022 28744 39028 28756
rect 38703 28716 39028 28744
rect 38703 28713 38715 28716
rect 38657 28707 38715 28713
rect 39022 28704 39028 28716
rect 39080 28704 39086 28756
rect 40678 28704 40684 28756
rect 40736 28744 40742 28756
rect 40773 28747 40831 28753
rect 40773 28744 40785 28747
rect 40736 28716 40785 28744
rect 40736 28704 40742 28716
rect 40773 28713 40785 28716
rect 40819 28713 40831 28747
rect 40773 28707 40831 28713
rect 42794 28704 42800 28756
rect 42852 28704 42858 28756
rect 44634 28704 44640 28756
rect 44692 28744 44698 28756
rect 44729 28747 44787 28753
rect 44729 28744 44741 28747
rect 44692 28716 44741 28744
rect 44692 28704 44698 28716
rect 44729 28713 44741 28716
rect 44775 28713 44787 28747
rect 44729 28707 44787 28713
rect 45557 28747 45615 28753
rect 45557 28713 45569 28747
rect 45603 28744 45615 28747
rect 46106 28744 46112 28756
rect 45603 28716 46112 28744
rect 45603 28713 45615 28716
rect 45557 28707 45615 28713
rect 46106 28704 46112 28716
rect 46164 28704 46170 28756
rect 48130 28704 48136 28756
rect 48188 28704 48194 28756
rect 48314 28704 48320 28756
rect 48372 28744 48378 28756
rect 48593 28747 48651 28753
rect 48593 28744 48605 28747
rect 48372 28716 48605 28744
rect 48372 28704 48378 28716
rect 48593 28713 48605 28716
rect 48639 28713 48651 28747
rect 48593 28707 48651 28713
rect 48869 28747 48927 28753
rect 48869 28713 48881 28747
rect 48915 28713 48927 28747
rect 48869 28707 48927 28713
rect 38010 28636 38016 28688
rect 38068 28636 38074 28688
rect 38396 28676 38424 28704
rect 39393 28679 39451 28685
rect 39393 28676 39405 28679
rect 38396 28648 39405 28676
rect 39393 28645 39405 28648
rect 39439 28645 39451 28679
rect 41785 28679 41843 28685
rect 41785 28676 41797 28679
rect 39393 28639 39451 28645
rect 41708 28648 41797 28676
rect 36725 28611 36783 28617
rect 36725 28608 36737 28611
rect 12584 28580 12940 28608
rect 36556 28580 36737 28608
rect 12584 28568 12590 28580
rect 10045 28543 10103 28549
rect 10045 28540 10057 28543
rect 10008 28512 10057 28540
rect 10008 28500 10014 28512
rect 10045 28509 10057 28512
rect 10091 28509 10103 28543
rect 10045 28503 10103 28509
rect 10413 28543 10471 28549
rect 10413 28509 10425 28543
rect 10459 28509 10471 28543
rect 10413 28503 10471 28509
rect 10060 28472 10088 28503
rect 11054 28500 11060 28552
rect 11112 28540 11118 28552
rect 11241 28543 11299 28549
rect 11241 28540 11253 28543
rect 11112 28512 11253 28540
rect 11112 28500 11118 28512
rect 11241 28509 11253 28512
rect 11287 28509 11299 28543
rect 11241 28503 11299 28509
rect 11330 28500 11336 28552
rect 11388 28500 11394 28552
rect 12912 28549 12940 28580
rect 36725 28577 36737 28580
rect 36771 28577 36783 28611
rect 36725 28571 36783 28577
rect 37001 28611 37059 28617
rect 37001 28577 37013 28611
rect 37047 28608 37059 28611
rect 38028 28608 38056 28636
rect 41708 28617 41736 28648
rect 41785 28645 41797 28648
rect 41831 28645 41843 28679
rect 45186 28676 45192 28688
rect 41785 28639 41843 28645
rect 44468 28648 45192 28676
rect 37047 28580 38056 28608
rect 41693 28611 41751 28617
rect 37047 28577 37059 28580
rect 37001 28571 37059 28577
rect 41693 28577 41705 28611
rect 41739 28577 41751 28611
rect 41693 28571 41751 28577
rect 42242 28568 42248 28620
rect 42300 28568 42306 28620
rect 42429 28611 42487 28617
rect 42429 28577 42441 28611
rect 42475 28608 42487 28611
rect 42794 28608 42800 28620
rect 42475 28580 42800 28608
rect 42475 28577 42487 28580
rect 42429 28571 42487 28577
rect 42794 28568 42800 28580
rect 42852 28568 42858 28620
rect 12897 28543 12955 28549
rect 12897 28509 12909 28543
rect 12943 28540 12955 28543
rect 12986 28540 12992 28552
rect 12943 28512 12992 28540
rect 12943 28509 12955 28512
rect 12897 28503 12955 28509
rect 12986 28500 12992 28512
rect 13044 28500 13050 28552
rect 38562 28500 38568 28552
rect 38620 28500 38626 28552
rect 38749 28543 38807 28549
rect 38749 28509 38761 28543
rect 38795 28540 38807 28543
rect 40957 28543 41015 28549
rect 38795 28512 39344 28540
rect 38795 28509 38807 28512
rect 38749 28503 38807 28509
rect 10229 28475 10287 28481
rect 10229 28472 10241 28475
rect 10060 28444 10241 28472
rect 10229 28441 10241 28444
rect 10275 28441 10287 28475
rect 10229 28435 10287 28441
rect 37458 28432 37464 28484
rect 37516 28432 37522 28484
rect 38654 28472 38660 28484
rect 38304 28444 38660 28472
rect 4617 28407 4675 28413
rect 4617 28373 4629 28407
rect 4663 28404 4675 28407
rect 4706 28404 4712 28416
rect 4663 28376 4712 28404
rect 4663 28373 4675 28376
rect 4617 28367 4675 28373
rect 4706 28364 4712 28376
rect 4764 28364 4770 28416
rect 5169 28407 5227 28413
rect 5169 28373 5181 28407
rect 5215 28404 5227 28407
rect 5350 28404 5356 28416
rect 5215 28376 5356 28404
rect 5215 28373 5227 28376
rect 5169 28367 5227 28373
rect 5350 28364 5356 28376
rect 5408 28364 5414 28416
rect 5534 28364 5540 28416
rect 5592 28404 5598 28416
rect 9122 28404 9128 28416
rect 5592 28376 9128 28404
rect 5592 28364 5598 28376
rect 9122 28364 9128 28376
rect 9180 28364 9186 28416
rect 9306 28364 9312 28416
rect 9364 28364 9370 28416
rect 12989 28407 13047 28413
rect 12989 28373 13001 28407
rect 13035 28404 13047 28407
rect 13354 28404 13360 28416
rect 13035 28376 13360 28404
rect 13035 28373 13047 28376
rect 12989 28367 13047 28373
rect 13354 28364 13360 28376
rect 13412 28404 13418 28416
rect 38304 28404 38332 28444
rect 38654 28432 38660 28444
rect 38712 28472 38718 28484
rect 39025 28475 39083 28481
rect 39025 28472 39037 28475
rect 38712 28444 39037 28472
rect 38712 28432 38718 28444
rect 39025 28441 39037 28444
rect 39071 28441 39083 28475
rect 39025 28435 39083 28441
rect 39316 28416 39344 28512
rect 40957 28509 40969 28543
rect 41003 28540 41015 28543
rect 41049 28543 41107 28549
rect 41049 28540 41061 28543
rect 41003 28512 41061 28540
rect 41003 28509 41015 28512
rect 40957 28503 41015 28509
rect 41049 28509 41061 28512
rect 41095 28509 41107 28543
rect 41049 28503 41107 28509
rect 42518 28500 42524 28552
rect 42576 28540 42582 28552
rect 42981 28543 43039 28549
rect 42981 28540 42993 28543
rect 42576 28512 42993 28540
rect 42576 28500 42582 28512
rect 42981 28509 42993 28512
rect 43027 28509 43039 28543
rect 44468 28540 44496 28648
rect 45186 28636 45192 28648
rect 45244 28676 45250 28688
rect 48148 28676 48176 28704
rect 48884 28676 48912 28707
rect 49142 28704 49148 28756
rect 49200 28744 49206 28756
rect 49237 28747 49295 28753
rect 49237 28744 49249 28747
rect 49200 28716 49249 28744
rect 49200 28704 49206 28716
rect 49237 28713 49249 28716
rect 49283 28713 49295 28747
rect 50154 28744 50160 28756
rect 49237 28707 49295 28713
rect 49620 28716 50160 28744
rect 49513 28679 49571 28685
rect 49513 28676 49525 28679
rect 45244 28648 45784 28676
rect 48148 28648 49525 28676
rect 45244 28636 45250 28648
rect 45646 28568 45652 28620
rect 45704 28568 45710 28620
rect 45756 28608 45784 28648
rect 49513 28645 49525 28648
rect 49559 28645 49571 28679
rect 49513 28639 49571 28645
rect 46566 28608 46572 28620
rect 45756 28580 46572 28608
rect 46566 28568 46572 28580
rect 46624 28568 46630 28620
rect 47397 28611 47455 28617
rect 47397 28577 47409 28611
rect 47443 28608 47455 28611
rect 47949 28611 48007 28617
rect 47949 28608 47961 28611
rect 47443 28580 47961 28608
rect 47443 28577 47455 28580
rect 47397 28571 47455 28577
rect 47949 28577 47961 28580
rect 47995 28577 48007 28611
rect 47949 28571 48007 28577
rect 48314 28568 48320 28620
rect 48372 28568 48378 28620
rect 44390 28512 44496 28540
rect 45097 28543 45155 28549
rect 42981 28503 43039 28509
rect 45097 28509 45109 28543
rect 45143 28509 45155 28543
rect 45097 28503 45155 28509
rect 43254 28432 43260 28484
rect 43312 28432 43318 28484
rect 45112 28472 45140 28503
rect 45186 28500 45192 28552
rect 45244 28500 45250 28552
rect 45373 28543 45431 28549
rect 45373 28509 45385 28543
rect 45419 28540 45431 28543
rect 45554 28540 45560 28552
rect 45419 28512 45560 28540
rect 45419 28509 45431 28512
rect 45373 28503 45431 28509
rect 45554 28500 45560 28512
rect 45612 28500 45618 28552
rect 48332 28540 48360 28568
rect 49620 28549 49648 28716
rect 50154 28704 50160 28716
rect 50212 28704 50218 28756
rect 51534 28704 51540 28756
rect 51592 28704 51598 28756
rect 51810 28704 51816 28756
rect 51868 28744 51874 28756
rect 51997 28747 52055 28753
rect 51997 28744 52009 28747
rect 51868 28716 52009 28744
rect 51868 28704 51874 28716
rect 51997 28713 52009 28716
rect 52043 28713 52055 28747
rect 51997 28707 52055 28713
rect 57146 28704 57152 28756
rect 57204 28704 57210 28756
rect 57422 28704 57428 28756
rect 57480 28744 57486 28756
rect 57517 28747 57575 28753
rect 57517 28744 57529 28747
rect 57480 28716 57529 28744
rect 57480 28704 57486 28716
rect 57517 28713 57529 28716
rect 57563 28713 57575 28747
rect 57517 28707 57575 28713
rect 49697 28679 49755 28685
rect 49697 28645 49709 28679
rect 49743 28676 49755 28679
rect 49878 28676 49884 28688
rect 49743 28648 49884 28676
rect 49743 28645 49755 28648
rect 49697 28639 49755 28645
rect 49878 28636 49884 28648
rect 49936 28636 49942 28688
rect 55214 28676 55220 28688
rect 51276 28648 55220 28676
rect 50157 28611 50215 28617
rect 50157 28577 50169 28611
rect 50203 28608 50215 28611
rect 50246 28608 50252 28620
rect 50203 28580 50252 28608
rect 50203 28577 50215 28580
rect 50157 28571 50215 28577
rect 50246 28568 50252 28580
rect 50304 28568 50310 28620
rect 49145 28543 49203 28549
rect 49145 28540 49157 28543
rect 48332 28512 49157 28540
rect 49145 28509 49157 28512
rect 49191 28509 49203 28543
rect 49145 28503 49203 28509
rect 49605 28543 49663 28549
rect 49605 28509 49617 28543
rect 49651 28509 49663 28543
rect 49605 28503 49663 28509
rect 49973 28543 50031 28549
rect 49973 28509 49985 28543
rect 50019 28540 50031 28543
rect 50614 28540 50620 28552
rect 50019 28512 50620 28540
rect 50019 28509 50031 28512
rect 49973 28503 50031 28509
rect 50614 28500 50620 28512
rect 50672 28500 50678 28552
rect 51276 28540 51304 28648
rect 55214 28636 55220 28648
rect 55272 28636 55278 28688
rect 52273 28611 52331 28617
rect 52273 28608 52285 28611
rect 51644 28580 52285 28608
rect 51644 28549 51672 28580
rect 52273 28577 52285 28580
rect 52319 28577 52331 28611
rect 52273 28571 52331 28577
rect 57425 28611 57483 28617
rect 57425 28577 57437 28611
rect 57471 28608 57483 28611
rect 57977 28611 58035 28617
rect 57977 28608 57989 28611
rect 57471 28580 57989 28608
rect 57471 28577 57483 28580
rect 57425 28571 57483 28577
rect 57977 28577 57989 28580
rect 58023 28577 58035 28611
rect 57977 28571 58035 28577
rect 51092 28512 51304 28540
rect 51537 28543 51595 28549
rect 45925 28475 45983 28481
rect 45925 28472 45937 28475
rect 45112 28444 45937 28472
rect 45925 28441 45937 28444
rect 45971 28441 45983 28475
rect 45925 28435 45983 28441
rect 13412 28376 38332 28404
rect 13412 28364 13418 28376
rect 38470 28364 38476 28416
rect 38528 28364 38534 28416
rect 39298 28364 39304 28416
rect 39356 28364 39362 28416
rect 42153 28407 42211 28413
rect 42153 28373 42165 28407
rect 42199 28404 42211 28407
rect 43070 28404 43076 28416
rect 42199 28376 43076 28404
rect 42199 28373 42211 28376
rect 42153 28367 42211 28373
rect 43070 28364 43076 28376
rect 43128 28364 43134 28416
rect 45940 28404 45968 28435
rect 46566 28432 46572 28484
rect 46624 28432 46630 28484
rect 48038 28432 48044 28484
rect 48096 28472 48102 28484
rect 48853 28475 48911 28481
rect 48096 28444 48728 28472
rect 48096 28432 48102 28444
rect 48222 28404 48228 28416
rect 45940 28376 48228 28404
rect 48222 28364 48228 28376
rect 48280 28364 48286 28416
rect 48700 28413 48728 28444
rect 48853 28441 48865 28475
rect 48899 28472 48911 28475
rect 49053 28475 49111 28481
rect 48899 28444 49004 28472
rect 48899 28441 48911 28444
rect 48853 28435 48911 28441
rect 48685 28407 48743 28413
rect 48685 28373 48697 28407
rect 48731 28373 48743 28407
rect 48976 28404 49004 28444
rect 49053 28441 49065 28475
rect 49099 28472 49111 28475
rect 49099 28444 49280 28472
rect 49099 28441 49111 28444
rect 49053 28435 49111 28441
rect 49142 28404 49148 28416
rect 48976 28376 49148 28404
rect 48685 28367 48743 28373
rect 49142 28364 49148 28376
rect 49200 28364 49206 28416
rect 49252 28404 49280 28444
rect 49694 28432 49700 28484
rect 49752 28432 49758 28484
rect 49881 28475 49939 28481
rect 49881 28441 49893 28475
rect 49927 28472 49939 28475
rect 50706 28472 50712 28484
rect 49927 28444 50712 28472
rect 49927 28441 49939 28444
rect 49881 28435 49939 28441
rect 50706 28432 50712 28444
rect 50764 28432 50770 28484
rect 49970 28404 49976 28416
rect 49252 28376 49976 28404
rect 49970 28364 49976 28376
rect 50028 28364 50034 28416
rect 50062 28364 50068 28416
rect 50120 28404 50126 28416
rect 50433 28407 50491 28413
rect 50433 28404 50445 28407
rect 50120 28376 50445 28404
rect 50120 28364 50126 28376
rect 50433 28373 50445 28376
rect 50479 28373 50491 28407
rect 50433 28367 50491 28373
rect 50525 28407 50583 28413
rect 50525 28373 50537 28407
rect 50571 28404 50583 28407
rect 51092 28404 51120 28512
rect 51537 28509 51549 28543
rect 51583 28509 51595 28543
rect 51537 28503 51595 28509
rect 51629 28543 51687 28549
rect 51629 28509 51641 28543
rect 51675 28509 51687 28543
rect 51629 28503 51687 28509
rect 51552 28416 51580 28503
rect 51718 28500 51724 28552
rect 51776 28540 51782 28552
rect 51813 28543 51871 28549
rect 51813 28540 51825 28543
rect 51776 28512 51825 28540
rect 51776 28500 51782 28512
rect 51813 28509 51825 28512
rect 51859 28509 51871 28543
rect 51813 28503 51871 28509
rect 51905 28543 51963 28549
rect 51905 28509 51917 28543
rect 51951 28540 51963 28543
rect 51994 28540 52000 28552
rect 51951 28512 52000 28540
rect 51951 28509 51963 28512
rect 51905 28503 51963 28509
rect 50571 28376 51120 28404
rect 50571 28373 50583 28376
rect 50525 28367 50583 28373
rect 51534 28364 51540 28416
rect 51592 28364 51598 28416
rect 51718 28364 51724 28416
rect 51776 28404 51782 28416
rect 51920 28404 51948 28503
rect 51994 28500 52000 28512
rect 52052 28500 52058 28552
rect 52089 28543 52147 28549
rect 52089 28509 52101 28543
rect 52135 28540 52147 28543
rect 52178 28540 52184 28552
rect 52135 28512 52184 28540
rect 52135 28509 52147 28512
rect 52089 28503 52147 28509
rect 52178 28500 52184 28512
rect 52236 28500 52242 28552
rect 52365 28543 52423 28549
rect 52365 28509 52377 28543
rect 52411 28540 52423 28543
rect 52546 28540 52552 28552
rect 52411 28512 52552 28540
rect 52411 28509 52423 28512
rect 52365 28503 52423 28509
rect 52546 28500 52552 28512
rect 52604 28500 52610 28552
rect 53193 28543 53251 28549
rect 53193 28509 53205 28543
rect 53239 28509 53251 28543
rect 53193 28503 53251 28509
rect 53377 28543 53435 28549
rect 53377 28509 53389 28543
rect 53423 28540 53435 28543
rect 53650 28540 53656 28552
rect 53423 28512 53656 28540
rect 53423 28509 53435 28512
rect 53377 28503 53435 28509
rect 53208 28416 53236 28503
rect 53650 28500 53656 28512
rect 53708 28500 53714 28552
rect 55858 28500 55864 28552
rect 55916 28540 55922 28552
rect 56410 28540 56416 28552
rect 55916 28512 56416 28540
rect 55916 28500 55922 28512
rect 56410 28500 56416 28512
rect 56468 28540 56474 28552
rect 57606 28540 57612 28552
rect 56468 28512 57612 28540
rect 56468 28500 56474 28512
rect 57606 28500 57612 28512
rect 57664 28500 57670 28552
rect 57698 28500 57704 28552
rect 57756 28500 57762 28552
rect 57790 28500 57796 28552
rect 57848 28540 57854 28552
rect 57885 28543 57943 28549
rect 57885 28540 57897 28543
rect 57848 28512 57897 28540
rect 57848 28500 57854 28512
rect 57885 28509 57897 28512
rect 57931 28509 57943 28543
rect 57885 28503 57943 28509
rect 58069 28543 58127 28549
rect 58069 28509 58081 28543
rect 58115 28509 58127 28543
rect 58069 28503 58127 28509
rect 58084 28472 58112 28503
rect 58342 28500 58348 28552
rect 58400 28500 58406 28552
rect 58253 28475 58311 28481
rect 58253 28472 58265 28475
rect 56612 28444 58265 28472
rect 56612 28416 56640 28444
rect 58253 28441 58265 28444
rect 58299 28441 58311 28475
rect 58253 28435 58311 28441
rect 51776 28376 51948 28404
rect 51776 28364 51782 28376
rect 53190 28364 53196 28416
rect 53248 28364 53254 28416
rect 53282 28364 53288 28416
rect 53340 28364 53346 28416
rect 56594 28364 56600 28416
rect 56652 28364 56658 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 3970 28160 3976 28212
rect 4028 28160 4034 28212
rect 4062 28160 4068 28212
rect 4120 28200 4126 28212
rect 4893 28203 4951 28209
rect 4893 28200 4905 28203
rect 4120 28172 4905 28200
rect 4120 28160 4126 28172
rect 4893 28169 4905 28172
rect 4939 28200 4951 28203
rect 6362 28200 6368 28212
rect 4939 28172 6368 28200
rect 4939 28169 4951 28172
rect 4893 28163 4951 28169
rect 6362 28160 6368 28172
rect 6420 28160 6426 28212
rect 7098 28160 7104 28212
rect 7156 28200 7162 28212
rect 8021 28203 8079 28209
rect 8021 28200 8033 28203
rect 7156 28172 8033 28200
rect 7156 28160 7162 28172
rect 8021 28169 8033 28172
rect 8067 28169 8079 28203
rect 8021 28163 8079 28169
rect 8220 28172 8708 28200
rect 4080 28104 4660 28132
rect 2682 28024 2688 28076
rect 2740 28024 2746 28076
rect 4080 28073 4108 28104
rect 4632 28073 4660 28104
rect 3881 28067 3939 28073
rect 3881 28033 3893 28067
rect 3927 28033 3939 28067
rect 3881 28027 3939 28033
rect 4065 28067 4123 28073
rect 4065 28033 4077 28067
rect 4111 28033 4123 28067
rect 4065 28027 4123 28033
rect 4433 28067 4491 28073
rect 4433 28033 4445 28067
rect 4479 28033 4491 28067
rect 4433 28027 4491 28033
rect 4617 28067 4675 28073
rect 4617 28033 4629 28067
rect 4663 28064 4675 28067
rect 4798 28064 4804 28076
rect 4663 28036 4804 28064
rect 4663 28033 4675 28036
rect 4617 28027 4675 28033
rect 1578 27956 1584 28008
rect 1636 27956 1642 28008
rect 3418 27956 3424 28008
rect 3476 27956 3482 28008
rect 3896 27928 3924 28027
rect 4448 27996 4476 28027
rect 4798 28024 4804 28036
rect 4856 28024 4862 28076
rect 8220 28073 8248 28172
rect 8386 28092 8392 28144
rect 8444 28132 8450 28144
rect 8573 28135 8631 28141
rect 8573 28132 8585 28135
rect 8444 28104 8585 28132
rect 8444 28092 8450 28104
rect 8573 28101 8585 28104
rect 8619 28101 8631 28135
rect 8680 28132 8708 28172
rect 8754 28160 8760 28212
rect 8812 28200 8818 28212
rect 9033 28203 9091 28209
rect 9033 28200 9045 28203
rect 8812 28172 9045 28200
rect 8812 28160 8818 28172
rect 9033 28169 9045 28172
rect 9079 28169 9091 28203
rect 9033 28163 9091 28169
rect 9122 28160 9128 28212
rect 9180 28160 9186 28212
rect 10226 28160 10232 28212
rect 10284 28200 10290 28212
rect 10781 28203 10839 28209
rect 10781 28200 10793 28203
rect 10284 28172 10793 28200
rect 10284 28160 10290 28172
rect 10781 28169 10793 28172
rect 10827 28169 10839 28203
rect 10781 28163 10839 28169
rect 38470 28160 38476 28212
rect 38528 28160 38534 28212
rect 38562 28160 38568 28212
rect 38620 28200 38626 28212
rect 39117 28203 39175 28209
rect 39117 28200 39129 28203
rect 38620 28172 39129 28200
rect 38620 28160 38626 28172
rect 39117 28169 39129 28172
rect 39163 28169 39175 28203
rect 39117 28163 39175 28169
rect 39206 28160 39212 28212
rect 39264 28160 39270 28212
rect 40034 28160 40040 28212
rect 40092 28160 40098 28212
rect 41233 28203 41291 28209
rect 41233 28200 41245 28203
rect 40604 28172 41245 28200
rect 11330 28132 11336 28144
rect 8680 28104 8892 28132
rect 8573 28095 8631 28101
rect 8205 28067 8263 28073
rect 8205 28033 8217 28067
rect 8251 28033 8263 28067
rect 8205 28027 8263 28033
rect 8478 28024 8484 28076
rect 8536 28024 8542 28076
rect 8864 28073 8892 28104
rect 9324 28104 11336 28132
rect 9324 28073 9352 28104
rect 11330 28092 11336 28104
rect 11388 28092 11394 28144
rect 8849 28067 8907 28073
rect 8849 28033 8861 28067
rect 8895 28064 8907 28067
rect 9309 28067 9367 28073
rect 9309 28064 9321 28067
rect 8895 28036 9321 28064
rect 8895 28033 8907 28036
rect 8849 28027 8907 28033
rect 9309 28033 9321 28036
rect 9355 28033 9367 28067
rect 9309 28027 9367 28033
rect 9585 28067 9643 28073
rect 9585 28033 9597 28067
rect 9631 28064 9643 28067
rect 9858 28064 9864 28076
rect 9631 28036 9864 28064
rect 9631 28033 9643 28036
rect 9585 28027 9643 28033
rect 9858 28024 9864 28036
rect 9916 28024 9922 28076
rect 12621 28067 12679 28073
rect 12621 28033 12633 28067
rect 12667 28064 12679 28067
rect 13078 28064 13084 28076
rect 12667 28036 13084 28064
rect 12667 28033 12679 28036
rect 12621 28027 12679 28033
rect 13078 28024 13084 28036
rect 13136 28064 13142 28076
rect 13136 28036 13492 28064
rect 13136 28024 13142 28036
rect 4982 27996 4988 28008
rect 4448 27968 4988 27996
rect 4982 27956 4988 27968
rect 5040 27956 5046 28008
rect 8389 27999 8447 28005
rect 8389 27965 8401 27999
rect 8435 27965 8447 27999
rect 8662 27996 8668 28008
rect 8389 27959 8447 27965
rect 8588 27968 8668 27996
rect 4154 27928 4160 27940
rect 3896 27900 4160 27928
rect 4154 27888 4160 27900
rect 4212 27928 4218 27940
rect 8404 27928 8432 27959
rect 8588 27928 8616 27968
rect 8662 27956 8668 27968
rect 8720 27956 8726 28008
rect 8938 27956 8944 28008
rect 8996 27996 9002 28008
rect 9401 27999 9459 28005
rect 9401 27996 9413 27999
rect 8996 27968 9413 27996
rect 8996 27956 9002 27968
rect 9401 27965 9413 27968
rect 9447 27996 9459 27999
rect 10134 27996 10140 28008
rect 9447 27968 10140 27996
rect 9447 27965 9459 27968
rect 9401 27959 9459 27965
rect 10134 27956 10140 27968
rect 10192 27996 10198 28008
rect 11054 27996 11060 28008
rect 10192 27968 11060 27996
rect 10192 27956 10198 27968
rect 11054 27956 11060 27968
rect 11112 27956 11118 28008
rect 12894 27956 12900 28008
rect 12952 27956 12958 28008
rect 13464 27937 13492 28036
rect 38102 28024 38108 28076
rect 38160 28024 38166 28076
rect 38488 28073 38516 28160
rect 39025 28135 39083 28141
rect 39025 28101 39037 28135
rect 39071 28132 39083 28135
rect 39224 28132 39252 28160
rect 39071 28104 39252 28132
rect 40052 28132 40080 28160
rect 40604 28141 40632 28172
rect 41233 28169 41245 28172
rect 41279 28169 41291 28203
rect 41233 28163 41291 28169
rect 43254 28160 43260 28212
rect 43312 28200 43318 28212
rect 43349 28203 43407 28209
rect 43349 28200 43361 28203
rect 43312 28172 43361 28200
rect 43312 28160 43318 28172
rect 43349 28169 43361 28172
rect 43395 28169 43407 28203
rect 43622 28200 43628 28212
rect 43349 28163 43407 28169
rect 43456 28172 43628 28200
rect 40589 28135 40647 28141
rect 40589 28132 40601 28135
rect 40052 28104 40172 28132
rect 39071 28101 39083 28104
rect 39025 28095 39083 28101
rect 38289 28067 38347 28073
rect 38289 28033 38301 28067
rect 38335 28033 38347 28067
rect 38289 28027 38347 28033
rect 38473 28067 38531 28073
rect 38473 28033 38485 28067
rect 38519 28033 38531 28067
rect 39853 28067 39911 28073
rect 39853 28064 39865 28067
rect 38473 28027 38531 28033
rect 38580 28036 39865 28064
rect 38304 27996 38332 28027
rect 38580 27996 38608 28036
rect 39853 28033 39865 28036
rect 39899 28033 39911 28067
rect 39853 28027 39911 28033
rect 40034 28024 40040 28076
rect 40092 28024 40098 28076
rect 40144 28073 40172 28104
rect 40236 28104 40601 28132
rect 40236 28076 40264 28104
rect 40589 28101 40601 28104
rect 40635 28101 40647 28135
rect 43456 28132 43484 28172
rect 43622 28160 43628 28172
rect 43680 28160 43686 28212
rect 44634 28160 44640 28212
rect 44692 28160 44698 28212
rect 45186 28160 45192 28212
rect 45244 28200 45250 28212
rect 45281 28203 45339 28209
rect 45281 28200 45293 28203
rect 45244 28172 45293 28200
rect 45244 28160 45250 28172
rect 45281 28169 45293 28172
rect 45327 28169 45339 28203
rect 45281 28163 45339 28169
rect 49050 28160 49056 28212
rect 49108 28160 49114 28212
rect 49694 28160 49700 28212
rect 49752 28160 49758 28212
rect 50154 28160 50160 28212
rect 50212 28160 50218 28212
rect 53834 28160 53840 28212
rect 53892 28200 53898 28212
rect 55677 28203 55735 28209
rect 55677 28200 55689 28203
rect 53892 28172 55689 28200
rect 53892 28160 53898 28172
rect 55677 28169 55689 28172
rect 55723 28169 55735 28203
rect 55677 28163 55735 28169
rect 57698 28160 57704 28212
rect 57756 28200 57762 28212
rect 57885 28203 57943 28209
rect 57885 28200 57897 28203
rect 57756 28172 57897 28200
rect 57756 28160 57762 28172
rect 57885 28169 57897 28172
rect 57931 28169 57943 28203
rect 57885 28163 57943 28169
rect 58802 28160 58808 28212
rect 58860 28160 58866 28212
rect 44652 28132 44680 28160
rect 40589 28095 40647 28101
rect 41156 28104 42196 28132
rect 40129 28067 40187 28073
rect 40129 28033 40141 28067
rect 40175 28033 40187 28067
rect 40129 28027 40187 28033
rect 38304 27968 38608 27996
rect 39666 27956 39672 28008
rect 39724 27956 39730 28008
rect 40144 27996 40172 28027
rect 40218 28024 40224 28076
rect 40276 28024 40282 28076
rect 40402 28024 40408 28076
rect 40460 28024 40466 28076
rect 40678 28024 40684 28076
rect 40736 28064 40742 28076
rect 41156 28073 41184 28104
rect 40773 28067 40831 28073
rect 40773 28064 40785 28067
rect 40736 28036 40785 28064
rect 40736 28024 40742 28036
rect 40773 28033 40785 28036
rect 40819 28033 40831 28067
rect 40773 28027 40831 28033
rect 40865 28067 40923 28073
rect 40865 28033 40877 28067
rect 40911 28064 40923 28067
rect 41141 28067 41199 28073
rect 41141 28064 41153 28067
rect 40911 28036 41153 28064
rect 40911 28033 40923 28036
rect 40865 28027 40923 28033
rect 41141 28033 41153 28036
rect 41187 28033 41199 28067
rect 41141 28027 41199 28033
rect 41322 28024 41328 28076
rect 41380 28024 41386 28076
rect 41966 28024 41972 28076
rect 42024 28024 42030 28076
rect 40310 27996 40316 28008
rect 40144 27968 40316 27996
rect 40310 27956 40316 27968
rect 40368 27956 40374 28008
rect 41877 27999 41935 28005
rect 41877 27996 41889 27999
rect 41386 27968 41889 27996
rect 4212 27900 5396 27928
rect 8404 27900 8616 27928
rect 13449 27931 13507 27937
rect 4212 27888 4218 27900
rect 5368 27872 5396 27900
rect 13449 27897 13461 27931
rect 13495 27928 13507 27931
rect 41386 27928 41414 27968
rect 41877 27965 41889 27968
rect 41923 27965 41935 27999
rect 41877 27959 41935 27965
rect 13495 27900 41414 27928
rect 13495 27897 13507 27900
rect 13449 27891 13507 27897
rect 2774 27820 2780 27872
rect 2832 27860 2838 27872
rect 2869 27863 2927 27869
rect 2869 27860 2881 27863
rect 2832 27832 2881 27860
rect 2832 27820 2838 27832
rect 2869 27829 2881 27832
rect 2915 27829 2927 27863
rect 2869 27823 2927 27829
rect 4525 27863 4583 27869
rect 4525 27829 4537 27863
rect 4571 27860 4583 27863
rect 4614 27860 4620 27872
rect 4571 27832 4620 27860
rect 4571 27829 4583 27832
rect 4525 27823 4583 27829
rect 4614 27820 4620 27832
rect 4672 27820 4678 27872
rect 5350 27820 5356 27872
rect 5408 27860 5414 27872
rect 6086 27860 6092 27872
rect 5408 27832 6092 27860
rect 5408 27820 5414 27832
rect 6086 27820 6092 27832
rect 6144 27820 6150 27872
rect 6825 27863 6883 27869
rect 6825 27829 6837 27863
rect 6871 27860 6883 27863
rect 7377 27863 7435 27869
rect 7377 27860 7389 27863
rect 6871 27832 7389 27860
rect 6871 27829 6883 27832
rect 6825 27823 6883 27829
rect 7377 27829 7389 27832
rect 7423 27860 7435 27863
rect 7650 27860 7656 27872
rect 7423 27832 7656 27860
rect 7423 27829 7435 27832
rect 7377 27823 7435 27829
rect 7650 27820 7656 27832
rect 7708 27820 7714 27872
rect 8481 27863 8539 27869
rect 8481 27829 8493 27863
rect 8527 27860 8539 27863
rect 8849 27863 8907 27869
rect 8849 27860 8861 27863
rect 8527 27832 8861 27860
rect 8527 27829 8539 27832
rect 8481 27823 8539 27829
rect 8849 27829 8861 27832
rect 8895 27860 8907 27863
rect 9585 27863 9643 27869
rect 9585 27860 9597 27863
rect 8895 27832 9597 27860
rect 8895 27829 8907 27832
rect 8849 27823 8907 27829
rect 9585 27829 9597 27832
rect 9631 27860 9643 27863
rect 10318 27860 10324 27872
rect 9631 27832 10324 27860
rect 9631 27829 9643 27832
rect 9585 27823 9643 27829
rect 10318 27820 10324 27832
rect 10376 27860 10382 27872
rect 11238 27860 11244 27872
rect 10376 27832 11244 27860
rect 10376 27820 10382 27832
rect 11238 27820 11244 27832
rect 11296 27820 11302 27872
rect 37918 27820 37924 27872
rect 37976 27860 37982 27872
rect 38197 27863 38255 27869
rect 38197 27860 38209 27863
rect 37976 27832 38209 27860
rect 37976 27820 37982 27832
rect 38197 27829 38209 27832
rect 38243 27829 38255 27863
rect 38197 27823 38255 27829
rect 40218 27820 40224 27872
rect 40276 27860 40282 27872
rect 40313 27863 40371 27869
rect 40313 27860 40325 27863
rect 40276 27832 40325 27860
rect 40276 27820 40282 27832
rect 40313 27829 40325 27832
rect 40359 27829 40371 27863
rect 40313 27823 40371 27829
rect 40402 27820 40408 27872
rect 40460 27860 40466 27872
rect 40589 27863 40647 27869
rect 40589 27860 40601 27863
rect 40460 27832 40601 27860
rect 40460 27820 40466 27832
rect 40589 27829 40601 27832
rect 40635 27829 40647 27863
rect 42168 27860 42196 28104
rect 43272 28104 43484 28132
rect 43548 28104 44680 28132
rect 43272 28073 43300 28104
rect 42245 28067 42303 28073
rect 42245 28033 42257 28067
rect 42291 28033 42303 28067
rect 42245 28027 42303 28033
rect 43257 28067 43315 28073
rect 43257 28033 43269 28067
rect 43303 28033 43315 28067
rect 43257 28027 43315 28033
rect 42260 27996 42288 28027
rect 43438 28024 43444 28076
rect 43496 28024 43502 28076
rect 43548 27996 43576 28104
rect 46382 28092 46388 28144
rect 46440 28092 46446 28144
rect 46845 28135 46903 28141
rect 46845 28101 46857 28135
rect 46891 28132 46903 28135
rect 47118 28132 47124 28144
rect 46891 28104 47124 28132
rect 46891 28101 46903 28104
rect 46845 28095 46903 28101
rect 47118 28092 47124 28104
rect 47176 28092 47182 28144
rect 47305 28135 47363 28141
rect 47305 28101 47317 28135
rect 47351 28132 47363 28135
rect 49068 28132 49096 28160
rect 47351 28104 47532 28132
rect 47351 28101 47363 28104
rect 47305 28095 47363 28101
rect 43717 28067 43775 28073
rect 43717 28033 43729 28067
rect 43763 28033 43775 28067
rect 43717 28027 43775 28033
rect 42260 27968 43576 27996
rect 43622 27956 43628 28008
rect 43680 27996 43686 28008
rect 43732 27996 43760 28027
rect 47210 28024 47216 28076
rect 47268 28024 47274 28076
rect 47397 28067 47455 28073
rect 47397 28033 47409 28067
rect 47443 28033 47455 28067
rect 47397 28027 47455 28033
rect 43993 27999 44051 28005
rect 43993 27996 44005 27999
rect 43680 27968 44005 27996
rect 43680 27956 43686 27968
rect 43993 27965 44005 27968
rect 44039 27965 44051 27999
rect 43993 27959 44051 27965
rect 44634 27956 44640 28008
rect 44692 27996 44698 28008
rect 45373 27999 45431 28005
rect 45373 27996 45385 27999
rect 44692 27968 45385 27996
rect 44692 27956 44698 27968
rect 45373 27965 45385 27968
rect 45419 27965 45431 27999
rect 45373 27959 45431 27965
rect 47118 27956 47124 28008
rect 47176 27956 47182 28008
rect 47412 27860 47440 28027
rect 47504 27996 47532 28104
rect 47596 28104 49096 28132
rect 49513 28135 49571 28141
rect 47596 28076 47624 28104
rect 49513 28101 49525 28135
rect 49559 28132 49571 28135
rect 50172 28132 50200 28160
rect 49559 28104 50200 28132
rect 49559 28101 49571 28104
rect 49513 28095 49571 28101
rect 47578 28024 47584 28076
rect 47636 28024 47642 28076
rect 47854 28024 47860 28076
rect 47912 28024 47918 28076
rect 48501 28067 48559 28073
rect 48501 28064 48513 28067
rect 47956 28036 48513 28064
rect 47956 27996 47984 28036
rect 48501 28033 48513 28036
rect 48547 28064 48559 28067
rect 49145 28067 49203 28073
rect 49145 28064 49157 28067
rect 48547 28036 49157 28064
rect 48547 28033 48559 28036
rect 48501 28027 48559 28033
rect 49145 28033 49157 28036
rect 49191 28033 49203 28067
rect 49145 28027 49203 28033
rect 49234 28024 49240 28076
rect 49292 28064 49298 28076
rect 49620 28073 49648 28104
rect 51902 28092 51908 28144
rect 51960 28132 51966 28144
rect 56502 28132 56508 28144
rect 51960 28104 56508 28132
rect 51960 28092 51966 28104
rect 49329 28067 49387 28073
rect 49329 28064 49341 28067
rect 49292 28036 49341 28064
rect 49292 28024 49298 28036
rect 49329 28033 49341 28036
rect 49375 28033 49387 28067
rect 49329 28027 49387 28033
rect 49605 28067 49663 28073
rect 49605 28033 49617 28067
rect 49651 28064 49663 28067
rect 49789 28067 49847 28073
rect 49651 28036 49685 28064
rect 49651 28033 49663 28036
rect 49605 28027 49663 28033
rect 49789 28033 49801 28067
rect 49835 28064 49847 28067
rect 50154 28064 50160 28076
rect 49835 28036 50160 28064
rect 49835 28033 49847 28036
rect 49789 28027 49847 28033
rect 47504 27968 47984 27996
rect 48133 27999 48191 28005
rect 48133 27965 48145 27999
rect 48179 27965 48191 27999
rect 48133 27959 48191 27965
rect 47581 27931 47639 27937
rect 47581 27897 47593 27931
rect 47627 27928 47639 27931
rect 47762 27928 47768 27940
rect 47627 27900 47768 27928
rect 47627 27897 47639 27900
rect 47581 27891 47639 27897
rect 47762 27888 47768 27900
rect 47820 27888 47826 27940
rect 47946 27888 47952 27940
rect 48004 27928 48010 27940
rect 48148 27928 48176 27959
rect 48222 27956 48228 28008
rect 48280 27996 48286 28008
rect 48409 27999 48467 28005
rect 48409 27996 48421 27999
rect 48280 27968 48421 27996
rect 48280 27956 48286 27968
rect 48409 27965 48421 27968
rect 48455 27965 48467 27999
rect 48409 27959 48467 27965
rect 49418 27956 49424 28008
rect 49476 27996 49482 28008
rect 49804 27996 49832 28027
rect 50154 28024 50160 28036
rect 50212 28024 50218 28076
rect 51166 28024 51172 28076
rect 51224 28064 51230 28076
rect 52362 28064 52368 28076
rect 51224 28036 52368 28064
rect 51224 28024 51230 28036
rect 52362 28024 52368 28036
rect 52420 28024 52426 28076
rect 52546 28024 52552 28076
rect 52604 28064 52610 28076
rect 53484 28073 53512 28104
rect 52733 28067 52791 28073
rect 52733 28064 52745 28067
rect 52604 28036 52745 28064
rect 52604 28024 52610 28036
rect 52733 28033 52745 28036
rect 52779 28033 52791 28067
rect 52733 28027 52791 28033
rect 53469 28067 53527 28073
rect 53469 28033 53481 28067
rect 53515 28033 53527 28067
rect 53469 28027 53527 28033
rect 53736 28067 53794 28073
rect 53736 28033 53748 28067
rect 53782 28064 53794 28067
rect 54018 28064 54024 28076
rect 53782 28036 54024 28064
rect 53782 28033 53794 28036
rect 53736 28027 53794 28033
rect 54018 28024 54024 28036
rect 54076 28024 54082 28076
rect 56152 28073 56180 28104
rect 56502 28092 56508 28104
rect 56560 28092 56566 28144
rect 56778 28092 56784 28144
rect 56836 28132 56842 28144
rect 58820 28132 58848 28160
rect 56836 28104 58848 28132
rect 56836 28092 56842 28104
rect 56410 28073 56416 28076
rect 55953 28067 56011 28073
rect 55953 28033 55965 28067
rect 55999 28033 56011 28067
rect 55953 28027 56011 28033
rect 56137 28067 56195 28073
rect 56137 28033 56149 28067
rect 56183 28033 56195 28067
rect 56137 28027 56195 28033
rect 56404 28027 56416 28073
rect 49476 27968 49832 27996
rect 52273 27999 52331 28005
rect 49476 27956 49482 27968
rect 52273 27965 52285 27999
rect 52319 27996 52331 27999
rect 52457 27999 52515 28005
rect 52457 27996 52469 27999
rect 52319 27968 52469 27996
rect 52319 27965 52331 27968
rect 52273 27959 52331 27965
rect 52457 27965 52469 27968
rect 52503 27965 52515 27999
rect 52457 27959 52515 27965
rect 52914 27956 52920 28008
rect 52972 27996 52978 28008
rect 53285 27999 53343 28005
rect 53285 27996 53297 27999
rect 52972 27968 53297 27996
rect 52972 27956 52978 27968
rect 53285 27965 53297 27968
rect 53331 27965 53343 27999
rect 54941 27999 54999 28005
rect 54941 27996 54953 27999
rect 53285 27959 53343 27965
rect 54864 27968 54953 27996
rect 54864 27937 54892 27968
rect 54941 27965 54953 27968
rect 54987 27965 54999 27999
rect 54941 27959 54999 27965
rect 55674 27956 55680 28008
rect 55732 27956 55738 28008
rect 48004 27900 48176 27928
rect 54849 27931 54907 27937
rect 48004 27888 48010 27900
rect 54849 27897 54861 27931
rect 54895 27897 54907 27931
rect 55968 27928 55996 28027
rect 56410 28024 56416 28027
rect 56468 28024 56474 28076
rect 58437 27999 58495 28005
rect 58437 27965 58449 27999
rect 58483 27965 58495 27999
rect 58437 27959 58495 27965
rect 54849 27891 54907 27897
rect 55600 27900 55996 27928
rect 57517 27931 57575 27937
rect 48130 27860 48136 27872
rect 42168 27832 48136 27860
rect 40589 27823 40647 27829
rect 48130 27820 48136 27832
rect 48188 27820 48194 27872
rect 48222 27820 48228 27872
rect 48280 27860 48286 27872
rect 49970 27860 49976 27872
rect 48280 27832 49976 27860
rect 48280 27820 48286 27832
rect 49970 27820 49976 27832
rect 50028 27820 50034 27872
rect 51626 27820 51632 27872
rect 51684 27820 51690 27872
rect 55030 27820 55036 27872
rect 55088 27860 55094 27872
rect 55600 27869 55628 27900
rect 57517 27897 57529 27931
rect 57563 27928 57575 27931
rect 58452 27928 58480 27959
rect 57563 27900 58480 27928
rect 57563 27897 57575 27900
rect 57517 27891 57575 27897
rect 55585 27863 55643 27869
rect 55585 27860 55597 27863
rect 55088 27832 55597 27860
rect 55088 27820 55094 27832
rect 55585 27829 55597 27832
rect 55631 27829 55643 27863
rect 55585 27823 55643 27829
rect 55858 27820 55864 27872
rect 55916 27820 55922 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 3329 27659 3387 27665
rect 3329 27625 3341 27659
rect 3375 27656 3387 27659
rect 3418 27656 3424 27668
rect 3375 27628 3424 27656
rect 3375 27625 3387 27628
rect 3329 27619 3387 27625
rect 3418 27616 3424 27628
rect 3476 27616 3482 27668
rect 4614 27656 4620 27668
rect 4172 27628 4620 27656
rect 3234 27548 3240 27600
rect 3292 27548 3298 27600
rect 3145 27523 3203 27529
rect 3145 27489 3157 27523
rect 3191 27520 3203 27523
rect 3252 27520 3280 27548
rect 3191 27492 3280 27520
rect 3191 27489 3203 27492
rect 3145 27483 3203 27489
rect 3234 27412 3240 27464
rect 3292 27412 3298 27464
rect 3418 27412 3424 27464
rect 3476 27412 3482 27464
rect 3973 27455 4031 27461
rect 3973 27421 3985 27455
rect 4019 27452 4031 27455
rect 4172 27452 4200 27628
rect 4614 27616 4620 27628
rect 4672 27616 4678 27668
rect 10962 27616 10968 27668
rect 11020 27656 11026 27668
rect 11330 27656 11336 27668
rect 11020 27628 11336 27656
rect 11020 27616 11026 27628
rect 11330 27616 11336 27628
rect 11388 27616 11394 27668
rect 39666 27656 39672 27668
rect 14108 27628 15056 27656
rect 4249 27591 4307 27597
rect 4249 27557 4261 27591
rect 4295 27557 4307 27591
rect 4249 27551 4307 27557
rect 13449 27591 13507 27597
rect 13449 27557 13461 27591
rect 13495 27588 13507 27591
rect 14108 27588 14136 27628
rect 13495 27560 14136 27588
rect 15028 27588 15056 27628
rect 38856 27628 39672 27656
rect 15473 27591 15531 27597
rect 15028 27560 15148 27588
rect 13495 27557 13507 27560
rect 13449 27551 13507 27557
rect 4019 27424 4200 27452
rect 4264 27452 4292 27551
rect 6822 27480 6828 27532
rect 6880 27520 6886 27532
rect 7285 27523 7343 27529
rect 7285 27520 7297 27523
rect 6880 27492 7297 27520
rect 6880 27480 6886 27492
rect 7285 27489 7297 27492
rect 7331 27489 7343 27523
rect 7285 27483 7343 27489
rect 8386 27480 8392 27532
rect 8444 27520 8450 27532
rect 8846 27520 8852 27532
rect 8444 27492 8852 27520
rect 8444 27480 8450 27492
rect 8846 27480 8852 27492
rect 8904 27480 8910 27532
rect 9769 27523 9827 27529
rect 9769 27489 9781 27523
rect 9815 27520 9827 27523
rect 10410 27520 10416 27532
rect 9815 27492 10416 27520
rect 9815 27489 9827 27492
rect 9769 27483 9827 27489
rect 10410 27480 10416 27492
rect 10468 27480 10474 27532
rect 13464 27520 13492 27551
rect 12820 27492 13492 27520
rect 14016 27492 14228 27520
rect 12820 27464 12848 27492
rect 5454 27455 5512 27461
rect 5454 27452 5466 27455
rect 4264 27424 5466 27452
rect 4019 27421 4031 27424
rect 3973 27415 4031 27421
rect 5454 27421 5466 27424
rect 5500 27421 5512 27455
rect 5454 27415 5512 27421
rect 5626 27412 5632 27464
rect 5684 27452 5690 27464
rect 5721 27455 5779 27461
rect 5721 27452 5733 27455
rect 5684 27424 5733 27452
rect 5684 27412 5690 27424
rect 5721 27421 5733 27424
rect 5767 27421 5779 27455
rect 5721 27415 5779 27421
rect 6454 27412 6460 27464
rect 6512 27412 6518 27464
rect 6546 27412 6552 27464
rect 6604 27452 6610 27464
rect 7009 27455 7067 27461
rect 7009 27452 7021 27455
rect 6604 27424 7021 27452
rect 6604 27412 6610 27424
rect 7009 27421 7021 27424
rect 7055 27421 7067 27455
rect 7009 27415 7067 27421
rect 7466 27412 7472 27464
rect 7524 27412 7530 27464
rect 10045 27455 10103 27461
rect 10045 27421 10057 27455
rect 10091 27452 10103 27455
rect 10226 27452 10232 27464
rect 10091 27424 10232 27452
rect 10091 27421 10103 27424
rect 10045 27415 10103 27421
rect 10226 27412 10232 27424
rect 10284 27452 10290 27464
rect 10689 27455 10747 27461
rect 10689 27452 10701 27455
rect 10284 27424 10701 27452
rect 10284 27412 10290 27424
rect 10689 27421 10701 27424
rect 10735 27421 10747 27455
rect 10689 27415 10747 27421
rect 12342 27412 12348 27464
rect 12400 27452 12406 27464
rect 12400 27424 12572 27452
rect 12400 27412 12406 27424
rect 2406 27344 2412 27396
rect 2464 27344 2470 27396
rect 2866 27344 2872 27396
rect 2924 27344 2930 27396
rect 4065 27387 4123 27393
rect 4065 27353 4077 27387
rect 4111 27384 4123 27387
rect 4154 27384 4160 27396
rect 4111 27356 4160 27384
rect 4111 27353 4123 27356
rect 4065 27347 4123 27353
rect 4154 27344 4160 27356
rect 4212 27344 4218 27396
rect 4249 27387 4307 27393
rect 4249 27353 4261 27387
rect 4295 27384 4307 27387
rect 5258 27384 5264 27396
rect 4295 27356 5264 27384
rect 4295 27353 4307 27356
rect 4249 27347 4307 27353
rect 5258 27344 5264 27356
rect 5316 27344 5322 27396
rect 6641 27387 6699 27393
rect 6641 27353 6653 27387
rect 6687 27384 6699 27387
rect 6825 27387 6883 27393
rect 6825 27384 6837 27387
rect 6687 27356 6837 27384
rect 6687 27353 6699 27356
rect 6641 27347 6699 27353
rect 6825 27353 6837 27356
rect 6871 27384 6883 27387
rect 7650 27384 7656 27396
rect 6871 27356 7656 27384
rect 6871 27353 6883 27356
rect 6825 27347 6883 27353
rect 7650 27344 7656 27356
rect 7708 27384 7714 27396
rect 10413 27387 10471 27393
rect 7708 27356 8064 27384
rect 7708 27344 7714 27356
rect 1397 27319 1455 27325
rect 1397 27285 1409 27319
rect 1443 27316 1455 27319
rect 2682 27316 2688 27328
rect 1443 27288 2688 27316
rect 1443 27285 1455 27288
rect 1397 27279 1455 27285
rect 2682 27276 2688 27288
rect 2740 27276 2746 27328
rect 4341 27319 4399 27325
rect 4341 27285 4353 27319
rect 4387 27316 4399 27319
rect 4798 27316 4804 27328
rect 4387 27288 4804 27316
rect 4387 27285 4399 27288
rect 4341 27279 4399 27285
rect 4798 27276 4804 27288
rect 4856 27316 4862 27328
rect 5166 27316 5172 27328
rect 4856 27288 5172 27316
rect 4856 27276 4862 27288
rect 5166 27276 5172 27288
rect 5224 27276 5230 27328
rect 6270 27276 6276 27328
rect 6328 27276 6334 27328
rect 6730 27276 6736 27328
rect 6788 27316 6794 27328
rect 8036 27325 8064 27356
rect 10413 27353 10425 27387
rect 10459 27384 10471 27387
rect 11238 27384 11244 27396
rect 10459 27356 11244 27384
rect 10459 27353 10471 27356
rect 10413 27347 10471 27353
rect 11238 27344 11244 27356
rect 11296 27344 11302 27396
rect 11330 27344 11336 27396
rect 11388 27384 11394 27396
rect 12078 27387 12136 27393
rect 12078 27384 12090 27387
rect 11388 27356 12090 27384
rect 11388 27344 11394 27356
rect 12078 27353 12090 27356
rect 12124 27353 12136 27387
rect 12078 27347 12136 27353
rect 7193 27319 7251 27325
rect 7193 27316 7205 27319
rect 6788 27288 7205 27316
rect 6788 27276 6794 27288
rect 7193 27285 7205 27288
rect 7239 27285 7251 27319
rect 7193 27279 7251 27285
rect 8021 27319 8079 27325
rect 8021 27285 8033 27319
rect 8067 27316 8079 27319
rect 8202 27316 8208 27328
rect 8067 27288 8208 27316
rect 8067 27285 8079 27288
rect 8021 27279 8079 27285
rect 8202 27276 8208 27288
rect 8260 27276 8266 27328
rect 11974 27276 11980 27328
rect 12032 27316 12038 27328
rect 12437 27319 12495 27325
rect 12437 27316 12449 27319
rect 12032 27288 12449 27316
rect 12032 27276 12038 27288
rect 12437 27285 12449 27288
rect 12483 27285 12495 27319
rect 12544 27316 12572 27424
rect 12618 27412 12624 27464
rect 12676 27412 12682 27464
rect 12802 27412 12808 27464
rect 12860 27412 12866 27464
rect 12894 27412 12900 27464
rect 12952 27452 12958 27464
rect 12989 27455 13047 27461
rect 12989 27452 13001 27455
rect 12952 27424 13001 27452
rect 12952 27412 12958 27424
rect 12989 27421 13001 27424
rect 13035 27421 13047 27455
rect 12989 27415 13047 27421
rect 13170 27412 13176 27464
rect 13228 27412 13234 27464
rect 13081 27387 13139 27393
rect 13081 27353 13093 27387
rect 13127 27384 13139 27387
rect 14016 27384 14044 27492
rect 14093 27455 14151 27461
rect 14093 27421 14105 27455
rect 14139 27421 14151 27455
rect 14200 27452 14228 27492
rect 14349 27455 14407 27461
rect 14349 27452 14361 27455
rect 14200 27424 14361 27452
rect 14093 27415 14151 27421
rect 14349 27421 14361 27424
rect 14395 27421 14407 27455
rect 15120 27452 15148 27560
rect 15473 27557 15485 27591
rect 15519 27588 15531 27591
rect 38105 27591 38163 27597
rect 15519 27560 31754 27588
rect 15519 27557 15531 27560
rect 15473 27551 15531 27557
rect 31726 27520 31754 27560
rect 38105 27557 38117 27591
rect 38151 27588 38163 27591
rect 38856 27588 38884 27628
rect 39666 27616 39672 27628
rect 39724 27616 39730 27668
rect 40034 27616 40040 27668
rect 40092 27616 40098 27668
rect 40310 27616 40316 27668
rect 40368 27616 40374 27668
rect 42978 27616 42984 27668
rect 43036 27616 43042 27668
rect 43438 27616 43444 27668
rect 43496 27656 43502 27668
rect 43533 27659 43591 27665
rect 43533 27656 43545 27659
rect 43496 27628 43545 27656
rect 43496 27616 43502 27628
rect 43533 27625 43545 27628
rect 43579 27656 43591 27659
rect 43714 27656 43720 27668
rect 43579 27628 43720 27656
rect 43579 27625 43591 27628
rect 43533 27619 43591 27625
rect 43714 27616 43720 27628
rect 43772 27616 43778 27668
rect 43993 27659 44051 27665
rect 43993 27625 44005 27659
rect 44039 27656 44051 27659
rect 44039 27628 45876 27656
rect 44039 27625 44051 27628
rect 43993 27619 44051 27625
rect 38151 27560 38884 27588
rect 38933 27591 38991 27597
rect 38151 27557 38163 27560
rect 38105 27551 38163 27557
rect 38933 27557 38945 27591
rect 38979 27588 38991 27591
rect 40052 27588 40080 27616
rect 38979 27560 40080 27588
rect 38979 27557 38991 27560
rect 38933 27551 38991 27557
rect 38197 27523 38255 27529
rect 31726 27492 38148 27520
rect 24581 27455 24639 27461
rect 24581 27452 24593 27455
rect 15120 27424 24593 27452
rect 14349 27415 14407 27421
rect 24581 27421 24593 27424
rect 24627 27452 24639 27455
rect 25777 27455 25835 27461
rect 25777 27452 25789 27455
rect 24627 27424 25789 27452
rect 24627 27421 24639 27424
rect 24581 27415 24639 27421
rect 25777 27421 25789 27424
rect 25823 27452 25835 27455
rect 25823 27424 26234 27452
rect 25823 27421 25835 27424
rect 25777 27415 25835 27421
rect 13127 27356 14044 27384
rect 13127 27353 13139 27356
rect 13081 27347 13139 27353
rect 13354 27316 13360 27328
rect 12544 27288 13360 27316
rect 12437 27279 12495 27285
rect 13354 27276 13360 27288
rect 13412 27316 13418 27328
rect 13817 27319 13875 27325
rect 13817 27316 13829 27319
rect 13412 27288 13829 27316
rect 13412 27276 13418 27288
rect 13817 27285 13829 27288
rect 13863 27316 13875 27319
rect 14108 27316 14136 27415
rect 25314 27344 25320 27396
rect 25372 27344 25378 27396
rect 26206 27384 26234 27424
rect 37918 27412 37924 27464
rect 37976 27412 37982 27464
rect 38010 27412 38016 27464
rect 38068 27412 38074 27464
rect 38120 27452 38148 27492
rect 38197 27489 38209 27523
rect 38243 27520 38255 27523
rect 39206 27520 39212 27532
rect 38243 27492 39212 27520
rect 38243 27489 38255 27492
rect 38197 27483 38255 27489
rect 38470 27452 38476 27464
rect 38120 27424 38476 27452
rect 38470 27412 38476 27424
rect 38528 27412 38534 27464
rect 38654 27412 38660 27464
rect 38712 27412 38718 27464
rect 38764 27461 38792 27492
rect 39206 27480 39212 27492
rect 39264 27480 39270 27532
rect 40037 27523 40095 27529
rect 40037 27520 40049 27523
rect 39408 27492 40049 27520
rect 39408 27464 39436 27492
rect 40037 27489 40049 27492
rect 40083 27489 40095 27523
rect 40037 27483 40095 27489
rect 40129 27523 40187 27529
rect 40129 27489 40141 27523
rect 40175 27520 40187 27523
rect 40328 27520 40356 27616
rect 40175 27492 40356 27520
rect 40405 27523 40463 27529
rect 40175 27489 40187 27492
rect 40129 27483 40187 27489
rect 40405 27489 40417 27523
rect 40451 27520 40463 27523
rect 40494 27520 40500 27532
rect 40451 27492 40500 27520
rect 40451 27489 40463 27492
rect 40405 27483 40463 27489
rect 40494 27480 40500 27492
rect 40552 27480 40558 27532
rect 38749 27455 38807 27461
rect 38749 27421 38761 27455
rect 38795 27421 38807 27455
rect 38749 27415 38807 27421
rect 39390 27412 39396 27464
rect 39448 27412 39454 27464
rect 39850 27412 39856 27464
rect 39908 27452 39914 27464
rect 39945 27455 40003 27461
rect 39945 27452 39957 27455
rect 39908 27424 39957 27452
rect 39908 27412 39914 27424
rect 39945 27421 39957 27424
rect 39991 27421 40003 27455
rect 39945 27415 40003 27421
rect 40218 27412 40224 27464
rect 40276 27452 40282 27464
rect 40313 27455 40371 27461
rect 40313 27452 40325 27455
rect 40276 27424 40325 27452
rect 40276 27412 40282 27424
rect 40313 27421 40325 27424
rect 40359 27452 40371 27455
rect 40678 27452 40684 27464
rect 40359 27424 40684 27452
rect 40359 27421 40371 27424
rect 40313 27415 40371 27421
rect 40678 27412 40684 27424
rect 40736 27412 40742 27464
rect 42996 27452 43024 27616
rect 43898 27520 43904 27532
rect 43456 27492 43904 27520
rect 43456 27461 43484 27492
rect 43898 27480 43904 27492
rect 43956 27480 43962 27532
rect 43633 27462 43691 27463
rect 43441 27455 43499 27461
rect 43441 27452 43453 27455
rect 42996 27424 43453 27452
rect 43441 27421 43453 27424
rect 43487 27421 43499 27455
rect 43441 27415 43499 27421
rect 43633 27457 43852 27462
rect 43633 27423 43645 27457
rect 43679 27452 43852 27457
rect 44008 27452 44036 27619
rect 45848 27600 45876 27628
rect 46382 27616 46388 27668
rect 46440 27656 46446 27668
rect 47305 27659 47363 27665
rect 47305 27656 47317 27659
rect 46440 27628 47317 27656
rect 46440 27616 46446 27628
rect 47305 27625 47317 27628
rect 47351 27656 47363 27659
rect 47673 27659 47731 27665
rect 47673 27656 47685 27659
rect 47351 27628 47685 27656
rect 47351 27625 47363 27628
rect 47305 27619 47363 27625
rect 47673 27625 47685 27628
rect 47719 27656 47731 27659
rect 47946 27656 47952 27668
rect 47719 27628 47952 27656
rect 47719 27625 47731 27628
rect 47673 27619 47731 27625
rect 47946 27616 47952 27628
rect 48004 27616 48010 27668
rect 52549 27659 52607 27665
rect 52549 27625 52561 27659
rect 52595 27656 52607 27659
rect 52914 27656 52920 27668
rect 52595 27628 52920 27656
rect 52595 27625 52607 27628
rect 52549 27619 52607 27625
rect 52914 27616 52920 27628
rect 52972 27616 52978 27668
rect 53190 27616 53196 27668
rect 53248 27616 53254 27668
rect 54018 27616 54024 27668
rect 54076 27616 54082 27668
rect 55401 27659 55459 27665
rect 55401 27625 55413 27659
rect 55447 27656 55459 27659
rect 55674 27656 55680 27668
rect 55447 27628 55680 27656
rect 55447 27625 55459 27628
rect 55401 27619 55459 27625
rect 55674 27616 55680 27628
rect 55732 27616 55738 27668
rect 56410 27616 56416 27668
rect 56468 27616 56474 27668
rect 58342 27616 58348 27668
rect 58400 27616 58406 27668
rect 44910 27588 44916 27600
rect 44468 27560 44916 27588
rect 44468 27461 44496 27560
rect 44910 27548 44916 27560
rect 44968 27588 44974 27600
rect 45097 27591 45155 27597
rect 45097 27588 45109 27591
rect 44968 27560 45109 27588
rect 44968 27548 44974 27560
rect 45097 27557 45109 27560
rect 45143 27557 45155 27591
rect 45097 27551 45155 27557
rect 45830 27548 45836 27600
rect 45888 27548 45894 27600
rect 46014 27548 46020 27600
rect 46072 27588 46078 27600
rect 50614 27588 50620 27600
rect 46072 27560 50620 27588
rect 46072 27548 46078 27560
rect 45756 27492 49648 27520
rect 44453 27455 44511 27461
rect 44453 27452 44465 27455
rect 43679 27434 44036 27452
rect 43679 27423 43691 27434
rect 43824 27424 44036 27434
rect 44100 27424 44465 27452
rect 43633 27417 43691 27423
rect 26206 27356 43668 27384
rect 13863 27288 14136 27316
rect 13863 27285 13875 27288
rect 13817 27279 13875 27285
rect 38654 27276 38660 27328
rect 38712 27316 38718 27328
rect 39206 27316 39212 27328
rect 38712 27288 39212 27316
rect 38712 27276 38718 27288
rect 39206 27276 39212 27288
rect 39264 27276 39270 27328
rect 39298 27276 39304 27328
rect 39356 27316 39362 27328
rect 39853 27319 39911 27325
rect 39853 27316 39865 27319
rect 39356 27288 39865 27316
rect 39356 27276 39362 27288
rect 39853 27285 39865 27288
rect 39899 27285 39911 27319
rect 39853 27279 39911 27285
rect 42150 27276 42156 27328
rect 42208 27276 42214 27328
rect 42886 27276 42892 27328
rect 42944 27316 42950 27328
rect 43530 27316 43536 27328
rect 42944 27288 43536 27316
rect 42944 27276 42950 27288
rect 43530 27276 43536 27288
rect 43588 27276 43594 27328
rect 43640 27316 43668 27356
rect 44100 27316 44128 27424
rect 44453 27421 44465 27424
rect 44499 27421 44511 27455
rect 44453 27415 44511 27421
rect 44818 27412 44824 27464
rect 44876 27452 44882 27464
rect 45005 27455 45063 27461
rect 45005 27452 45017 27455
rect 44876 27424 45017 27452
rect 44876 27412 44882 27424
rect 45005 27421 45017 27424
rect 45051 27421 45063 27455
rect 45005 27415 45063 27421
rect 45020 27384 45048 27415
rect 45646 27412 45652 27464
rect 45704 27452 45710 27464
rect 45756 27461 45784 27492
rect 45741 27455 45799 27461
rect 45741 27452 45753 27455
rect 45704 27424 45753 27452
rect 45704 27412 45710 27424
rect 45741 27421 45753 27424
rect 45787 27421 45799 27455
rect 45741 27415 45799 27421
rect 45922 27412 45928 27464
rect 45980 27412 45986 27464
rect 46109 27455 46167 27461
rect 46109 27421 46121 27455
rect 46155 27452 46167 27455
rect 46474 27452 46480 27464
rect 46155 27424 46480 27452
rect 46155 27421 46167 27424
rect 46109 27415 46167 27421
rect 45278 27384 45284 27396
rect 45020 27356 45284 27384
rect 45278 27344 45284 27356
rect 45336 27384 45342 27396
rect 45833 27387 45891 27393
rect 45833 27384 45845 27387
rect 45336 27356 45845 27384
rect 45336 27344 45342 27356
rect 45833 27353 45845 27356
rect 45879 27353 45891 27387
rect 45833 27347 45891 27353
rect 43640 27288 44128 27316
rect 44726 27276 44732 27328
rect 44784 27276 44790 27328
rect 45738 27276 45744 27328
rect 45796 27316 45802 27328
rect 46124 27316 46152 27415
rect 46474 27412 46480 27424
rect 46532 27412 46538 27464
rect 47762 27412 47768 27464
rect 47820 27452 47826 27464
rect 47949 27455 48007 27461
rect 47949 27452 47961 27455
rect 47820 27424 47961 27452
rect 47820 27412 47826 27424
rect 47949 27421 47961 27424
rect 47995 27421 48007 27455
rect 47949 27415 48007 27421
rect 48130 27412 48136 27464
rect 48188 27452 48194 27464
rect 48225 27455 48283 27461
rect 48225 27452 48237 27455
rect 48188 27424 48237 27452
rect 48188 27412 48194 27424
rect 48225 27421 48237 27424
rect 48271 27421 48283 27455
rect 48225 27415 48283 27421
rect 48314 27412 48320 27464
rect 48372 27412 48378 27464
rect 48501 27455 48559 27461
rect 48501 27421 48513 27455
rect 48547 27452 48559 27455
rect 48590 27452 48596 27464
rect 48547 27424 48596 27452
rect 48547 27421 48559 27424
rect 48501 27415 48559 27421
rect 48041 27387 48099 27393
rect 48041 27353 48053 27387
rect 48087 27384 48099 27387
rect 48516 27384 48544 27415
rect 48590 27412 48596 27424
rect 48648 27452 48654 27464
rect 49050 27452 49056 27464
rect 48648 27424 49056 27452
rect 48648 27412 48654 27424
rect 49050 27412 49056 27424
rect 49108 27412 49114 27464
rect 49620 27393 49648 27492
rect 49896 27461 49924 27560
rect 50614 27548 50620 27560
rect 50672 27548 50678 27600
rect 53837 27591 53895 27597
rect 53837 27557 53849 27591
rect 53883 27588 53895 27591
rect 54036 27588 54064 27616
rect 56505 27591 56563 27597
rect 56505 27588 56517 27591
rect 53883 27560 54064 27588
rect 56152 27560 56517 27588
rect 53883 27557 53895 27560
rect 53837 27551 53895 27557
rect 56152 27532 56180 27560
rect 56505 27557 56517 27560
rect 56551 27588 56563 27591
rect 56778 27588 56784 27600
rect 56551 27560 56784 27588
rect 56551 27557 56563 27560
rect 56505 27551 56563 27557
rect 56778 27548 56784 27560
rect 56836 27548 56842 27600
rect 57977 27591 58035 27597
rect 57977 27557 57989 27591
rect 58023 27557 58035 27591
rect 57977 27551 58035 27557
rect 53745 27523 53803 27529
rect 53745 27489 53757 27523
rect 53791 27520 53803 27523
rect 54113 27523 54171 27529
rect 54113 27520 54125 27523
rect 53791 27492 54125 27520
rect 53791 27489 53803 27492
rect 53745 27483 53803 27489
rect 54113 27489 54125 27492
rect 54159 27489 54171 27523
rect 54113 27483 54171 27489
rect 54757 27523 54815 27529
rect 54757 27489 54769 27523
rect 54803 27520 54815 27523
rect 54941 27523 54999 27529
rect 54941 27520 54953 27523
rect 54803 27492 54953 27520
rect 54803 27489 54815 27492
rect 54757 27483 54815 27489
rect 54941 27489 54953 27492
rect 54987 27489 54999 27523
rect 54941 27483 54999 27489
rect 56134 27480 56140 27532
rect 56192 27480 56198 27532
rect 56321 27523 56379 27529
rect 56321 27489 56333 27523
rect 56367 27520 56379 27523
rect 56689 27523 56747 27529
rect 56689 27520 56701 27523
rect 56367 27492 56701 27520
rect 56367 27489 56379 27492
rect 56321 27483 56379 27489
rect 56689 27489 56701 27492
rect 56735 27489 56747 27523
rect 56870 27520 56876 27532
rect 56689 27483 56747 27489
rect 56796 27492 56876 27520
rect 49789 27455 49847 27461
rect 49789 27421 49801 27455
rect 49835 27421 49847 27455
rect 49789 27415 49847 27421
rect 49881 27455 49939 27461
rect 49881 27421 49893 27455
rect 49927 27421 49939 27455
rect 49881 27415 49939 27421
rect 48087 27356 48544 27384
rect 49605 27387 49663 27393
rect 48087 27353 48099 27356
rect 48041 27347 48099 27353
rect 49605 27353 49617 27387
rect 49651 27384 49663 27387
rect 49694 27384 49700 27396
rect 49651 27356 49700 27384
rect 49651 27353 49663 27356
rect 49605 27347 49663 27353
rect 49694 27344 49700 27356
rect 49752 27344 49758 27396
rect 49804 27384 49832 27415
rect 49970 27412 49976 27464
rect 50028 27452 50034 27464
rect 50341 27455 50399 27461
rect 50341 27452 50353 27455
rect 50028 27424 50353 27452
rect 50028 27412 50034 27424
rect 50341 27421 50353 27424
rect 50387 27452 50399 27455
rect 50982 27452 50988 27464
rect 50387 27424 50988 27452
rect 50387 27421 50399 27424
rect 50341 27415 50399 27421
rect 50982 27412 50988 27424
rect 51040 27412 51046 27464
rect 51169 27455 51227 27461
rect 51169 27421 51181 27455
rect 51215 27452 51227 27455
rect 51902 27452 51908 27464
rect 51215 27424 51908 27452
rect 51215 27421 51227 27424
rect 51169 27415 51227 27421
rect 51902 27412 51908 27424
rect 51960 27412 51966 27464
rect 53101 27455 53159 27461
rect 53101 27452 53113 27455
rect 53024 27424 53113 27452
rect 51442 27393 51448 27396
rect 50249 27387 50307 27393
rect 50249 27384 50261 27387
rect 49804 27356 50261 27384
rect 50249 27353 50261 27356
rect 50295 27384 50307 27387
rect 50295 27356 50936 27384
rect 50295 27353 50307 27356
rect 50249 27347 50307 27353
rect 50908 27328 50936 27356
rect 51436 27347 51448 27393
rect 51442 27344 51448 27347
rect 51500 27344 51506 27396
rect 53024 27328 53052 27424
rect 53101 27421 53113 27424
rect 53147 27421 53159 27455
rect 53101 27415 53159 27421
rect 53285 27455 53343 27461
rect 53285 27421 53297 27455
rect 53331 27452 53343 27455
rect 53834 27452 53840 27464
rect 53331 27424 53840 27452
rect 53331 27421 53343 27424
rect 53285 27415 53343 27421
rect 53834 27412 53840 27424
rect 53892 27412 53898 27464
rect 53929 27455 53987 27461
rect 53929 27421 53941 27455
rect 53975 27421 53987 27455
rect 53929 27415 53987 27421
rect 54021 27455 54079 27461
rect 54021 27421 54033 27455
rect 54067 27421 54079 27455
rect 54021 27415 54079 27421
rect 45796 27288 46152 27316
rect 45796 27276 45802 27288
rect 48682 27276 48688 27328
rect 48740 27276 48746 27328
rect 48774 27276 48780 27328
rect 48832 27316 48838 27328
rect 48961 27319 49019 27325
rect 48961 27316 48973 27319
rect 48832 27288 48973 27316
rect 48832 27276 48838 27288
rect 48961 27285 48973 27288
rect 49007 27316 49019 27319
rect 49234 27316 49240 27328
rect 49007 27288 49240 27316
rect 49007 27285 49019 27288
rect 48961 27279 49019 27285
rect 49234 27276 49240 27288
rect 49292 27276 49298 27328
rect 50890 27276 50896 27328
rect 50948 27276 50954 27328
rect 53006 27276 53012 27328
rect 53064 27276 53070 27328
rect 53834 27276 53840 27328
rect 53892 27316 53898 27328
rect 53944 27316 53972 27415
rect 54036 27384 54064 27415
rect 54846 27412 54852 27464
rect 54904 27412 54910 27464
rect 55030 27412 55036 27464
rect 55088 27412 55094 27464
rect 55309 27455 55367 27461
rect 55309 27421 55321 27455
rect 55355 27421 55367 27455
rect 55309 27415 55367 27421
rect 55493 27455 55551 27461
rect 55493 27421 55505 27455
rect 55539 27452 55551 27455
rect 55858 27452 55864 27464
rect 55539 27424 55864 27452
rect 55539 27421 55551 27424
rect 55493 27415 55551 27421
rect 55324 27384 55352 27415
rect 55858 27412 55864 27424
rect 55916 27452 55922 27464
rect 56410 27452 56416 27464
rect 55916 27424 56416 27452
rect 55916 27412 55922 27424
rect 56410 27412 56416 27424
rect 56468 27412 56474 27464
rect 56594 27412 56600 27464
rect 56652 27412 56658 27464
rect 56796 27452 56824 27492
rect 56870 27480 56876 27492
rect 56928 27480 56934 27532
rect 57333 27523 57391 27529
rect 57333 27489 57345 27523
rect 57379 27520 57391 27523
rect 57517 27523 57575 27529
rect 57517 27520 57529 27523
rect 57379 27492 57529 27520
rect 57379 27489 57391 27492
rect 57333 27483 57391 27489
rect 57517 27489 57529 27492
rect 57563 27489 57575 27523
rect 57517 27483 57575 27489
rect 56704 27424 56824 27452
rect 57425 27455 57483 27461
rect 56704 27384 56732 27424
rect 57425 27421 57437 27455
rect 57471 27421 57483 27455
rect 57425 27415 57483 27421
rect 57609 27455 57667 27461
rect 57609 27421 57621 27455
rect 57655 27452 57667 27455
rect 57698 27452 57704 27464
rect 57655 27424 57704 27452
rect 57655 27421 57667 27424
rect 57609 27415 57667 27421
rect 54036 27356 56732 27384
rect 54938 27316 54944 27328
rect 53892 27288 54944 27316
rect 53892 27276 53898 27288
rect 54938 27276 54944 27288
rect 54996 27316 55002 27328
rect 56134 27316 56140 27328
rect 54996 27288 56140 27316
rect 54996 27276 55002 27288
rect 56134 27276 56140 27288
rect 56192 27276 56198 27328
rect 56318 27276 56324 27328
rect 56376 27316 56382 27328
rect 57440 27316 57468 27415
rect 57698 27412 57704 27424
rect 57756 27412 57762 27464
rect 57793 27455 57851 27461
rect 57793 27421 57805 27455
rect 57839 27421 57851 27455
rect 57992 27452 58020 27551
rect 58069 27455 58127 27461
rect 58069 27452 58081 27455
rect 57992 27424 58081 27452
rect 57793 27415 57851 27421
rect 58069 27421 58081 27424
rect 58115 27421 58127 27455
rect 58069 27415 58127 27421
rect 58529 27455 58587 27461
rect 58529 27421 58541 27455
rect 58575 27452 58587 27455
rect 58894 27452 58900 27464
rect 58575 27424 58900 27452
rect 58575 27421 58587 27424
rect 58529 27415 58587 27421
rect 57808 27384 57836 27415
rect 58894 27412 58900 27424
rect 58952 27412 58958 27464
rect 58710 27384 58716 27396
rect 57808 27356 58716 27384
rect 58710 27344 58716 27356
rect 58768 27344 58774 27396
rect 56376 27288 57468 27316
rect 56376 27276 56382 27288
rect 58158 27276 58164 27328
rect 58216 27276 58222 27328
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 2685 27115 2743 27121
rect 2685 27081 2697 27115
rect 2731 27112 2743 27115
rect 2866 27112 2872 27124
rect 2731 27084 2872 27112
rect 2731 27081 2743 27084
rect 2685 27075 2743 27081
rect 2866 27072 2872 27084
rect 2924 27072 2930 27124
rect 3418 27072 3424 27124
rect 3476 27112 3482 27124
rect 3881 27115 3939 27121
rect 3881 27112 3893 27115
rect 3476 27084 3893 27112
rect 3476 27072 3482 27084
rect 3881 27081 3893 27084
rect 3927 27081 3939 27115
rect 3881 27075 3939 27081
rect 4154 27072 4160 27124
rect 4212 27112 4218 27124
rect 4617 27115 4675 27121
rect 4617 27112 4629 27115
rect 4212 27084 4629 27112
rect 4212 27072 4218 27084
rect 4617 27081 4629 27084
rect 4663 27112 4675 27115
rect 4706 27112 4712 27124
rect 4663 27084 4712 27112
rect 4663 27081 4675 27084
rect 4617 27075 4675 27081
rect 4706 27072 4712 27084
rect 4764 27072 4770 27124
rect 8941 27115 8999 27121
rect 8941 27081 8953 27115
rect 8987 27081 8999 27115
rect 8941 27075 8999 27081
rect 2777 27047 2835 27053
rect 2777 27013 2789 27047
rect 2823 27013 2835 27047
rect 4065 27047 4123 27053
rect 4065 27044 4077 27047
rect 2777 27007 2835 27013
rect 3068 27016 4077 27044
rect 2133 26979 2191 26985
rect 2133 26945 2145 26979
rect 2179 26976 2191 26979
rect 2792 26976 2820 27007
rect 3068 26985 3096 27016
rect 4065 27013 4077 27016
rect 4111 27013 4123 27047
rect 4065 27007 4123 27013
rect 4801 27047 4859 27053
rect 4801 27013 4813 27047
rect 4847 27044 4859 27047
rect 4847 27016 5120 27044
rect 4847 27013 4859 27016
rect 4801 27007 4859 27013
rect 2179 26948 2820 26976
rect 3053 26979 3111 26985
rect 2179 26945 2191 26948
rect 2133 26939 2191 26945
rect 3053 26945 3065 26979
rect 3099 26945 3111 26979
rect 3053 26939 3111 26945
rect 3973 26979 4031 26985
rect 3973 26945 3985 26979
rect 4019 26945 4031 26979
rect 3973 26939 4031 26945
rect 4157 26979 4215 26985
rect 4157 26945 4169 26979
rect 4203 26945 4215 26979
rect 4157 26939 4215 26945
rect 2774 26868 2780 26920
rect 2832 26868 2838 26920
rect 3237 26911 3295 26917
rect 3237 26877 3249 26911
rect 3283 26877 3295 26911
rect 3237 26871 3295 26877
rect 2682 26800 2688 26852
rect 2740 26840 2746 26852
rect 3252 26840 3280 26871
rect 2740 26812 3280 26840
rect 2740 26800 2746 26812
rect 3786 26800 3792 26852
rect 3844 26840 3850 26852
rect 3988 26840 4016 26939
rect 4172 26908 4200 26939
rect 4982 26936 4988 26988
rect 5040 26936 5046 26988
rect 5092 26976 5120 27016
rect 5166 27004 5172 27056
rect 5224 27044 5230 27056
rect 5997 27047 6055 27053
rect 5997 27044 6009 27047
rect 5224 27016 6009 27044
rect 5224 27004 5230 27016
rect 5997 27013 6009 27016
rect 6043 27013 6055 27047
rect 5997 27007 6055 27013
rect 6270 27004 6276 27056
rect 6328 27004 6334 27056
rect 6362 27004 6368 27056
rect 6420 27044 6426 27056
rect 7466 27044 7472 27056
rect 6420 27016 7472 27044
rect 6420 27004 6426 27016
rect 5626 26976 5632 26988
rect 5092 26948 5632 26976
rect 5626 26936 5632 26948
rect 5684 26936 5690 26988
rect 6086 26936 6092 26988
rect 6144 26976 6150 26988
rect 6181 26979 6239 26985
rect 6181 26976 6193 26979
rect 6144 26948 6193 26976
rect 6144 26936 6150 26948
rect 6181 26945 6193 26948
rect 6227 26945 6239 26979
rect 6181 26939 6239 26945
rect 4614 26908 4620 26920
rect 4172 26880 4620 26908
rect 4614 26868 4620 26880
rect 4672 26868 4678 26920
rect 6288 26908 6316 27004
rect 6641 26979 6699 26985
rect 6641 26945 6653 26979
rect 6687 26976 6699 26979
rect 7009 26979 7067 26985
rect 7009 26976 7021 26979
rect 6687 26948 7021 26976
rect 6687 26945 6699 26948
rect 6641 26939 6699 26945
rect 7009 26945 7021 26948
rect 7055 26945 7067 26979
rect 7009 26939 7067 26945
rect 6365 26911 6423 26917
rect 6365 26908 6377 26911
rect 6288 26880 6377 26908
rect 6365 26877 6377 26880
rect 6411 26877 6423 26911
rect 7024 26908 7052 26939
rect 7190 26936 7196 26988
rect 7248 26936 7254 26988
rect 7300 26985 7328 27016
rect 7466 27004 7472 27016
rect 7524 27004 7530 27056
rect 8956 27044 8984 27075
rect 9950 27072 9956 27124
rect 10008 27112 10014 27124
rect 10597 27115 10655 27121
rect 10597 27112 10609 27115
rect 10008 27084 10609 27112
rect 10008 27072 10014 27084
rect 10597 27081 10609 27084
rect 10643 27081 10655 27115
rect 10597 27075 10655 27081
rect 11330 27072 11336 27124
rect 11388 27072 11394 27124
rect 12802 27112 12808 27124
rect 12084 27084 12808 27112
rect 12084 27053 12112 27084
rect 12802 27072 12808 27084
rect 12860 27072 12866 27124
rect 38010 27072 38016 27124
rect 38068 27112 38074 27124
rect 38473 27115 38531 27121
rect 38473 27112 38485 27115
rect 38068 27084 38485 27112
rect 38068 27072 38074 27084
rect 38473 27081 38485 27084
rect 38519 27081 38531 27115
rect 38473 27075 38531 27081
rect 38562 27072 38568 27124
rect 38620 27112 38626 27124
rect 42886 27112 42892 27124
rect 38620 27084 42892 27112
rect 38620 27072 38626 27084
rect 42886 27072 42892 27084
rect 42944 27072 42950 27124
rect 42978 27072 42984 27124
rect 43036 27072 43042 27124
rect 43070 27072 43076 27124
rect 43128 27072 43134 27124
rect 46106 27112 46112 27124
rect 43456 27084 46112 27112
rect 10321 27047 10379 27053
rect 10321 27044 10333 27047
rect 7576 27016 8984 27044
rect 9048 27016 10333 27044
rect 7285 26979 7343 26985
rect 7285 26945 7297 26979
rect 7331 26945 7343 26979
rect 7576 26976 7604 27016
rect 7834 26985 7840 26988
rect 7828 26976 7840 26985
rect 7285 26939 7343 26945
rect 7484 26948 7604 26976
rect 7795 26948 7840 26976
rect 7484 26908 7512 26948
rect 7828 26939 7840 26948
rect 7834 26936 7840 26939
rect 7892 26936 7898 26988
rect 8202 26936 8208 26988
rect 8260 26976 8266 26988
rect 9048 26976 9076 27016
rect 10321 27013 10333 27016
rect 10367 27044 10379 27047
rect 11057 27047 11115 27053
rect 11057 27044 11069 27047
rect 10367 27016 11069 27044
rect 10367 27013 10379 27016
rect 10321 27007 10379 27013
rect 11057 27013 11069 27016
rect 11103 27044 11115 27047
rect 12069 27047 12127 27053
rect 12069 27044 12081 27047
rect 11103 27016 12081 27044
rect 11103 27013 11115 27016
rect 11057 27007 11115 27013
rect 12069 27013 12081 27016
rect 12115 27013 12127 27047
rect 25314 27044 25320 27056
rect 12069 27007 12127 27013
rect 12406 27016 25320 27044
rect 8260 26948 9076 26976
rect 8260 26936 8266 26948
rect 9766 26936 9772 26988
rect 9824 26976 9830 26988
rect 10137 26979 10195 26985
rect 10137 26976 10149 26979
rect 9824 26948 10149 26976
rect 9824 26936 9830 26948
rect 10137 26945 10149 26948
rect 10183 26945 10195 26979
rect 10137 26939 10195 26945
rect 10410 26936 10416 26988
rect 10468 26936 10474 26988
rect 11149 26979 11207 26985
rect 11149 26945 11161 26979
rect 11195 26976 11207 26979
rect 11514 26976 11520 26988
rect 11195 26948 11520 26976
rect 11195 26945 11207 26948
rect 11149 26939 11207 26945
rect 11514 26936 11520 26948
rect 11572 26936 11578 26988
rect 11698 26936 11704 26988
rect 11756 26976 11762 26988
rect 11885 26979 11943 26985
rect 11885 26976 11897 26979
rect 11756 26948 11897 26976
rect 11756 26936 11762 26948
rect 11885 26945 11897 26948
rect 11931 26945 11943 26979
rect 11885 26939 11943 26945
rect 7024 26880 7512 26908
rect 7561 26911 7619 26917
rect 6365 26871 6423 26877
rect 7561 26877 7573 26911
rect 7607 26877 7619 26911
rect 7561 26871 7619 26877
rect 5074 26840 5080 26852
rect 3844 26812 5080 26840
rect 3844 26800 3850 26812
rect 5074 26800 5080 26812
rect 5132 26800 5138 26852
rect 7377 26843 7435 26849
rect 5184 26812 7236 26840
rect 2961 26775 3019 26781
rect 2961 26741 2973 26775
rect 3007 26772 3019 26775
rect 3326 26772 3332 26784
rect 3007 26744 3332 26772
rect 3007 26741 3019 26744
rect 2961 26735 3019 26741
rect 3326 26732 3332 26744
rect 3384 26772 3390 26784
rect 5184 26772 5212 26812
rect 3384 26744 5212 26772
rect 3384 26732 3390 26744
rect 5810 26732 5816 26784
rect 5868 26732 5874 26784
rect 6178 26732 6184 26784
rect 6236 26772 6242 26784
rect 6457 26775 6515 26781
rect 6457 26772 6469 26775
rect 6236 26744 6469 26772
rect 6236 26732 6242 26744
rect 6457 26741 6469 26744
rect 6503 26741 6515 26775
rect 6457 26735 6515 26741
rect 6546 26732 6552 26784
rect 6604 26732 6610 26784
rect 7098 26732 7104 26784
rect 7156 26732 7162 26784
rect 7208 26772 7236 26812
rect 7377 26809 7389 26843
rect 7423 26840 7435 26843
rect 7576 26840 7604 26871
rect 12406 26840 12434 27016
rect 25314 27004 25320 27016
rect 25372 27004 25378 27056
rect 38102 27004 38108 27056
rect 38160 27044 38166 27056
rect 39390 27044 39396 27056
rect 38160 27016 39396 27044
rect 38160 27004 38166 27016
rect 39390 27004 39396 27016
rect 39448 27004 39454 27056
rect 39669 27047 39727 27053
rect 39669 27013 39681 27047
rect 39715 27044 39727 27047
rect 40497 27047 40555 27053
rect 40497 27044 40509 27047
rect 39715 27016 40509 27044
rect 39715 27013 39727 27016
rect 39669 27007 39727 27013
rect 40497 27013 40509 27016
rect 40543 27013 40555 27047
rect 42150 27044 42156 27056
rect 41722 27016 42156 27044
rect 40497 27007 40555 27013
rect 42150 27004 42156 27016
rect 42208 27004 42214 27056
rect 42996 27044 43024 27072
rect 43346 27044 43352 27056
rect 42812 27016 43024 27044
rect 43180 27016 43352 27044
rect 38657 26979 38715 26985
rect 38657 26945 38669 26979
rect 38703 26976 38715 26979
rect 38746 26976 38752 26988
rect 38703 26948 38752 26976
rect 38703 26945 38715 26948
rect 38657 26939 38715 26945
rect 38746 26936 38752 26948
rect 38804 26936 38810 26988
rect 38838 26936 38844 26988
rect 38896 26936 38902 26988
rect 38933 26979 38991 26985
rect 38933 26945 38945 26979
rect 38979 26945 38991 26979
rect 39850 26976 39856 26988
rect 38933 26939 38991 26945
rect 39132 26948 39856 26976
rect 36909 26911 36967 26917
rect 36909 26877 36921 26911
rect 36955 26908 36967 26911
rect 37274 26908 37280 26920
rect 36955 26880 37280 26908
rect 36955 26877 36967 26880
rect 36909 26871 36967 26877
rect 37274 26868 37280 26880
rect 37332 26868 37338 26920
rect 38948 26908 38976 26939
rect 38672 26880 38976 26908
rect 38672 26852 38700 26880
rect 7423 26812 7604 26840
rect 8496 26812 10548 26840
rect 7423 26809 7435 26812
rect 7377 26803 7435 26809
rect 8496 26772 8524 26812
rect 10520 26784 10548 26812
rect 10612 26812 12434 26840
rect 38381 26843 38439 26849
rect 10612 26784 10640 26812
rect 38381 26809 38393 26843
rect 38427 26840 38439 26843
rect 38654 26840 38660 26852
rect 38427 26812 38660 26840
rect 38427 26809 38439 26812
rect 38381 26803 38439 26809
rect 38654 26800 38660 26812
rect 38712 26800 38718 26852
rect 39132 26784 39160 26948
rect 39850 26936 39856 26948
rect 39908 26936 39914 26988
rect 39942 26936 39948 26988
rect 40000 26936 40006 26988
rect 40037 26979 40095 26985
rect 40037 26945 40049 26979
rect 40083 26976 40095 26979
rect 40126 26976 40132 26988
rect 40083 26948 40132 26976
rect 40083 26945 40095 26948
rect 40037 26939 40095 26945
rect 40126 26936 40132 26948
rect 40184 26936 40190 26988
rect 42426 26976 42432 26988
rect 41984 26948 42432 26976
rect 40218 26868 40224 26920
rect 40276 26868 40282 26920
rect 7208 26744 8524 26772
rect 9950 26732 9956 26784
rect 10008 26732 10014 26784
rect 10502 26732 10508 26784
rect 10560 26732 10566 26784
rect 10594 26732 10600 26784
rect 10652 26732 10658 26784
rect 11698 26732 11704 26784
rect 11756 26732 11762 26784
rect 12529 26775 12587 26781
rect 12529 26741 12541 26775
rect 12575 26772 12587 26775
rect 13354 26772 13360 26784
rect 12575 26744 13360 26772
rect 12575 26741 12587 26744
rect 12529 26735 12587 26741
rect 13354 26732 13360 26744
rect 13412 26732 13418 26784
rect 36262 26732 36268 26784
rect 36320 26732 36326 26784
rect 36722 26732 36728 26784
rect 36780 26772 36786 26784
rect 37458 26772 37464 26784
rect 36780 26744 37464 26772
rect 36780 26732 36786 26744
rect 37458 26732 37464 26744
rect 37516 26732 37522 26784
rect 39114 26732 39120 26784
rect 39172 26732 39178 26784
rect 40678 26732 40684 26784
rect 40736 26772 40742 26784
rect 41984 26781 42012 26948
rect 42426 26936 42432 26948
rect 42484 26936 42490 26988
rect 42610 26936 42616 26988
rect 42668 26936 42674 26988
rect 42812 26985 42840 27016
rect 42797 26979 42855 26985
rect 42797 26945 42809 26979
rect 42843 26945 42855 26979
rect 42797 26939 42855 26945
rect 42981 26979 43039 26985
rect 42981 26945 42993 26979
rect 43027 26976 43039 26979
rect 43180 26976 43208 27016
rect 43346 27004 43352 27016
rect 43404 27004 43410 27056
rect 43456 27053 43484 27084
rect 46106 27072 46112 27084
rect 46164 27072 46170 27124
rect 46474 27072 46480 27124
rect 46532 27112 46538 27124
rect 46845 27115 46903 27121
rect 46845 27112 46857 27115
rect 46532 27084 46857 27112
rect 46532 27072 46538 27084
rect 46845 27081 46857 27084
rect 46891 27112 46903 27115
rect 46891 27084 48314 27112
rect 46891 27081 46903 27084
rect 46845 27075 46903 27081
rect 43441 27047 43499 27053
rect 43441 27013 43453 27047
rect 43487 27013 43499 27047
rect 43441 27007 43499 27013
rect 43530 27004 43536 27056
rect 43588 27053 43594 27056
rect 43588 27047 43617 27053
rect 43605 27013 43617 27047
rect 43588 27007 43617 27013
rect 43588 27004 43594 27007
rect 43714 27004 43720 27056
rect 43772 27004 43778 27056
rect 43809 27047 43867 27053
rect 43809 27013 43821 27047
rect 43855 27044 43867 27047
rect 43990 27044 43996 27056
rect 43855 27016 43996 27044
rect 43855 27013 43867 27016
rect 43809 27007 43867 27013
rect 43990 27004 43996 27016
rect 44048 27004 44054 27056
rect 44910 27004 44916 27056
rect 44968 27004 44974 27056
rect 45922 27004 45928 27056
rect 45980 27044 45986 27056
rect 46201 27047 46259 27053
rect 46201 27044 46213 27047
rect 45980 27016 46213 27044
rect 45980 27004 45986 27016
rect 46201 27013 46213 27016
rect 46247 27044 46259 27047
rect 47210 27044 47216 27056
rect 46247 27016 46428 27044
rect 46247 27013 46259 27016
rect 46201 27007 46259 27013
rect 43027 26948 43208 26976
rect 43027 26945 43039 26948
rect 42981 26939 43039 26945
rect 43254 26936 43260 26988
rect 43312 26936 43318 26988
rect 43732 26976 43760 27004
rect 43732 26948 43852 26976
rect 43824 26917 43852 26948
rect 43898 26936 43904 26988
rect 43956 26976 43962 26988
rect 44085 26979 44143 26985
rect 44085 26976 44097 26979
rect 43956 26948 44097 26976
rect 43956 26936 43962 26948
rect 44085 26945 44097 26948
rect 44131 26945 44143 26979
rect 44085 26939 44143 26945
rect 45738 26936 45744 26988
rect 45796 26936 45802 26988
rect 45833 26979 45891 26985
rect 45833 26945 45845 26979
rect 45879 26976 45891 26979
rect 45940 26976 45968 27004
rect 45879 26948 45968 26976
rect 45879 26945 45891 26948
rect 45833 26939 45891 26945
rect 46014 26936 46020 26988
rect 46072 26976 46078 26988
rect 46400 26985 46428 27016
rect 46483 27016 47216 27044
rect 46293 26979 46351 26985
rect 46293 26976 46305 26979
rect 46072 26948 46305 26976
rect 46072 26936 46078 26948
rect 46293 26945 46305 26948
rect 46339 26945 46351 26979
rect 46293 26939 46351 26945
rect 46385 26979 46443 26985
rect 46385 26945 46397 26979
rect 46431 26945 46443 26979
rect 46385 26939 46443 26945
rect 42889 26911 42947 26917
rect 42889 26877 42901 26911
rect 42935 26908 42947 26911
rect 43717 26911 43775 26917
rect 43717 26908 43729 26911
rect 42935 26900 43208 26908
rect 43364 26900 43729 26908
rect 42935 26880 43729 26900
rect 42935 26877 42947 26880
rect 42889 26871 42947 26877
rect 43180 26872 43392 26880
rect 43717 26877 43729 26880
rect 43763 26877 43775 26911
rect 43717 26871 43775 26877
rect 43809 26911 43867 26917
rect 43809 26877 43821 26911
rect 43855 26877 43867 26911
rect 46483 26908 46511 27016
rect 47210 27004 47216 27016
rect 47268 27004 47274 27056
rect 48286 27044 48314 27084
rect 51442 27072 51448 27124
rect 51500 27072 51506 27124
rect 51534 27072 51540 27124
rect 51592 27112 51598 27124
rect 54110 27112 54116 27124
rect 51592 27084 54116 27112
rect 51592 27072 51598 27084
rect 49970 27044 49976 27056
rect 48286 27016 49976 27044
rect 49970 27004 49976 27016
rect 50028 27004 50034 27056
rect 46566 26936 46572 26988
rect 46624 26936 46630 26988
rect 47670 26936 47676 26988
rect 47728 26976 47734 26988
rect 47949 26979 48007 26985
rect 47949 26976 47961 26979
rect 47728 26948 47961 26976
rect 47728 26936 47734 26948
rect 47949 26945 47961 26948
rect 47995 26945 48007 26979
rect 47949 26939 48007 26945
rect 48041 26979 48099 26985
rect 48041 26945 48053 26979
rect 48087 26945 48099 26979
rect 48041 26939 48099 26945
rect 43809 26871 43867 26877
rect 44100 26880 46511 26908
rect 48056 26908 48084 26939
rect 48222 26936 48228 26988
rect 48280 26936 48286 26988
rect 48774 26936 48780 26988
rect 48832 26936 48838 26988
rect 49421 26979 49479 26985
rect 49421 26945 49433 26979
rect 49467 26976 49479 26979
rect 49694 26976 49700 26988
rect 49467 26948 49700 26976
rect 49467 26945 49479 26948
rect 49421 26939 49479 26945
rect 49694 26936 49700 26948
rect 49752 26936 49758 26988
rect 50890 26936 50896 26988
rect 50948 26936 50954 26988
rect 51644 26976 51672 27084
rect 54110 27072 54116 27084
rect 54168 27072 54174 27124
rect 54570 27072 54576 27124
rect 54628 27072 54634 27124
rect 58158 27072 58164 27124
rect 58216 27072 58222 27124
rect 52178 27044 52184 27056
rect 51736 27016 52184 27044
rect 51736 26985 51764 27016
rect 52178 27004 52184 27016
rect 52236 27044 52242 27056
rect 58176 27044 58204 27072
rect 52236 27016 58204 27044
rect 52236 27004 52242 27016
rect 51184 26948 51672 26976
rect 51721 26979 51779 26985
rect 48792 26908 48820 26936
rect 48056 26880 48820 26908
rect 49789 26911 49847 26917
rect 43732 26840 43760 26871
rect 43993 26843 44051 26849
rect 43993 26840 44005 26843
rect 43732 26812 44005 26840
rect 43993 26809 44005 26812
rect 44039 26809 44051 26843
rect 43993 26803 44051 26809
rect 41969 26775 42027 26781
rect 41969 26772 41981 26775
rect 40736 26744 41981 26772
rect 40736 26732 40742 26744
rect 41969 26741 41981 26744
rect 42015 26741 42027 26775
rect 41969 26735 42027 26741
rect 42334 26732 42340 26784
rect 42392 26772 42398 26784
rect 42429 26775 42487 26781
rect 42429 26772 42441 26775
rect 42392 26744 42441 26772
rect 42392 26732 42398 26744
rect 42429 26741 42441 26744
rect 42475 26772 42487 26775
rect 44100 26772 44128 26880
rect 49789 26877 49801 26911
rect 49835 26877 49847 26911
rect 49789 26871 49847 26877
rect 45830 26800 45836 26852
rect 45888 26840 45894 26852
rect 45925 26843 45983 26849
rect 45925 26840 45937 26843
rect 45888 26812 45937 26840
rect 45888 26800 45894 26812
rect 45925 26809 45937 26812
rect 45971 26809 45983 26843
rect 45925 26803 45983 26809
rect 46014 26800 46020 26852
rect 46072 26800 46078 26852
rect 46569 26843 46627 26849
rect 46569 26809 46581 26843
rect 46615 26840 46627 26843
rect 47302 26840 47308 26852
rect 46615 26812 47308 26840
rect 46615 26809 46627 26812
rect 46569 26803 46627 26809
rect 47302 26800 47308 26812
rect 47360 26800 47366 26852
rect 49804 26840 49832 26871
rect 50154 26868 50160 26920
rect 50212 26868 50218 26920
rect 51184 26917 51212 26948
rect 51721 26945 51733 26979
rect 51767 26945 51779 26979
rect 51721 26939 51779 26945
rect 53469 26979 53527 26985
rect 53469 26945 53481 26979
rect 53515 26945 53527 26979
rect 53469 26939 53527 26945
rect 53653 26979 53711 26985
rect 53653 26945 53665 26979
rect 53699 26976 53711 26979
rect 53926 26976 53932 26988
rect 53699 26948 53932 26976
rect 53699 26945 53711 26948
rect 53653 26939 53711 26945
rect 51169 26911 51227 26917
rect 51169 26877 51181 26911
rect 51215 26877 51227 26911
rect 51169 26871 51227 26877
rect 51445 26911 51503 26917
rect 51445 26877 51457 26911
rect 51491 26908 51503 26911
rect 51626 26908 51632 26920
rect 51491 26880 51632 26908
rect 51491 26877 51503 26880
rect 51445 26871 51503 26877
rect 51626 26868 51632 26880
rect 51684 26868 51690 26920
rect 53484 26908 53512 26939
rect 53926 26936 53932 26948
rect 53984 26936 53990 26988
rect 54846 26936 54852 26988
rect 54904 26976 54910 26988
rect 56689 26979 56747 26985
rect 56689 26976 56701 26979
rect 54904 26948 56701 26976
rect 54904 26936 54910 26948
rect 56336 26920 56364 26948
rect 56689 26945 56701 26948
rect 56735 26945 56747 26979
rect 56689 26939 56747 26945
rect 56873 26979 56931 26985
rect 56873 26945 56885 26979
rect 56919 26976 56931 26979
rect 57146 26976 57152 26988
rect 56919 26948 57152 26976
rect 56919 26945 56931 26948
rect 56873 26939 56931 26945
rect 57146 26936 57152 26948
rect 57204 26976 57210 26988
rect 57885 26979 57943 26985
rect 57885 26976 57897 26979
rect 57204 26948 57897 26976
rect 57204 26936 57210 26948
rect 57885 26945 57897 26948
rect 57931 26945 57943 26979
rect 57885 26939 57943 26945
rect 54478 26908 54484 26920
rect 53484 26880 54484 26908
rect 54478 26868 54484 26880
rect 54536 26868 54542 26920
rect 56042 26868 56048 26920
rect 56100 26868 56106 26920
rect 56318 26868 56324 26920
rect 56376 26868 56382 26920
rect 56781 26911 56839 26917
rect 56781 26877 56793 26911
rect 56827 26908 56839 26911
rect 57517 26911 57575 26917
rect 57517 26908 57529 26911
rect 56827 26880 57529 26908
rect 56827 26877 56839 26880
rect 56781 26871 56839 26877
rect 57517 26877 57529 26880
rect 57563 26877 57575 26911
rect 57517 26871 57575 26877
rect 58529 26911 58587 26917
rect 58529 26877 58541 26911
rect 58575 26877 58587 26911
rect 58529 26871 58587 26877
rect 51718 26840 51724 26852
rect 48286 26812 51724 26840
rect 42475 26744 44128 26772
rect 46032 26772 46060 26800
rect 47213 26775 47271 26781
rect 47213 26772 47225 26775
rect 46032 26744 47225 26772
rect 42475 26741 42487 26744
rect 42429 26735 42487 26741
rect 47213 26741 47225 26744
rect 47259 26741 47271 26775
rect 47213 26735 47271 26741
rect 47578 26732 47584 26784
rect 47636 26772 47642 26784
rect 48286 26772 48314 26812
rect 51718 26800 51724 26812
rect 51776 26800 51782 26852
rect 53650 26840 53656 26852
rect 53300 26812 53656 26840
rect 47636 26744 48314 26772
rect 48409 26775 48467 26781
rect 47636 26732 47642 26744
rect 48409 26741 48421 26775
rect 48455 26772 48467 26775
rect 48498 26772 48504 26784
rect 48455 26744 48504 26772
rect 48455 26741 48467 26744
rect 48409 26735 48467 26741
rect 48498 26732 48504 26744
rect 48556 26732 48562 26784
rect 48774 26732 48780 26784
rect 48832 26732 48838 26784
rect 50798 26732 50804 26784
rect 50856 26732 50862 26784
rect 51626 26732 51632 26784
rect 51684 26772 51690 26784
rect 53300 26772 53328 26812
rect 53650 26800 53656 26812
rect 53708 26800 53714 26852
rect 51684 26744 53328 26772
rect 51684 26732 51690 26744
rect 53374 26732 53380 26784
rect 53432 26772 53438 26784
rect 53561 26775 53619 26781
rect 53561 26772 53573 26775
rect 53432 26744 53573 26772
rect 53432 26732 53438 26744
rect 53561 26741 53573 26744
rect 53607 26741 53619 26775
rect 53561 26735 53619 26741
rect 55398 26732 55404 26784
rect 55456 26732 55462 26784
rect 56962 26732 56968 26784
rect 57020 26732 57026 26784
rect 58544 26772 58572 26871
rect 58544 26744 58940 26772
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 5718 26528 5724 26580
rect 5776 26568 5782 26580
rect 6546 26568 6552 26580
rect 5776 26540 6552 26568
rect 5776 26528 5782 26540
rect 6546 26528 6552 26540
rect 6604 26568 6610 26580
rect 6733 26571 6791 26577
rect 6733 26568 6745 26571
rect 6604 26540 6745 26568
rect 6604 26528 6610 26540
rect 6733 26537 6745 26540
rect 6779 26537 6791 26571
rect 6733 26531 6791 26537
rect 7834 26528 7840 26580
rect 7892 26568 7898 26580
rect 7929 26571 7987 26577
rect 7929 26568 7941 26571
rect 7892 26540 7941 26568
rect 7892 26528 7898 26540
rect 7929 26537 7941 26540
rect 7975 26537 7987 26571
rect 7929 26531 7987 26537
rect 9674 26528 9680 26580
rect 9732 26568 9738 26580
rect 10045 26571 10103 26577
rect 10045 26568 10057 26571
rect 9732 26540 10057 26568
rect 9732 26528 9738 26540
rect 10045 26537 10057 26540
rect 10091 26568 10103 26571
rect 10134 26568 10140 26580
rect 10091 26540 10140 26568
rect 10091 26537 10103 26540
rect 10045 26531 10103 26537
rect 10134 26528 10140 26540
rect 10192 26528 10198 26580
rect 35345 26571 35403 26577
rect 35345 26537 35357 26571
rect 35391 26568 35403 26571
rect 40129 26571 40187 26577
rect 40129 26568 40141 26571
rect 35391 26540 40141 26568
rect 35391 26537 35403 26540
rect 35345 26531 35403 26537
rect 6086 26460 6092 26512
rect 6144 26500 6150 26512
rect 6365 26503 6423 26509
rect 6365 26500 6377 26503
rect 6144 26472 6377 26500
rect 6144 26460 6150 26472
rect 6365 26469 6377 26472
rect 6411 26500 6423 26503
rect 9214 26500 9220 26512
rect 6411 26472 9220 26500
rect 6411 26469 6423 26472
rect 6365 26463 6423 26469
rect 9214 26460 9220 26472
rect 9272 26500 9278 26512
rect 10594 26500 10600 26512
rect 9272 26472 10600 26500
rect 9272 26460 9278 26472
rect 10594 26460 10600 26472
rect 10652 26460 10658 26512
rect 12345 26503 12403 26509
rect 12345 26469 12357 26503
rect 12391 26469 12403 26503
rect 12345 26463 12403 26469
rect 3234 26392 3240 26444
rect 3292 26432 3298 26444
rect 3292 26404 4016 26432
rect 3292 26392 3298 26404
rect 3988 26376 4016 26404
rect 7098 26392 7104 26444
rect 7156 26392 7162 26444
rect 7466 26392 7472 26444
rect 7524 26432 7530 26444
rect 8205 26435 8263 26441
rect 8205 26432 8217 26435
rect 7524 26404 8217 26432
rect 7524 26392 7530 26404
rect 8205 26401 8217 26404
rect 8251 26432 8263 26435
rect 8386 26432 8392 26444
rect 8251 26404 8392 26432
rect 8251 26401 8263 26404
rect 8205 26395 8263 26401
rect 8386 26392 8392 26404
rect 8444 26392 8450 26444
rect 1394 26324 1400 26376
rect 1452 26364 1458 26376
rect 2593 26367 2651 26373
rect 2593 26364 2605 26367
rect 1452 26336 2605 26364
rect 1452 26324 1458 26336
rect 2593 26333 2605 26336
rect 2639 26364 2651 26367
rect 2869 26367 2927 26373
rect 2869 26364 2881 26367
rect 2639 26336 2881 26364
rect 2639 26333 2651 26336
rect 2593 26327 2651 26333
rect 2869 26333 2881 26336
rect 2915 26333 2927 26367
rect 2869 26327 2927 26333
rect 3513 26367 3571 26373
rect 3513 26333 3525 26367
rect 3559 26364 3571 26367
rect 3789 26367 3847 26373
rect 3789 26364 3801 26367
rect 3559 26336 3801 26364
rect 3559 26333 3571 26336
rect 3513 26327 3571 26333
rect 3789 26333 3801 26336
rect 3835 26333 3847 26367
rect 3789 26327 3847 26333
rect 3970 26324 3976 26376
rect 4028 26324 4034 26376
rect 4614 26324 4620 26376
rect 4672 26324 4678 26376
rect 4801 26367 4859 26373
rect 4801 26333 4813 26367
rect 4847 26364 4859 26367
rect 5166 26364 5172 26376
rect 4847 26336 5172 26364
rect 4847 26333 4859 26336
rect 4801 26327 4859 26333
rect 5166 26324 5172 26336
rect 5224 26324 5230 26376
rect 7116 26364 7144 26392
rect 7653 26367 7711 26373
rect 7653 26364 7665 26367
rect 7116 26336 7665 26364
rect 7653 26333 7665 26336
rect 7699 26333 7711 26367
rect 7653 26327 7711 26333
rect 10137 26367 10195 26373
rect 10137 26333 10149 26367
rect 10183 26333 10195 26367
rect 10137 26327 10195 26333
rect 1578 26256 1584 26308
rect 1636 26256 1642 26308
rect 4632 26296 4660 26324
rect 5442 26296 5448 26308
rect 4632 26268 5448 26296
rect 5442 26256 5448 26268
rect 5500 26256 5506 26308
rect 7558 26256 7564 26308
rect 7616 26296 7622 26308
rect 7929 26299 7987 26305
rect 7929 26296 7941 26299
rect 7616 26268 7941 26296
rect 7616 26256 7622 26268
rect 7929 26265 7941 26268
rect 7975 26265 7987 26299
rect 7929 26259 7987 26265
rect 10152 26240 10180 26327
rect 10962 26324 10968 26376
rect 11020 26364 11026 26376
rect 11330 26364 11336 26376
rect 11020 26336 11336 26364
rect 11020 26324 11026 26336
rect 11330 26324 11336 26336
rect 11388 26324 11394 26376
rect 12161 26367 12219 26373
rect 12161 26333 12173 26367
rect 12207 26333 12219 26367
rect 12360 26364 12388 26463
rect 35452 26444 35480 26540
rect 40129 26537 40141 26540
rect 40175 26568 40187 26571
rect 40218 26568 40224 26580
rect 40175 26540 40224 26568
rect 40175 26537 40187 26540
rect 40129 26531 40187 26537
rect 40218 26528 40224 26540
rect 40276 26528 40282 26580
rect 40586 26528 40592 26580
rect 40644 26568 40650 26580
rect 42245 26571 42303 26577
rect 42245 26568 42257 26571
rect 40644 26540 42257 26568
rect 40644 26528 40650 26540
rect 42245 26537 42257 26540
rect 42291 26537 42303 26571
rect 42245 26531 42303 26537
rect 42426 26528 42432 26580
rect 42484 26528 42490 26580
rect 42794 26528 42800 26580
rect 42852 26568 42858 26580
rect 43073 26571 43131 26577
rect 43073 26568 43085 26571
rect 42852 26540 43085 26568
rect 42852 26528 42858 26540
rect 43073 26537 43085 26540
rect 43119 26537 43131 26571
rect 43073 26531 43131 26537
rect 46201 26571 46259 26577
rect 46201 26537 46213 26571
rect 46247 26568 46259 26571
rect 46382 26568 46388 26580
rect 46247 26540 46388 26568
rect 46247 26537 46259 26540
rect 46201 26531 46259 26537
rect 46382 26528 46388 26540
rect 46440 26528 46446 26580
rect 47854 26528 47860 26580
rect 47912 26528 47918 26580
rect 48498 26577 48504 26580
rect 48488 26571 48504 26577
rect 48488 26537 48500 26571
rect 48488 26531 48504 26537
rect 48498 26528 48504 26531
rect 48556 26528 48562 26580
rect 49973 26571 50031 26577
rect 49973 26537 49985 26571
rect 50019 26568 50031 26571
rect 50154 26568 50160 26580
rect 50019 26540 50160 26568
rect 50019 26537 50031 26540
rect 49973 26531 50031 26537
rect 50154 26528 50160 26540
rect 50212 26528 50218 26580
rect 51629 26571 51687 26577
rect 51629 26568 51641 26571
rect 51046 26540 51641 26568
rect 39114 26460 39120 26512
rect 39172 26460 39178 26512
rect 39206 26460 39212 26512
rect 39264 26500 39270 26512
rect 39393 26503 39451 26509
rect 39393 26500 39405 26503
rect 39264 26472 39405 26500
rect 39264 26460 39270 26472
rect 39393 26469 39405 26472
rect 39439 26469 39451 26503
rect 39393 26463 39451 26469
rect 39942 26460 39948 26512
rect 40000 26500 40006 26512
rect 40497 26503 40555 26509
rect 40497 26500 40509 26503
rect 40000 26472 40509 26500
rect 40000 26460 40006 26472
rect 40497 26469 40509 26472
rect 40543 26469 40555 26503
rect 40497 26463 40555 26469
rect 41049 26503 41107 26509
rect 41049 26469 41061 26503
rect 41095 26500 41107 26503
rect 41690 26500 41696 26512
rect 41095 26472 41696 26500
rect 41095 26469 41107 26472
rect 41049 26463 41107 26469
rect 35434 26392 35440 26444
rect 35492 26392 35498 26444
rect 37185 26435 37243 26441
rect 37185 26401 37197 26435
rect 37231 26432 37243 26435
rect 37277 26435 37335 26441
rect 37277 26432 37289 26435
rect 37231 26404 37289 26432
rect 37231 26401 37243 26404
rect 37185 26395 37243 26401
rect 37277 26401 37289 26404
rect 37323 26401 37335 26435
rect 40310 26432 40316 26444
rect 37277 26395 37335 26401
rect 37844 26404 38516 26432
rect 37844 26376 37872 26404
rect 13642 26367 13700 26373
rect 13642 26364 13654 26367
rect 12360 26336 13654 26364
rect 12161 26327 12219 26333
rect 13642 26333 13654 26336
rect 13688 26333 13700 26367
rect 13642 26327 13700 26333
rect 13909 26367 13967 26373
rect 13909 26333 13921 26367
rect 13955 26333 13967 26367
rect 13909 26327 13967 26333
rect 10870 26256 10876 26308
rect 10928 26296 10934 26308
rect 11606 26296 11612 26308
rect 10928 26268 11612 26296
rect 10928 26256 10934 26268
rect 11606 26256 11612 26268
rect 11664 26256 11670 26308
rect 12176 26296 12204 26327
rect 12618 26296 12624 26308
rect 12176 26268 12624 26296
rect 12618 26256 12624 26268
rect 12676 26256 12682 26308
rect 13924 26296 13952 26327
rect 37826 26324 37832 26376
rect 37884 26324 37890 26376
rect 38102 26324 38108 26376
rect 38160 26364 38166 26376
rect 38488 26373 38516 26404
rect 38672 26404 40316 26432
rect 38672 26373 38700 26404
rect 40310 26392 40316 26404
rect 40368 26392 40374 26444
rect 40512 26432 40540 26463
rect 41690 26460 41696 26472
rect 41748 26460 41754 26512
rect 41208 26435 41266 26441
rect 41208 26432 41220 26435
rect 40512 26404 41220 26432
rect 41208 26401 41220 26404
rect 41254 26401 41266 26435
rect 41208 26395 41266 26401
rect 42334 26392 42340 26444
rect 42392 26392 42398 26444
rect 38197 26367 38255 26373
rect 38197 26364 38209 26367
rect 38160 26336 38209 26364
rect 38160 26324 38166 26336
rect 38197 26333 38209 26336
rect 38243 26333 38255 26367
rect 38197 26327 38255 26333
rect 38473 26367 38531 26373
rect 38473 26333 38485 26367
rect 38519 26333 38531 26367
rect 38473 26327 38531 26333
rect 38657 26367 38715 26373
rect 38657 26333 38669 26367
rect 38703 26333 38715 26367
rect 38657 26327 38715 26333
rect 38841 26367 38899 26373
rect 38841 26333 38853 26367
rect 38887 26364 38899 26367
rect 39206 26364 39212 26376
rect 38887 26336 39212 26364
rect 38887 26333 38899 26336
rect 38841 26327 38899 26333
rect 39206 26324 39212 26336
rect 39264 26324 39270 26376
rect 40402 26324 40408 26376
rect 40460 26324 40466 26376
rect 41693 26367 41751 26373
rect 41693 26333 41705 26367
rect 41739 26364 41751 26367
rect 42352 26364 42380 26392
rect 42444 26373 42472 26528
rect 51046 26512 51074 26540
rect 51629 26537 51641 26540
rect 51675 26568 51687 26571
rect 51902 26568 51908 26580
rect 51675 26540 51908 26568
rect 51675 26537 51687 26540
rect 51629 26531 51687 26537
rect 51902 26528 51908 26540
rect 51960 26528 51966 26580
rect 53742 26528 53748 26580
rect 53800 26528 53806 26580
rect 53834 26528 53840 26580
rect 53892 26568 53898 26580
rect 53929 26571 53987 26577
rect 53929 26568 53941 26571
rect 53892 26540 53941 26568
rect 53892 26528 53898 26540
rect 53929 26537 53941 26540
rect 53975 26537 53987 26571
rect 53929 26531 53987 26537
rect 54478 26528 54484 26580
rect 54536 26568 54542 26580
rect 54573 26571 54631 26577
rect 54573 26568 54585 26571
rect 54536 26540 54585 26568
rect 54536 26528 54542 26540
rect 54573 26537 54585 26540
rect 54619 26537 54631 26571
rect 54573 26531 54631 26537
rect 54754 26528 54760 26580
rect 54812 26568 54818 26580
rect 54938 26568 54944 26580
rect 54812 26540 54944 26568
rect 54812 26528 54818 26540
rect 54938 26528 54944 26540
rect 54996 26528 55002 26580
rect 56042 26528 56048 26580
rect 56100 26568 56106 26580
rect 56689 26571 56747 26577
rect 56689 26568 56701 26571
rect 56100 26540 56701 26568
rect 56100 26528 56106 26540
rect 56689 26537 56701 26540
rect 56735 26537 56747 26571
rect 56689 26531 56747 26537
rect 58161 26571 58219 26577
rect 58161 26537 58173 26571
rect 58207 26568 58219 26571
rect 58912 26568 58940 26744
rect 58207 26540 58940 26568
rect 58207 26537 58219 26540
rect 58161 26531 58219 26537
rect 44818 26460 44824 26512
rect 44876 26460 44882 26512
rect 44928 26472 46980 26500
rect 44928 26432 44956 26472
rect 45373 26435 45431 26441
rect 45373 26432 45385 26435
rect 43180 26404 44036 26432
rect 43180 26373 43208 26404
rect 44008 26376 44036 26404
rect 44652 26404 44956 26432
rect 45020 26404 45385 26432
rect 41739 26336 42380 26364
rect 42429 26367 42487 26373
rect 41739 26333 41751 26336
rect 41693 26327 41751 26333
rect 42429 26333 42441 26367
rect 42475 26333 42487 26367
rect 42429 26327 42487 26333
rect 43165 26367 43223 26373
rect 43165 26333 43177 26367
rect 43211 26333 43223 26367
rect 43165 26327 43223 26333
rect 43257 26367 43315 26373
rect 43257 26333 43269 26367
rect 43303 26364 43315 26367
rect 43898 26364 43904 26376
rect 43303 26336 43904 26364
rect 43303 26333 43315 26336
rect 43257 26327 43315 26333
rect 43898 26324 43904 26336
rect 43956 26324 43962 26376
rect 43990 26324 43996 26376
rect 44048 26324 44054 26376
rect 44450 26324 44456 26376
rect 44508 26364 44514 26376
rect 44652 26373 44680 26404
rect 45020 26373 45048 26404
rect 45373 26401 45385 26404
rect 45419 26401 45431 26435
rect 45646 26432 45652 26444
rect 45373 26395 45431 26401
rect 45572 26404 45652 26432
rect 44545 26367 44603 26373
rect 44545 26364 44557 26367
rect 44508 26336 44557 26364
rect 44508 26324 44514 26336
rect 44545 26333 44557 26336
rect 44591 26333 44603 26367
rect 44545 26327 44603 26333
rect 44637 26367 44695 26373
rect 44637 26333 44649 26367
rect 44683 26333 44695 26367
rect 44637 26327 44695 26333
rect 44821 26367 44879 26373
rect 44821 26333 44833 26367
rect 44867 26364 44879 26367
rect 45005 26367 45063 26373
rect 45005 26364 45017 26367
rect 44867 26336 45017 26364
rect 44867 26333 44879 26336
rect 44821 26327 44879 26333
rect 45005 26333 45017 26336
rect 45051 26333 45063 26367
rect 45005 26327 45063 26333
rect 45186 26324 45192 26376
rect 45244 26324 45250 26376
rect 45281 26367 45339 26373
rect 45281 26333 45293 26367
rect 45327 26364 45339 26367
rect 45477 26367 45535 26373
rect 45370 26364 45376 26366
rect 45327 26336 45376 26364
rect 45327 26333 45339 26336
rect 45281 26327 45339 26333
rect 45370 26314 45376 26336
rect 45428 26314 45434 26366
rect 45477 26333 45489 26367
rect 45523 26364 45535 26367
rect 45572 26364 45600 26404
rect 45646 26392 45652 26404
rect 45704 26432 45710 26444
rect 45704 26404 46244 26432
rect 45704 26392 45710 26404
rect 45523 26336 45600 26364
rect 46109 26367 46167 26373
rect 45523 26333 45535 26336
rect 45477 26327 45535 26333
rect 46109 26333 46121 26367
rect 46155 26333 46167 26367
rect 46216 26364 46244 26404
rect 46952 26376 46980 26472
rect 51046 26460 51080 26512
rect 51132 26460 51138 26512
rect 53650 26500 53656 26512
rect 53576 26472 53656 26500
rect 47118 26392 47124 26444
rect 47176 26432 47182 26444
rect 48225 26435 48283 26441
rect 48225 26432 48237 26435
rect 47176 26404 48237 26432
rect 47176 26392 47182 26404
rect 48225 26401 48237 26404
rect 48271 26432 48283 26435
rect 48498 26432 48504 26444
rect 48271 26404 48504 26432
rect 48271 26401 48283 26404
rect 48225 26395 48283 26401
rect 48498 26392 48504 26404
rect 48556 26432 48562 26444
rect 51046 26432 51074 26460
rect 48556 26404 51074 26432
rect 53377 26435 53435 26441
rect 48556 26392 48562 26404
rect 53377 26401 53389 26435
rect 53423 26432 53435 26435
rect 53466 26432 53472 26444
rect 53423 26404 53472 26432
rect 53423 26401 53435 26404
rect 53377 26395 53435 26401
rect 53466 26392 53472 26404
rect 53524 26392 53530 26444
rect 46293 26367 46351 26373
rect 46293 26364 46305 26367
rect 46216 26336 46305 26364
rect 46109 26327 46167 26333
rect 46293 26333 46305 26336
rect 46339 26333 46351 26367
rect 46293 26327 46351 26333
rect 14277 26299 14335 26305
rect 14277 26296 14289 26299
rect 13372 26268 14289 26296
rect 13372 26240 13400 26268
rect 14277 26265 14289 26268
rect 14323 26265 14335 26299
rect 14277 26259 14335 26265
rect 35710 26256 35716 26308
rect 35768 26256 35774 26308
rect 36722 26256 36728 26308
rect 36780 26256 36786 26308
rect 38013 26299 38071 26305
rect 38013 26296 38025 26299
rect 37568 26268 38025 26296
rect 3878 26188 3884 26240
rect 3936 26188 3942 26240
rect 4798 26188 4804 26240
rect 4856 26188 4862 26240
rect 7742 26188 7748 26240
rect 7800 26188 7806 26240
rect 10134 26188 10140 26240
rect 10192 26188 10198 26240
rect 10318 26188 10324 26240
rect 10376 26228 10382 26240
rect 12342 26228 12348 26240
rect 10376 26200 12348 26228
rect 10376 26188 10382 26200
rect 12342 26188 12348 26200
rect 12400 26228 12406 26240
rect 12529 26231 12587 26237
rect 12529 26228 12541 26231
rect 12400 26200 12541 26228
rect 12400 26188 12406 26200
rect 12529 26197 12541 26200
rect 12575 26197 12587 26231
rect 12529 26191 12587 26197
rect 13354 26188 13360 26240
rect 13412 26188 13418 26240
rect 37090 26188 37096 26240
rect 37148 26228 37154 26240
rect 37568 26228 37596 26268
rect 38013 26265 38025 26268
rect 38059 26265 38071 26299
rect 38013 26259 38071 26265
rect 38746 26256 38752 26308
rect 38804 26296 38810 26308
rect 39114 26296 39120 26308
rect 38804 26268 39120 26296
rect 38804 26256 38810 26268
rect 39114 26256 39120 26268
rect 39172 26256 39178 26308
rect 41417 26299 41475 26305
rect 41417 26265 41429 26299
rect 41463 26296 41475 26299
rect 42981 26299 43039 26305
rect 42981 26296 42993 26299
rect 41463 26268 42993 26296
rect 41463 26265 41475 26268
rect 41417 26259 41475 26265
rect 42981 26265 42993 26268
rect 43027 26296 43039 26299
rect 45097 26299 45155 26305
rect 45097 26296 45109 26299
rect 43027 26268 45109 26296
rect 43027 26265 43039 26268
rect 42981 26259 43039 26265
rect 45097 26265 45109 26268
rect 45143 26265 45155 26299
rect 45097 26259 45155 26265
rect 37148 26200 37596 26228
rect 37148 26188 37154 26200
rect 37918 26188 37924 26240
rect 37976 26188 37982 26240
rect 38838 26188 38844 26240
rect 38896 26228 38902 26240
rect 38933 26231 38991 26237
rect 38933 26228 38945 26231
rect 38896 26200 38945 26228
rect 38896 26188 38902 26200
rect 38933 26197 38945 26200
rect 38979 26228 38991 26231
rect 40770 26228 40776 26240
rect 38979 26200 40776 26228
rect 38979 26197 38991 26200
rect 38933 26191 38991 26197
rect 40770 26188 40776 26200
rect 40828 26188 40834 26240
rect 41325 26231 41383 26237
rect 41325 26197 41337 26231
rect 41371 26228 41383 26231
rect 42061 26231 42119 26237
rect 42061 26228 42073 26231
rect 41371 26200 42073 26228
rect 41371 26197 41383 26200
rect 41325 26191 41383 26197
rect 42061 26197 42073 26200
rect 42107 26228 42119 26231
rect 42150 26228 42156 26240
rect 42107 26200 42156 26228
rect 42107 26197 42119 26200
rect 42061 26191 42119 26197
rect 42150 26188 42156 26200
rect 42208 26188 42214 26240
rect 43346 26188 43352 26240
rect 43404 26228 43410 26240
rect 45738 26228 45744 26240
rect 43404 26200 45744 26228
rect 43404 26188 43410 26200
rect 45738 26188 45744 26200
rect 45796 26228 45802 26240
rect 46124 26228 46152 26327
rect 46382 26324 46388 26376
rect 46440 26324 46446 26376
rect 46934 26324 46940 26376
rect 46992 26364 46998 26376
rect 47213 26367 47271 26373
rect 47213 26364 47225 26367
rect 46992 26336 47225 26364
rect 46992 26324 46998 26336
rect 47213 26333 47225 26336
rect 47259 26333 47271 26367
rect 47213 26327 47271 26333
rect 47302 26324 47308 26376
rect 47360 26364 47366 26376
rect 47489 26367 47547 26373
rect 47489 26364 47501 26367
rect 47360 26336 47501 26364
rect 47360 26324 47366 26336
rect 47489 26333 47501 26336
rect 47535 26364 47547 26367
rect 47765 26367 47823 26373
rect 47765 26364 47777 26367
rect 47535 26336 47777 26364
rect 47535 26333 47547 26336
rect 47489 26327 47547 26333
rect 47765 26333 47777 26336
rect 47811 26333 47823 26367
rect 47765 26327 47823 26333
rect 48038 26324 48044 26376
rect 48096 26324 48102 26376
rect 51810 26324 51816 26376
rect 51868 26324 51874 26376
rect 52730 26324 52736 26376
rect 52788 26324 52794 26376
rect 46474 26256 46480 26308
rect 46532 26256 46538 26308
rect 48056 26296 48084 26324
rect 47320 26268 48084 26296
rect 46842 26228 46848 26240
rect 45796 26200 46848 26228
rect 45796 26188 45802 26200
rect 46842 26188 46848 26200
rect 46900 26188 46906 26240
rect 47320 26237 47348 26268
rect 48406 26256 48412 26308
rect 48464 26296 48470 26308
rect 48464 26268 48990 26296
rect 48464 26256 48470 26268
rect 49786 26256 49792 26308
rect 49844 26296 49850 26308
rect 50157 26299 50215 26305
rect 50157 26296 50169 26299
rect 49844 26268 50169 26296
rect 49844 26256 49850 26268
rect 50157 26265 50169 26268
rect 50203 26265 50215 26299
rect 51828 26296 51856 26324
rect 52822 26296 52828 26308
rect 51828 26268 52828 26296
rect 50157 26259 50215 26265
rect 52822 26256 52828 26268
rect 52880 26296 52886 26308
rect 53469 26299 53527 26305
rect 53469 26296 53481 26299
rect 52880 26268 53481 26296
rect 52880 26256 52886 26268
rect 53469 26265 53481 26268
rect 53515 26265 53527 26299
rect 53576 26296 53604 26472
rect 53650 26460 53656 26472
rect 53708 26460 53714 26512
rect 55306 26500 55312 26512
rect 55140 26472 55312 26500
rect 55140 26441 55168 26472
rect 55306 26460 55312 26472
rect 55364 26460 55370 26512
rect 55125 26435 55183 26441
rect 55125 26401 55137 26435
rect 55171 26401 55183 26435
rect 55125 26395 55183 26401
rect 56502 26392 56508 26444
rect 56560 26432 56566 26444
rect 56781 26435 56839 26441
rect 56781 26432 56793 26435
rect 56560 26404 56793 26432
rect 56560 26392 56566 26404
rect 56781 26401 56793 26404
rect 56827 26401 56839 26435
rect 56781 26395 56839 26401
rect 53742 26324 53748 26376
rect 53800 26324 53806 26376
rect 53834 26324 53840 26376
rect 53892 26324 53898 26376
rect 54113 26367 54171 26373
rect 54113 26333 54125 26367
rect 54159 26333 54171 26367
rect 54113 26327 54171 26333
rect 53653 26299 53711 26305
rect 53653 26296 53665 26299
rect 53576 26268 53665 26296
rect 53469 26259 53527 26265
rect 53653 26265 53665 26268
rect 53699 26265 53711 26299
rect 53653 26259 53711 26265
rect 54128 26240 54156 26327
rect 54478 26324 54484 26376
rect 54536 26324 54542 26376
rect 54570 26324 54576 26376
rect 54628 26324 54634 26376
rect 54665 26367 54723 26373
rect 54665 26333 54677 26367
rect 54711 26333 54723 26367
rect 54665 26327 54723 26333
rect 54849 26367 54907 26373
rect 54849 26333 54861 26367
rect 54895 26364 54907 26367
rect 54895 26336 55076 26364
rect 54895 26333 54907 26336
rect 54849 26327 54907 26333
rect 54202 26256 54208 26308
rect 54260 26256 54266 26308
rect 54389 26299 54447 26305
rect 54389 26265 54401 26299
rect 54435 26296 54447 26299
rect 54588 26296 54616 26324
rect 54435 26268 54616 26296
rect 54435 26265 54447 26268
rect 54389 26259 54447 26265
rect 47305 26231 47363 26237
rect 47305 26197 47317 26231
rect 47351 26197 47363 26231
rect 47305 26191 47363 26197
rect 47670 26188 47676 26240
rect 47728 26188 47734 26240
rect 53742 26188 53748 26240
rect 53800 26228 53806 26240
rect 54110 26228 54116 26240
rect 53800 26200 54116 26228
rect 53800 26188 53806 26200
rect 54110 26188 54116 26200
rect 54168 26188 54174 26240
rect 54294 26188 54300 26240
rect 54352 26188 54358 26240
rect 54680 26228 54708 26327
rect 55048 26240 55076 26336
rect 55214 26324 55220 26376
rect 55272 26364 55278 26376
rect 55309 26367 55367 26373
rect 55309 26364 55321 26367
rect 55272 26336 55321 26364
rect 55272 26324 55278 26336
rect 55309 26333 55321 26336
rect 55355 26364 55367 26367
rect 56520 26364 56548 26392
rect 55355 26336 56548 26364
rect 58437 26367 58495 26373
rect 55355 26333 55367 26336
rect 55309 26327 55367 26333
rect 58437 26333 58449 26367
rect 58483 26364 58495 26367
rect 58894 26364 58900 26376
rect 58483 26336 58900 26364
rect 58483 26333 58495 26336
rect 58437 26327 58495 26333
rect 58894 26324 58900 26336
rect 58952 26324 58958 26376
rect 57054 26305 57060 26308
rect 55125 26299 55183 26305
rect 55125 26265 55137 26299
rect 55171 26296 55183 26299
rect 55554 26299 55612 26305
rect 55554 26296 55566 26299
rect 55171 26268 55566 26296
rect 55171 26265 55183 26268
rect 55125 26259 55183 26265
rect 55554 26265 55566 26268
rect 55600 26265 55612 26299
rect 55554 26259 55612 26265
rect 57048 26259 57060 26305
rect 57054 26256 57060 26259
rect 57112 26256 57118 26308
rect 54846 26228 54852 26240
rect 54680 26200 54852 26228
rect 54846 26188 54852 26200
rect 54904 26188 54910 26240
rect 55030 26188 55036 26240
rect 55088 26188 55094 26240
rect 58250 26188 58256 26240
rect 58308 26188 58314 26240
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 1394 25984 1400 26036
rect 1452 25984 1458 26036
rect 5442 25984 5448 26036
rect 5500 25984 5506 26036
rect 7377 26027 7435 26033
rect 7377 25993 7389 26027
rect 7423 26024 7435 26027
rect 7742 26024 7748 26036
rect 7423 25996 7748 26024
rect 7423 25993 7435 25996
rect 7377 25987 7435 25993
rect 7742 25984 7748 25996
rect 7800 26024 7806 26036
rect 8297 26027 8355 26033
rect 8297 26024 8309 26027
rect 7800 25996 8309 26024
rect 7800 25984 7806 25996
rect 8297 25993 8309 25996
rect 8343 25993 8355 26027
rect 9674 26024 9680 26036
rect 8297 25987 8355 25993
rect 8588 25996 9680 26024
rect 2406 25916 2412 25968
rect 2464 25916 2470 25968
rect 7193 25959 7251 25965
rect 7193 25925 7205 25959
rect 7239 25956 7251 25959
rect 7239 25928 7880 25956
rect 7239 25925 7251 25928
rect 7193 25919 7251 25925
rect 7852 25900 7880 25928
rect 8588 25900 8616 25996
rect 9674 25984 9680 25996
rect 9732 26024 9738 26036
rect 10045 26027 10103 26033
rect 9732 25996 9996 26024
rect 9732 25984 9738 25996
rect 9766 25956 9772 25968
rect 9232 25928 9444 25956
rect 3878 25848 3884 25900
rect 3936 25848 3942 25900
rect 4332 25891 4390 25897
rect 4332 25857 4344 25891
rect 4378 25888 4390 25891
rect 4614 25888 4620 25900
rect 4378 25860 4620 25888
rect 4378 25857 4390 25860
rect 4332 25851 4390 25857
rect 4614 25848 4620 25860
rect 4672 25848 4678 25900
rect 7469 25891 7527 25897
rect 7469 25857 7481 25891
rect 7515 25857 7527 25891
rect 7469 25851 7527 25857
rect 2869 25823 2927 25829
rect 2869 25789 2881 25823
rect 2915 25820 2927 25823
rect 2915 25792 3096 25820
rect 2915 25789 2927 25792
rect 2869 25783 2927 25789
rect 3068 25752 3096 25792
rect 3142 25780 3148 25832
rect 3200 25780 3206 25832
rect 4062 25780 4068 25832
rect 4120 25780 4126 25832
rect 3418 25752 3424 25764
rect 3068 25724 3424 25752
rect 3418 25712 3424 25724
rect 3476 25712 3482 25764
rect 7484 25696 7512 25851
rect 7834 25848 7840 25900
rect 7892 25848 7898 25900
rect 8478 25848 8484 25900
rect 8536 25848 8542 25900
rect 8570 25848 8576 25900
rect 8628 25848 8634 25900
rect 8662 25848 8668 25900
rect 8720 25888 8726 25900
rect 8757 25891 8815 25897
rect 8757 25888 8769 25891
rect 8720 25860 8769 25888
rect 8720 25848 8726 25860
rect 8757 25857 8769 25860
rect 8803 25888 8815 25891
rect 9030 25888 9036 25900
rect 8803 25860 9036 25888
rect 8803 25857 8815 25860
rect 8757 25851 8815 25857
rect 9030 25848 9036 25860
rect 9088 25848 9094 25900
rect 8505 25820 8533 25848
rect 9232 25820 9260 25928
rect 9309 25891 9367 25897
rect 9309 25857 9321 25891
rect 9355 25857 9367 25891
rect 9309 25851 9367 25857
rect 8505 25792 9260 25820
rect 3234 25644 3240 25696
rect 3292 25644 3298 25696
rect 7190 25644 7196 25696
rect 7248 25644 7254 25696
rect 7466 25644 7472 25696
rect 7524 25644 7530 25696
rect 8754 25644 8760 25696
rect 8812 25644 8818 25696
rect 9122 25644 9128 25696
rect 9180 25644 9186 25696
rect 9232 25684 9260 25792
rect 9324 25752 9352 25851
rect 9416 25820 9444 25928
rect 9508 25928 9772 25956
rect 9508 25897 9536 25928
rect 9766 25916 9772 25928
rect 9824 25916 9830 25968
rect 9493 25891 9551 25897
rect 9493 25857 9505 25891
rect 9539 25857 9551 25891
rect 9493 25851 9551 25857
rect 9677 25891 9735 25897
rect 9677 25857 9689 25891
rect 9723 25857 9735 25891
rect 9968 25888 9996 25996
rect 10045 25993 10057 26027
rect 10091 26024 10103 26027
rect 10410 26024 10416 26036
rect 10091 25996 10416 26024
rect 10091 25993 10103 25996
rect 10045 25987 10103 25993
rect 10410 25984 10416 25996
rect 10468 25984 10474 26036
rect 10505 26027 10563 26033
rect 10505 25993 10517 26027
rect 10551 26024 10563 26027
rect 10870 26024 10876 26036
rect 10551 25996 10876 26024
rect 10551 25993 10563 25996
rect 10505 25987 10563 25993
rect 10870 25984 10876 25996
rect 10928 25984 10934 26036
rect 10962 25984 10968 26036
rect 11020 25984 11026 26036
rect 11514 25984 11520 26036
rect 11572 25984 11578 26036
rect 11701 26027 11759 26033
rect 11701 25993 11713 26027
rect 11747 26024 11759 26027
rect 11882 26024 11888 26036
rect 11747 25996 11888 26024
rect 11747 25993 11759 25996
rect 11701 25987 11759 25993
rect 11882 25984 11888 25996
rect 11940 26024 11946 26036
rect 12529 26027 12587 26033
rect 11940 25996 12204 26024
rect 11940 25984 11946 25996
rect 10321 25891 10379 25897
rect 10321 25888 10333 25891
rect 9968 25860 10333 25888
rect 9677 25851 9735 25857
rect 10321 25857 10333 25860
rect 10367 25857 10379 25891
rect 10321 25851 10379 25857
rect 9692 25820 9720 25851
rect 10410 25848 10416 25900
rect 10468 25888 10474 25900
rect 10505 25891 10563 25897
rect 10505 25888 10517 25891
rect 10468 25860 10517 25888
rect 10468 25848 10474 25860
rect 10505 25857 10517 25860
rect 10551 25888 10563 25891
rect 10689 25891 10747 25897
rect 10689 25888 10701 25891
rect 10551 25860 10701 25888
rect 10551 25857 10563 25860
rect 10505 25851 10563 25857
rect 10689 25857 10701 25860
rect 10735 25857 10747 25891
rect 10689 25851 10747 25857
rect 10781 25891 10839 25897
rect 10781 25857 10793 25891
rect 10827 25888 10839 25891
rect 10980 25888 11008 25984
rect 11606 25916 11612 25968
rect 11664 25956 11670 25968
rect 12176 25965 12204 25996
rect 12529 25993 12541 26027
rect 12575 26024 12587 26027
rect 12618 26024 12624 26036
rect 12575 25996 12624 26024
rect 12575 25993 12587 25996
rect 12529 25987 12587 25993
rect 12618 25984 12624 25996
rect 12676 25984 12682 26036
rect 35710 25984 35716 26036
rect 35768 25984 35774 26036
rect 36262 25984 36268 26036
rect 36320 25984 36326 26036
rect 37090 26024 37096 26036
rect 36648 25996 37096 26024
rect 11793 25959 11851 25965
rect 11793 25956 11805 25959
rect 11664 25928 11805 25956
rect 11664 25916 11670 25928
rect 11793 25925 11805 25928
rect 11839 25925 11851 25959
rect 11793 25919 11851 25925
rect 12161 25959 12219 25965
rect 12161 25925 12173 25959
rect 12207 25925 12219 25959
rect 36280 25956 36308 25984
rect 12161 25919 12219 25925
rect 12391 25925 12449 25931
rect 10827 25860 11008 25888
rect 10827 25857 10839 25860
rect 10781 25851 10839 25857
rect 9416 25792 9720 25820
rect 9769 25823 9827 25829
rect 9646 25752 9674 25792
rect 9769 25789 9781 25823
rect 9815 25820 9827 25823
rect 10796 25820 10824 25851
rect 11146 25848 11152 25900
rect 11204 25848 11210 25900
rect 11330 25848 11336 25900
rect 11388 25848 11394 25900
rect 11885 25891 11943 25897
rect 11885 25857 11897 25891
rect 11931 25888 11943 25891
rect 12066 25888 12072 25900
rect 11931 25860 12072 25888
rect 11931 25857 11943 25860
rect 11885 25851 11943 25857
rect 9815 25792 10824 25820
rect 11241 25823 11299 25829
rect 9815 25789 9827 25792
rect 9769 25783 9827 25789
rect 11241 25789 11253 25823
rect 11287 25820 11299 25823
rect 11900 25820 11928 25851
rect 12066 25848 12072 25860
rect 12124 25888 12130 25900
rect 12391 25891 12403 25925
rect 12437 25891 12449 25925
rect 35452 25928 36308 25956
rect 12391 25888 12449 25891
rect 12124 25885 12449 25888
rect 12124 25860 12434 25885
rect 12124 25848 12130 25860
rect 14918 25848 14924 25900
rect 14976 25888 14982 25900
rect 35452 25897 35480 25928
rect 36648 25897 36676 25996
rect 37090 25984 37096 25996
rect 37148 25984 37154 26036
rect 37274 25984 37280 26036
rect 37332 25984 37338 26036
rect 37826 25984 37832 26036
rect 37884 25984 37890 26036
rect 37918 25984 37924 26036
rect 37976 25984 37982 26036
rect 39114 25984 39120 26036
rect 39172 25984 39178 26036
rect 45278 25984 45284 26036
rect 45336 26024 45342 26036
rect 46014 26024 46020 26036
rect 45336 25996 46020 26024
rect 45336 25984 45342 25996
rect 46014 25984 46020 25996
rect 46072 25984 46078 26036
rect 46934 25984 46940 26036
rect 46992 25984 46998 26036
rect 47857 26027 47915 26033
rect 47857 25993 47869 26027
rect 47903 26024 47915 26027
rect 48774 26024 48780 26036
rect 47903 25996 48780 26024
rect 47903 25993 47915 25996
rect 47857 25987 47915 25993
rect 48774 25984 48780 25996
rect 48832 26024 48838 26036
rect 48832 25996 49004 26024
rect 48832 25984 48838 25996
rect 36817 25959 36875 25965
rect 36817 25925 36829 25959
rect 36863 25956 36875 25959
rect 37366 25956 37372 25968
rect 36863 25928 37372 25956
rect 36863 25925 36875 25928
rect 36817 25919 36875 25925
rect 37366 25916 37372 25928
rect 37424 25916 37430 25968
rect 37642 25956 37648 25968
rect 37476 25928 37648 25956
rect 29825 25891 29883 25897
rect 29825 25888 29837 25891
rect 14976 25860 29837 25888
rect 14976 25848 14982 25860
rect 29825 25857 29837 25860
rect 29871 25857 29883 25891
rect 29825 25851 29883 25857
rect 35437 25891 35495 25897
rect 35437 25857 35449 25891
rect 35483 25857 35495 25891
rect 35437 25851 35495 25857
rect 35621 25891 35679 25897
rect 35621 25857 35633 25891
rect 35667 25888 35679 25891
rect 36449 25891 36507 25897
rect 36449 25888 36461 25891
rect 35667 25860 36461 25888
rect 35667 25857 35679 25860
rect 35621 25851 35679 25857
rect 36449 25857 36461 25860
rect 36495 25857 36507 25891
rect 36449 25851 36507 25857
rect 36633 25891 36691 25897
rect 36633 25857 36645 25891
rect 36679 25857 36691 25891
rect 36633 25851 36691 25857
rect 36906 25848 36912 25900
rect 36964 25848 36970 25900
rect 37090 25848 37096 25900
rect 37148 25888 37154 25900
rect 37476 25897 37504 25928
rect 37642 25916 37648 25928
rect 37700 25956 37706 25968
rect 37936 25956 37964 25984
rect 38838 25956 38844 25968
rect 37700 25928 37964 25956
rect 38028 25928 38844 25956
rect 37700 25916 37706 25928
rect 37277 25891 37335 25897
rect 37277 25888 37289 25891
rect 37148 25860 37289 25888
rect 37148 25848 37154 25860
rect 37277 25857 37289 25860
rect 37323 25857 37335 25891
rect 37277 25851 37335 25857
rect 37461 25891 37519 25897
rect 37461 25857 37473 25891
rect 37507 25857 37519 25891
rect 37461 25851 37519 25857
rect 37734 25848 37740 25900
rect 37792 25848 37798 25900
rect 37921 25891 37979 25897
rect 37921 25857 37933 25891
rect 37967 25886 37979 25891
rect 38028 25886 38056 25928
rect 38838 25916 38844 25928
rect 38896 25916 38902 25968
rect 40402 25956 40408 25968
rect 39776 25928 40408 25956
rect 39209 25900 39267 25903
rect 37967 25858 38056 25886
rect 37967 25857 37979 25858
rect 37921 25851 37979 25857
rect 39206 25848 39212 25900
rect 39264 25894 39270 25900
rect 39776 25897 39804 25928
rect 40402 25916 40408 25928
rect 40460 25916 40466 25968
rect 39264 25866 39303 25894
rect 39761 25891 39819 25897
rect 39264 25848 39270 25866
rect 39761 25857 39773 25891
rect 39807 25857 39819 25891
rect 39761 25851 39819 25857
rect 39945 25891 40003 25897
rect 39945 25857 39957 25891
rect 39991 25888 40003 25891
rect 42886 25888 42892 25900
rect 39991 25860 42892 25888
rect 39991 25857 40003 25860
rect 39945 25851 40003 25857
rect 42886 25848 42892 25860
rect 42944 25848 42950 25900
rect 44450 25848 44456 25900
rect 44508 25888 44514 25900
rect 45296 25897 45324 25984
rect 45373 25959 45431 25965
rect 45373 25925 45385 25959
rect 45419 25956 45431 25959
rect 45922 25956 45928 25968
rect 45419 25928 45928 25956
rect 45419 25925 45431 25928
rect 45373 25919 45431 25925
rect 45922 25916 45928 25928
rect 45980 25956 45986 25968
rect 47765 25959 47823 25965
rect 47765 25956 47777 25959
rect 45980 25928 47777 25956
rect 45980 25916 45986 25928
rect 47765 25925 47777 25928
rect 47811 25925 47823 25959
rect 47765 25919 47823 25925
rect 47964 25928 48176 25956
rect 47964 25900 47992 25928
rect 45281 25891 45339 25897
rect 45281 25888 45293 25891
rect 44508 25860 45293 25888
rect 44508 25848 44514 25860
rect 45281 25857 45293 25860
rect 45327 25857 45339 25891
rect 45281 25851 45339 25857
rect 45465 25891 45523 25897
rect 45465 25857 45477 25891
rect 45511 25857 45523 25891
rect 45465 25851 45523 25857
rect 11287 25792 11928 25820
rect 35529 25823 35587 25829
rect 11287 25789 11299 25792
rect 11241 25783 11299 25789
rect 35529 25789 35541 25823
rect 35575 25820 35587 25823
rect 36265 25823 36323 25829
rect 36265 25820 36277 25823
rect 35575 25792 36277 25820
rect 35575 25789 35587 25792
rect 35529 25783 35587 25789
rect 36265 25789 36277 25792
rect 36311 25789 36323 25823
rect 36265 25783 36323 25789
rect 36538 25780 36544 25832
rect 36596 25820 36602 25832
rect 36596 25792 44312 25820
rect 36596 25780 36602 25792
rect 10318 25752 10324 25764
rect 9324 25724 9444 25752
rect 9646 25724 10324 25752
rect 9309 25687 9367 25693
rect 9309 25684 9321 25687
rect 9232 25656 9321 25684
rect 9309 25653 9321 25656
rect 9355 25653 9367 25687
rect 9416 25684 9444 25724
rect 10318 25712 10324 25724
rect 10376 25712 10382 25764
rect 12069 25755 12127 25761
rect 12069 25721 12081 25755
rect 12115 25752 12127 25755
rect 12158 25752 12164 25764
rect 12115 25724 12164 25752
rect 12115 25721 12127 25724
rect 12069 25715 12127 25721
rect 12158 25712 12164 25724
rect 12216 25752 12222 25764
rect 12618 25752 12624 25764
rect 12216 25724 12624 25752
rect 12216 25712 12222 25724
rect 12618 25712 12624 25724
rect 12676 25752 12682 25764
rect 13170 25752 13176 25764
rect 12676 25724 13176 25752
rect 12676 25712 12682 25724
rect 13170 25712 13176 25724
rect 13228 25712 13234 25764
rect 13446 25712 13452 25764
rect 13504 25752 13510 25764
rect 13504 25724 26234 25752
rect 13504 25712 13510 25724
rect 9861 25687 9919 25693
rect 9861 25684 9873 25687
rect 9416 25656 9873 25684
rect 9309 25647 9367 25653
rect 9861 25653 9873 25656
rect 9907 25684 9919 25687
rect 10134 25684 10140 25696
rect 9907 25656 10140 25684
rect 9907 25653 9919 25656
rect 9861 25647 9919 25653
rect 10134 25644 10140 25656
rect 10192 25684 10198 25696
rect 11146 25684 11152 25696
rect 10192 25656 11152 25684
rect 10192 25644 10198 25656
rect 11146 25644 11152 25656
rect 11204 25644 11210 25696
rect 12342 25644 12348 25696
rect 12400 25644 12406 25696
rect 26206 25684 26234 25724
rect 31110 25712 31116 25764
rect 31168 25752 31174 25764
rect 31297 25755 31355 25761
rect 31297 25752 31309 25755
rect 31168 25724 31309 25752
rect 31168 25712 31174 25724
rect 31297 25721 31309 25724
rect 31343 25752 31355 25755
rect 44082 25752 44088 25764
rect 31343 25724 44088 25752
rect 31343 25721 31355 25724
rect 31297 25715 31355 25721
rect 44082 25712 44088 25724
rect 44140 25712 44146 25764
rect 44284 25752 44312 25792
rect 45186 25780 45192 25832
rect 45244 25820 45250 25832
rect 45480 25820 45508 25851
rect 45554 25848 45560 25900
rect 45612 25888 45618 25900
rect 46753 25891 46811 25897
rect 46753 25888 46765 25891
rect 45612 25860 46765 25888
rect 45612 25848 45618 25860
rect 46753 25857 46765 25860
rect 46799 25857 46811 25891
rect 46753 25851 46811 25857
rect 46937 25891 46995 25897
rect 46937 25857 46949 25891
rect 46983 25857 46995 25891
rect 46937 25851 46995 25857
rect 46474 25820 46480 25832
rect 45244 25792 46480 25820
rect 45244 25780 45250 25792
rect 46474 25780 46480 25792
rect 46532 25780 46538 25832
rect 46290 25752 46296 25764
rect 44284 25724 46296 25752
rect 46290 25712 46296 25724
rect 46348 25712 46354 25764
rect 46952 25752 46980 25851
rect 47946 25848 47952 25900
rect 48004 25848 48010 25900
rect 48038 25848 48044 25900
rect 48096 25848 48102 25900
rect 48148 25888 48176 25928
rect 48222 25916 48228 25968
rect 48280 25916 48286 25968
rect 48406 25888 48412 25900
rect 48148 25860 48412 25888
rect 48406 25848 48412 25860
rect 48464 25888 48470 25900
rect 48501 25891 48559 25897
rect 48501 25888 48513 25891
rect 48464 25860 48513 25888
rect 48464 25848 48470 25860
rect 48501 25857 48513 25860
rect 48547 25857 48559 25891
rect 48501 25851 48559 25857
rect 47670 25780 47676 25832
rect 47728 25820 47734 25832
rect 48133 25823 48191 25829
rect 48133 25820 48145 25823
rect 47728 25792 48145 25820
rect 47728 25780 47734 25792
rect 48133 25789 48145 25792
rect 48179 25789 48191 25823
rect 48133 25783 48191 25789
rect 47854 25752 47860 25764
rect 46952 25724 47860 25752
rect 47854 25712 47860 25724
rect 47912 25712 47918 25764
rect 48976 25761 49004 25996
rect 51258 25984 51264 26036
rect 51316 25984 51322 26036
rect 52457 26027 52515 26033
rect 52457 25993 52469 26027
rect 52503 26024 52515 26027
rect 52730 26024 52736 26036
rect 52503 25996 52736 26024
rect 52503 25993 52515 25996
rect 52457 25987 52515 25993
rect 52730 25984 52736 25996
rect 52788 25984 52794 26036
rect 53466 25984 53472 26036
rect 53524 25984 53530 26036
rect 54202 25984 54208 26036
rect 54260 26024 54266 26036
rect 54665 26027 54723 26033
rect 54665 26024 54677 26027
rect 54260 25996 54677 26024
rect 54260 25984 54266 25996
rect 54665 25993 54677 25996
rect 54711 25993 54723 26027
rect 54665 25987 54723 25993
rect 55306 25984 55312 26036
rect 55364 25984 55370 26036
rect 56965 26027 57023 26033
rect 56965 25993 56977 26027
rect 57011 26024 57023 26027
rect 57054 26024 57060 26036
rect 57011 25996 57060 26024
rect 57011 25993 57023 25996
rect 56965 25987 57023 25993
rect 57054 25984 57060 25996
rect 57112 25984 57118 26036
rect 58250 25984 58256 26036
rect 58308 25984 58314 26036
rect 50798 25916 50804 25968
rect 50856 25956 50862 25968
rect 50893 25959 50951 25965
rect 50893 25956 50905 25959
rect 50856 25928 50905 25956
rect 50856 25916 50862 25928
rect 50893 25925 50905 25928
rect 50939 25925 50951 25959
rect 50893 25919 50951 25925
rect 51074 25848 51080 25900
rect 51132 25848 51138 25900
rect 51276 25888 51304 25984
rect 53484 25956 53512 25984
rect 53834 25956 53840 25968
rect 53484 25928 53840 25956
rect 51350 25897 51356 25900
rect 51184 25860 51304 25888
rect 50154 25780 50160 25832
rect 50212 25820 50218 25832
rect 51184 25820 51212 25860
rect 51344 25851 51356 25897
rect 51350 25848 51356 25851
rect 51408 25848 51414 25900
rect 52454 25848 52460 25900
rect 52512 25888 52518 25900
rect 53668 25897 53696 25928
rect 53834 25916 53840 25928
rect 53892 25916 53898 25968
rect 57974 25956 57980 25968
rect 57256 25928 57980 25956
rect 53469 25891 53527 25897
rect 53469 25888 53481 25891
rect 52512 25860 53481 25888
rect 52512 25848 52518 25860
rect 53208 25832 53236 25860
rect 53469 25857 53481 25860
rect 53515 25857 53527 25891
rect 53469 25851 53527 25857
rect 53653 25891 53711 25897
rect 53653 25857 53665 25891
rect 53699 25857 53711 25891
rect 53653 25851 53711 25857
rect 54757 25891 54815 25897
rect 54757 25857 54769 25891
rect 54803 25888 54815 25891
rect 55398 25888 55404 25900
rect 54803 25860 55404 25888
rect 54803 25857 54815 25860
rect 54757 25851 54815 25857
rect 55398 25848 55404 25860
rect 55456 25888 55462 25900
rect 56045 25891 56103 25897
rect 56045 25888 56057 25891
rect 55456 25860 56057 25888
rect 55456 25848 55462 25860
rect 56045 25857 56057 25860
rect 56091 25857 56103 25891
rect 56045 25851 56103 25857
rect 56229 25891 56287 25897
rect 56229 25857 56241 25891
rect 56275 25857 56287 25891
rect 56229 25851 56287 25857
rect 50212 25792 51212 25820
rect 50212 25780 50218 25792
rect 53190 25780 53196 25832
rect 53248 25780 53254 25832
rect 53377 25823 53435 25829
rect 53377 25789 53389 25823
rect 53423 25820 53435 25823
rect 53561 25823 53619 25829
rect 53561 25820 53573 25823
rect 53423 25792 53573 25820
rect 53423 25789 53435 25792
rect 53377 25783 53435 25789
rect 53561 25789 53573 25792
rect 53607 25789 53619 25823
rect 53561 25783 53619 25789
rect 55953 25823 56011 25829
rect 55953 25789 55965 25823
rect 55999 25820 56011 25823
rect 56137 25823 56195 25829
rect 56137 25820 56149 25823
rect 55999 25792 56149 25820
rect 55999 25789 56011 25792
rect 55953 25783 56011 25789
rect 56137 25789 56149 25792
rect 56183 25789 56195 25823
rect 56244 25820 56272 25851
rect 56778 25848 56784 25900
rect 56836 25888 56842 25900
rect 57256 25897 57284 25928
rect 57974 25916 57980 25928
rect 58032 25916 58038 25968
rect 57149 25891 57207 25897
rect 57149 25888 57161 25891
rect 56836 25860 57161 25888
rect 56836 25848 56842 25860
rect 57149 25857 57161 25860
rect 57195 25857 57207 25891
rect 57149 25851 57207 25857
rect 57241 25891 57299 25897
rect 57241 25857 57253 25891
rect 57287 25857 57299 25891
rect 57241 25851 57299 25857
rect 57885 25891 57943 25897
rect 57885 25857 57897 25891
rect 57931 25857 57943 25891
rect 57885 25851 57943 25857
rect 58161 25891 58219 25897
rect 58161 25857 58173 25891
rect 58207 25888 58219 25891
rect 58268 25888 58296 25984
rect 58207 25860 58296 25888
rect 58207 25857 58219 25860
rect 58161 25851 58219 25857
rect 56318 25820 56324 25832
rect 56244 25792 56324 25820
rect 56137 25783 56195 25789
rect 56318 25780 56324 25792
rect 56376 25820 56382 25832
rect 56502 25820 56508 25832
rect 56376 25792 56508 25820
rect 56376 25780 56382 25792
rect 56502 25780 56508 25792
rect 56560 25780 56566 25832
rect 56962 25780 56968 25832
rect 57020 25780 57026 25832
rect 57900 25820 57928 25851
rect 58618 25848 58624 25900
rect 58676 25848 58682 25900
rect 58636 25820 58664 25848
rect 57900 25792 58664 25820
rect 48961 25755 49019 25761
rect 48961 25721 48973 25755
rect 49007 25752 49019 25755
rect 49142 25752 49148 25764
rect 49007 25724 49148 25752
rect 49007 25721 49019 25724
rect 48961 25715 49019 25721
rect 49142 25712 49148 25724
rect 49200 25712 49206 25764
rect 56870 25712 56876 25764
rect 56928 25752 56934 25764
rect 58253 25755 58311 25761
rect 58253 25752 58265 25755
rect 56928 25724 58265 25752
rect 56928 25712 56934 25724
rect 58253 25721 58265 25724
rect 58299 25721 58311 25755
rect 58253 25715 58311 25721
rect 37734 25684 37740 25696
rect 26206 25656 37740 25684
rect 37734 25644 37740 25656
rect 37792 25684 37798 25696
rect 38197 25687 38255 25693
rect 38197 25684 38209 25687
rect 37792 25656 38209 25684
rect 37792 25644 37798 25656
rect 38197 25653 38209 25656
rect 38243 25653 38255 25687
rect 38197 25647 38255 25653
rect 39390 25644 39396 25696
rect 39448 25684 39454 25696
rect 39945 25687 40003 25693
rect 39945 25684 39957 25687
rect 39448 25656 39957 25684
rect 39448 25644 39454 25656
rect 39945 25653 39957 25656
rect 39991 25653 40003 25687
rect 39945 25647 40003 25653
rect 41325 25687 41383 25693
rect 41325 25653 41337 25687
rect 41371 25684 41383 25687
rect 41414 25684 41420 25696
rect 41371 25656 41420 25684
rect 41371 25653 41383 25656
rect 41325 25647 41383 25653
rect 41414 25644 41420 25656
rect 41472 25644 41478 25696
rect 41598 25644 41604 25696
rect 41656 25684 41662 25696
rect 41785 25687 41843 25693
rect 41785 25684 41797 25687
rect 41656 25656 41797 25684
rect 41656 25644 41662 25656
rect 41785 25653 41797 25656
rect 41831 25684 41843 25687
rect 42702 25684 42708 25696
rect 41831 25656 42708 25684
rect 41831 25653 41843 25656
rect 41785 25647 41843 25653
rect 42702 25644 42708 25656
rect 42760 25684 42766 25696
rect 49418 25684 49424 25696
rect 42760 25656 49424 25684
rect 42760 25644 42766 25656
rect 49418 25644 49424 25656
rect 49476 25644 49482 25696
rect 49786 25644 49792 25696
rect 49844 25644 49850 25696
rect 52730 25644 52736 25696
rect 52788 25644 52794 25696
rect 58066 25644 58072 25696
rect 58124 25644 58130 25696
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 3418 25440 3424 25492
rect 3476 25440 3482 25492
rect 3786 25440 3792 25492
rect 3844 25440 3850 25492
rect 3881 25483 3939 25489
rect 3881 25449 3893 25483
rect 3927 25480 3939 25483
rect 4062 25480 4068 25492
rect 3927 25452 4068 25480
rect 3927 25449 3939 25452
rect 3881 25443 3939 25449
rect 4062 25440 4068 25452
rect 4120 25440 4126 25492
rect 4525 25483 4583 25489
rect 4525 25449 4537 25483
rect 4571 25480 4583 25483
rect 4614 25480 4620 25492
rect 4571 25452 4620 25480
rect 4571 25449 4583 25452
rect 4525 25443 4583 25449
rect 4614 25440 4620 25452
rect 4672 25440 4678 25492
rect 5718 25440 5724 25492
rect 5776 25440 5782 25492
rect 5810 25440 5816 25492
rect 5868 25440 5874 25492
rect 7466 25440 7472 25492
rect 7524 25440 7530 25492
rect 8754 25440 8760 25492
rect 8812 25480 8818 25492
rect 9766 25480 9772 25492
rect 8812 25452 9772 25480
rect 8812 25440 8818 25452
rect 9766 25440 9772 25452
rect 9824 25480 9830 25492
rect 10137 25483 10195 25489
rect 10137 25480 10149 25483
rect 9824 25452 10149 25480
rect 9824 25440 9830 25452
rect 10137 25449 10149 25452
rect 10183 25480 10195 25483
rect 10410 25480 10416 25492
rect 10183 25452 10416 25480
rect 10183 25449 10195 25452
rect 10137 25443 10195 25449
rect 10410 25440 10416 25452
rect 10468 25440 10474 25492
rect 11793 25483 11851 25489
rect 11793 25449 11805 25483
rect 11839 25480 11851 25483
rect 11882 25480 11888 25492
rect 11839 25452 11888 25480
rect 11839 25449 11851 25452
rect 11793 25443 11851 25449
rect 11882 25440 11888 25452
rect 11940 25440 11946 25492
rect 11992 25452 12204 25480
rect 2409 25415 2467 25421
rect 2409 25381 2421 25415
rect 2455 25412 2467 25415
rect 3326 25412 3332 25424
rect 2455 25384 3332 25412
rect 2455 25381 2467 25384
rect 2409 25375 2467 25381
rect 3326 25372 3332 25384
rect 3384 25372 3390 25424
rect 2593 25347 2651 25353
rect 2593 25313 2605 25347
rect 2639 25344 2651 25347
rect 3234 25344 3240 25356
rect 2639 25316 3240 25344
rect 2639 25313 2651 25316
rect 2593 25307 2651 25313
rect 3234 25304 3240 25316
rect 3292 25304 3298 25356
rect 3694 25304 3700 25356
rect 3752 25304 3758 25356
rect 3804 25344 3832 25440
rect 5537 25347 5595 25353
rect 3804 25316 4108 25344
rect 2317 25279 2375 25285
rect 2317 25245 2329 25279
rect 2363 25245 2375 25279
rect 2777 25279 2835 25285
rect 2777 25276 2789 25279
rect 2317 25239 2375 25245
rect 2608 25248 2789 25276
rect 2332 25140 2360 25239
rect 2608 25217 2636 25248
rect 2777 25245 2789 25248
rect 2823 25245 2835 25279
rect 3712 25276 3740 25304
rect 4080 25288 4108 25316
rect 4264 25316 5497 25344
rect 3789 25279 3847 25285
rect 3789 25276 3801 25279
rect 3712 25248 3801 25276
rect 2777 25239 2835 25245
rect 3789 25245 3801 25248
rect 3835 25245 3847 25279
rect 3789 25239 3847 25245
rect 4062 25236 4068 25288
rect 4120 25236 4126 25288
rect 4264 25285 4292 25316
rect 4249 25279 4307 25285
rect 4249 25245 4261 25279
rect 4295 25245 4307 25279
rect 4706 25276 4712 25288
rect 4249 25239 4307 25245
rect 4540 25248 4712 25276
rect 4540 25217 4568 25248
rect 4706 25236 4712 25248
rect 4764 25236 4770 25288
rect 4798 25236 4804 25288
rect 4856 25236 4862 25288
rect 5166 25236 5172 25288
rect 5224 25276 5230 25288
rect 5261 25279 5319 25285
rect 5261 25276 5273 25279
rect 5224 25248 5273 25276
rect 5224 25236 5230 25248
rect 5261 25245 5273 25248
rect 5307 25245 5319 25279
rect 5469 25276 5497 25316
rect 5537 25313 5549 25347
rect 5583 25344 5595 25347
rect 5828 25344 5856 25440
rect 5905 25415 5963 25421
rect 5905 25381 5917 25415
rect 5951 25381 5963 25415
rect 5905 25375 5963 25381
rect 5583 25316 5856 25344
rect 5583 25313 5595 25316
rect 5537 25307 5595 25313
rect 5626 25276 5632 25288
rect 5469 25248 5632 25276
rect 5261 25239 5319 25245
rect 2593 25211 2651 25217
rect 2593 25177 2605 25211
rect 2639 25177 2651 25211
rect 4525 25211 4583 25217
rect 2593 25171 2651 25177
rect 2746 25180 4108 25208
rect 2746 25140 2774 25180
rect 4080 25149 4108 25180
rect 4525 25177 4537 25211
rect 4571 25177 4583 25211
rect 4525 25171 4583 25177
rect 5077 25211 5135 25217
rect 5077 25177 5089 25211
rect 5123 25177 5135 25211
rect 5276 25208 5304 25239
rect 5626 25236 5632 25248
rect 5684 25236 5690 25288
rect 5813 25279 5871 25285
rect 5813 25245 5825 25279
rect 5859 25276 5871 25279
rect 5920 25276 5948 25375
rect 7282 25372 7288 25424
rect 7340 25372 7346 25424
rect 9122 25372 9128 25424
rect 9180 25372 9186 25424
rect 11146 25372 11152 25424
rect 11204 25412 11210 25424
rect 11992 25412 12020 25452
rect 11204 25384 12020 25412
rect 12176 25412 12204 25452
rect 12526 25440 12532 25492
rect 12584 25480 12590 25492
rect 13078 25480 13084 25492
rect 12584 25452 13084 25480
rect 12584 25440 12590 25452
rect 13078 25440 13084 25452
rect 13136 25480 13142 25492
rect 13630 25480 13636 25492
rect 13136 25452 13636 25480
rect 13136 25440 13142 25452
rect 13630 25440 13636 25452
rect 13688 25480 13694 25492
rect 13817 25483 13875 25489
rect 13817 25480 13829 25483
rect 13688 25452 13829 25480
rect 13688 25440 13694 25452
rect 13817 25449 13829 25452
rect 13863 25449 13875 25483
rect 13817 25443 13875 25449
rect 25314 25440 25320 25492
rect 25372 25480 25378 25492
rect 36538 25480 36544 25492
rect 25372 25452 26234 25480
rect 25372 25440 25378 25452
rect 26206 25412 26234 25452
rect 31726 25452 36544 25480
rect 31726 25412 31754 25452
rect 36538 25440 36544 25452
rect 36596 25440 36602 25492
rect 36906 25440 36912 25492
rect 36964 25480 36970 25492
rect 37093 25483 37151 25489
rect 37093 25480 37105 25483
rect 36964 25452 37105 25480
rect 36964 25440 36970 25452
rect 37093 25449 37105 25452
rect 37139 25449 37151 25483
rect 37093 25443 37151 25449
rect 37458 25440 37464 25492
rect 37516 25480 37522 25492
rect 38013 25483 38071 25489
rect 38013 25480 38025 25483
rect 37516 25452 38025 25480
rect 37516 25440 37522 25452
rect 38013 25449 38025 25452
rect 38059 25480 38071 25483
rect 38562 25480 38568 25492
rect 38059 25452 38568 25480
rect 38059 25449 38071 25452
rect 38013 25443 38071 25449
rect 38562 25440 38568 25452
rect 38620 25440 38626 25492
rect 39669 25483 39727 25489
rect 39669 25449 39681 25483
rect 39715 25480 39727 25483
rect 40402 25480 40408 25492
rect 39715 25452 40408 25480
rect 39715 25449 39727 25452
rect 39669 25443 39727 25449
rect 40402 25440 40408 25452
rect 40460 25440 40466 25492
rect 40957 25483 41015 25489
rect 40957 25480 40969 25483
rect 40512 25452 40969 25480
rect 37642 25412 37648 25424
rect 12176 25384 13124 25412
rect 26206 25384 31754 25412
rect 37016 25384 37648 25412
rect 11204 25372 11210 25384
rect 7300 25344 7328 25372
rect 7300 25316 7604 25344
rect 5859 25248 5948 25276
rect 7029 25279 7087 25285
rect 5859 25245 5871 25248
rect 5813 25239 5871 25245
rect 7029 25245 7041 25279
rect 7075 25276 7087 25279
rect 7190 25276 7196 25288
rect 7075 25248 7196 25276
rect 7075 25245 7087 25248
rect 7029 25239 7087 25245
rect 5828 25208 5856 25239
rect 7190 25236 7196 25248
rect 7248 25236 7254 25288
rect 7282 25236 7288 25288
rect 7340 25236 7346 25288
rect 7576 25285 7604 25316
rect 8570 25304 8576 25356
rect 8628 25304 8634 25356
rect 7377 25279 7435 25285
rect 7377 25245 7389 25279
rect 7423 25245 7435 25279
rect 7377 25239 7435 25245
rect 7561 25279 7619 25285
rect 7561 25245 7573 25279
rect 7607 25276 7619 25279
rect 7926 25276 7932 25288
rect 7607 25248 7932 25276
rect 7607 25245 7619 25248
rect 7561 25239 7619 25245
rect 7392 25208 7420 25239
rect 7926 25236 7932 25248
rect 7984 25236 7990 25288
rect 8478 25236 8484 25288
rect 8536 25276 8542 25288
rect 9140 25276 9168 25372
rect 9674 25304 9680 25356
rect 9732 25344 9738 25356
rect 9953 25347 10011 25353
rect 9953 25344 9965 25347
rect 9732 25316 9965 25344
rect 9732 25304 9738 25316
rect 9953 25313 9965 25316
rect 9999 25313 10011 25347
rect 9953 25307 10011 25313
rect 10152 25316 12020 25344
rect 10152 25285 10180 25316
rect 11992 25285 12020 25316
rect 12066 25304 12072 25356
rect 12124 25344 12130 25356
rect 12124 25316 12204 25344
rect 12124 25304 12130 25316
rect 12176 25285 12204 25316
rect 13096 25288 13124 25384
rect 9309 25279 9367 25285
rect 9309 25276 9321 25279
rect 8536 25248 9076 25276
rect 9140 25248 9321 25276
rect 8536 25236 8542 25248
rect 8018 25208 8024 25220
rect 5276 25180 5764 25208
rect 5828 25180 7420 25208
rect 7484 25180 8024 25208
rect 5077 25171 5135 25177
rect 2332 25112 2774 25140
rect 4065 25143 4123 25149
rect 4065 25109 4077 25143
rect 4111 25109 4123 25143
rect 4065 25103 4123 25109
rect 4706 25100 4712 25152
rect 4764 25140 4770 25152
rect 4893 25143 4951 25149
rect 4893 25140 4905 25143
rect 4764 25112 4905 25140
rect 4764 25100 4770 25112
rect 4893 25109 4905 25112
rect 4939 25109 4951 25143
rect 5092 25140 5120 25171
rect 5442 25140 5448 25152
rect 5092 25112 5448 25140
rect 4893 25103 4951 25109
rect 5442 25100 5448 25112
rect 5500 25100 5506 25152
rect 5534 25100 5540 25152
rect 5592 25100 5598 25152
rect 5736 25140 5764 25180
rect 7484 25140 7512 25180
rect 8018 25168 8024 25180
rect 8076 25208 8082 25220
rect 8757 25211 8815 25217
rect 8076 25180 8432 25208
rect 8076 25168 8082 25180
rect 5736 25112 7512 25140
rect 8294 25100 8300 25152
rect 8352 25100 8358 25152
rect 8404 25140 8432 25180
rect 8757 25177 8769 25211
rect 8803 25208 8815 25211
rect 8846 25208 8852 25220
rect 8803 25180 8852 25208
rect 8803 25177 8815 25180
rect 8757 25171 8815 25177
rect 8846 25168 8852 25180
rect 8904 25168 8910 25220
rect 9048 25208 9076 25248
rect 9309 25245 9321 25248
rect 9355 25245 9367 25279
rect 10137 25279 10195 25285
rect 10137 25276 10149 25279
rect 9309 25239 9367 25245
rect 9646 25248 10149 25276
rect 9646 25208 9674 25248
rect 10137 25245 10149 25248
rect 10183 25245 10195 25279
rect 10137 25239 10195 25245
rect 11885 25279 11943 25285
rect 11885 25245 11897 25279
rect 11931 25245 11943 25279
rect 11885 25239 11943 25245
rect 11977 25279 12035 25285
rect 11977 25245 11989 25279
rect 12023 25245 12035 25279
rect 11977 25239 12035 25245
rect 12161 25279 12219 25285
rect 12161 25245 12173 25279
rect 12207 25245 12219 25279
rect 12161 25239 12219 25245
rect 12897 25279 12955 25285
rect 12897 25245 12909 25279
rect 12943 25245 12955 25279
rect 12897 25239 12955 25245
rect 9048 25180 9674 25208
rect 9858 25168 9864 25220
rect 9916 25208 9922 25220
rect 10226 25208 10232 25220
rect 9916 25180 10232 25208
rect 9916 25168 9922 25180
rect 10226 25168 10232 25180
rect 10284 25168 10290 25220
rect 9033 25143 9091 25149
rect 9033 25140 9045 25143
rect 8404 25112 9045 25140
rect 9033 25109 9045 25112
rect 9079 25109 9091 25143
rect 9033 25103 9091 25109
rect 10318 25100 10324 25152
rect 10376 25100 10382 25152
rect 11900 25140 11928 25239
rect 12069 25211 12127 25217
rect 12069 25177 12081 25211
rect 12115 25208 12127 25211
rect 12710 25208 12716 25220
rect 12115 25180 12716 25208
rect 12115 25177 12127 25180
rect 12069 25171 12127 25177
rect 12710 25168 12716 25180
rect 12768 25208 12774 25220
rect 12912 25208 12940 25239
rect 13078 25236 13084 25288
rect 13136 25236 13142 25288
rect 13357 25279 13415 25285
rect 13357 25276 13369 25279
rect 13280 25248 13369 25276
rect 12768 25180 12940 25208
rect 12768 25168 12774 25180
rect 12526 25140 12532 25152
rect 11900 25112 12532 25140
rect 12526 25100 12532 25112
rect 12584 25100 12590 25152
rect 13280 25149 13308 25248
rect 13357 25245 13369 25248
rect 13403 25245 13415 25279
rect 13357 25239 13415 25245
rect 36814 25236 36820 25288
rect 36872 25236 36878 25288
rect 37016 25285 37044 25384
rect 37642 25372 37648 25384
rect 37700 25372 37706 25424
rect 40313 25415 40371 25421
rect 40313 25381 40325 25415
rect 40359 25412 40371 25415
rect 40512 25412 40540 25452
rect 40957 25449 40969 25452
rect 41003 25480 41015 25483
rect 41414 25480 41420 25492
rect 41003 25452 41420 25480
rect 41003 25449 41015 25452
rect 40957 25443 41015 25449
rect 41414 25440 41420 25452
rect 41472 25480 41478 25492
rect 42242 25480 42248 25492
rect 41472 25452 42248 25480
rect 41472 25440 41478 25452
rect 42242 25440 42248 25452
rect 42300 25440 42306 25492
rect 42610 25440 42616 25492
rect 42668 25480 42674 25492
rect 42668 25452 44036 25480
rect 42668 25440 42674 25452
rect 40359 25384 40540 25412
rect 40359 25381 40371 25384
rect 40313 25375 40371 25381
rect 40328 25344 40356 25375
rect 40770 25372 40776 25424
rect 40828 25412 40834 25424
rect 41506 25412 41512 25424
rect 40828 25384 41512 25412
rect 40828 25372 40834 25384
rect 41506 25372 41512 25384
rect 41564 25372 41570 25424
rect 44008 25412 44036 25452
rect 44082 25440 44088 25492
rect 44140 25480 44146 25492
rect 44637 25483 44695 25489
rect 44637 25480 44649 25483
rect 44140 25452 44649 25480
rect 44140 25440 44146 25452
rect 44637 25449 44649 25452
rect 44683 25480 44695 25483
rect 47302 25480 47308 25492
rect 44683 25452 47308 25480
rect 44683 25449 44695 25452
rect 44637 25443 44695 25449
rect 47302 25440 47308 25452
rect 47360 25480 47366 25492
rect 47946 25480 47952 25492
rect 47360 25452 47952 25480
rect 47360 25440 47366 25452
rect 47946 25440 47952 25452
rect 48004 25440 48010 25492
rect 48041 25483 48099 25489
rect 48041 25449 48053 25483
rect 48087 25480 48099 25483
rect 48130 25480 48136 25492
rect 48087 25452 48136 25480
rect 48087 25449 48099 25452
rect 48041 25443 48099 25449
rect 48130 25440 48136 25452
rect 48188 25440 48194 25492
rect 48406 25440 48412 25492
rect 48464 25480 48470 25492
rect 48501 25483 48559 25489
rect 48501 25480 48513 25483
rect 48464 25452 48513 25480
rect 48464 25440 48470 25452
rect 48501 25449 48513 25452
rect 48547 25449 48559 25483
rect 48501 25443 48559 25449
rect 51350 25440 51356 25492
rect 51408 25440 51414 25492
rect 51445 25483 51503 25489
rect 51445 25449 51457 25483
rect 51491 25480 51503 25483
rect 51626 25480 51632 25492
rect 51491 25452 51632 25480
rect 51491 25449 51503 25452
rect 51445 25443 51503 25449
rect 51626 25440 51632 25452
rect 51684 25440 51690 25492
rect 52730 25440 52736 25492
rect 52788 25440 52794 25492
rect 53098 25440 53104 25492
rect 53156 25480 53162 25492
rect 53742 25480 53748 25492
rect 53156 25452 53748 25480
rect 53156 25440 53162 25452
rect 53742 25440 53748 25452
rect 53800 25440 53806 25492
rect 44269 25415 44327 25421
rect 44269 25412 44281 25415
rect 44008 25384 44281 25412
rect 44269 25381 44281 25384
rect 44315 25381 44327 25415
rect 49418 25412 49424 25424
rect 44269 25375 44327 25381
rect 46676 25384 49424 25412
rect 37200 25316 37964 25344
rect 37001 25279 37059 25285
rect 37001 25245 37013 25279
rect 37047 25245 37059 25279
rect 37001 25239 37059 25245
rect 36909 25211 36967 25217
rect 36909 25177 36921 25211
rect 36955 25208 36967 25211
rect 37200 25208 37228 25316
rect 37277 25279 37335 25285
rect 37277 25245 37289 25279
rect 37323 25245 37335 25279
rect 37277 25239 37335 25245
rect 36955 25180 37228 25208
rect 36955 25177 36967 25180
rect 36909 25171 36967 25177
rect 13265 25143 13323 25149
rect 13265 25109 13277 25143
rect 13311 25109 13323 25143
rect 13265 25103 13323 25109
rect 13446 25100 13452 25152
rect 13504 25100 13510 25152
rect 37292 25140 37320 25239
rect 37458 25236 37464 25288
rect 37516 25236 37522 25288
rect 37553 25279 37611 25285
rect 37553 25245 37565 25279
rect 37599 25245 37611 25279
rect 37553 25239 37611 25245
rect 37568 25208 37596 25239
rect 37642 25236 37648 25288
rect 37700 25236 37706 25288
rect 37826 25236 37832 25288
rect 37884 25236 37890 25288
rect 37936 25285 37964 25316
rect 38764 25316 40356 25344
rect 38764 25285 38792 25316
rect 37921 25279 37979 25285
rect 37921 25245 37933 25279
rect 37967 25245 37979 25279
rect 37921 25239 37979 25245
rect 38749 25279 38807 25285
rect 38749 25245 38761 25279
rect 38795 25245 38807 25279
rect 38749 25239 38807 25245
rect 38930 25236 38936 25288
rect 38988 25236 38994 25288
rect 39500 25285 39528 25316
rect 40586 25304 40592 25356
rect 40644 25304 40650 25356
rect 40696 25316 42196 25344
rect 39301 25279 39359 25285
rect 39301 25245 39313 25279
rect 39347 25276 39359 25279
rect 39485 25279 39543 25285
rect 39485 25276 39497 25279
rect 39347 25248 39497 25276
rect 39347 25245 39359 25248
rect 39301 25239 39359 25245
rect 39485 25245 39497 25248
rect 39531 25245 39543 25279
rect 39485 25239 39543 25245
rect 39669 25279 39727 25285
rect 39669 25245 39681 25279
rect 39715 25245 39727 25279
rect 39669 25239 39727 25245
rect 37737 25211 37795 25217
rect 37737 25208 37749 25211
rect 37568 25180 37749 25208
rect 37737 25177 37749 25180
rect 37783 25177 37795 25211
rect 39684 25208 39712 25239
rect 40034 25236 40040 25288
rect 40092 25276 40098 25288
rect 40604 25276 40632 25304
rect 40092 25248 40632 25276
rect 40092 25236 40098 25248
rect 39945 25211 40003 25217
rect 39945 25208 39957 25211
rect 37737 25171 37795 25177
rect 38856 25180 39957 25208
rect 38856 25140 38884 25180
rect 39945 25177 39957 25180
rect 39991 25177 40003 25211
rect 39945 25171 40003 25177
rect 37292 25112 38884 25140
rect 38933 25143 38991 25149
rect 38933 25109 38945 25143
rect 38979 25140 38991 25143
rect 39206 25140 39212 25152
rect 38979 25112 39212 25140
rect 38979 25109 38991 25112
rect 38933 25103 38991 25109
rect 39206 25100 39212 25112
rect 39264 25140 39270 25152
rect 40696 25140 40724 25316
rect 41598 25236 41604 25288
rect 41656 25236 41662 25288
rect 41690 25236 41696 25288
rect 41748 25236 41754 25288
rect 41874 25236 41880 25288
rect 41932 25236 41938 25288
rect 42168 25285 42196 25316
rect 42518 25304 42524 25356
rect 42576 25304 42582 25356
rect 42153 25279 42211 25285
rect 42153 25245 42165 25279
rect 42199 25245 42211 25279
rect 44082 25276 44088 25288
rect 43930 25248 44088 25276
rect 42153 25239 42211 25245
rect 44082 25236 44088 25248
rect 44140 25236 44146 25288
rect 41046 25168 41052 25220
rect 41104 25208 41110 25220
rect 41141 25211 41199 25217
rect 41141 25208 41153 25211
rect 41104 25180 41153 25208
rect 41104 25168 41110 25180
rect 41141 25177 41153 25180
rect 41187 25208 41199 25211
rect 41233 25211 41291 25217
rect 41233 25208 41245 25211
rect 41187 25180 41245 25208
rect 41187 25177 41199 25180
rect 41141 25171 41199 25177
rect 41233 25177 41245 25180
rect 41279 25177 41291 25211
rect 41233 25171 41291 25177
rect 41449 25211 41507 25217
rect 41449 25177 41461 25211
rect 41495 25208 41507 25211
rect 41616 25208 41644 25236
rect 41495 25180 41644 25208
rect 41495 25177 41507 25180
rect 41449 25171 41507 25177
rect 41782 25168 41788 25220
rect 41840 25168 41846 25220
rect 42794 25168 42800 25220
rect 42852 25168 42858 25220
rect 44284 25208 44312 25375
rect 45649 25347 45707 25353
rect 45649 25313 45661 25347
rect 45695 25344 45707 25347
rect 46477 25347 46535 25353
rect 46477 25344 46489 25347
rect 45695 25316 46489 25344
rect 45695 25313 45707 25316
rect 45649 25307 45707 25313
rect 46477 25313 46489 25316
rect 46523 25313 46535 25347
rect 46477 25307 46535 25313
rect 44818 25236 44824 25288
rect 44876 25276 44882 25288
rect 45278 25276 45284 25288
rect 44876 25248 45284 25276
rect 44876 25236 44882 25248
rect 45278 25236 45284 25248
rect 45336 25276 45342 25288
rect 45741 25279 45799 25285
rect 45741 25276 45753 25279
rect 45336 25248 45753 25276
rect 45336 25236 45342 25248
rect 45741 25245 45753 25248
rect 45787 25245 45799 25279
rect 45741 25239 45799 25245
rect 45922 25236 45928 25288
rect 45980 25236 45986 25288
rect 46014 25236 46020 25288
rect 46072 25236 46078 25288
rect 46109 25279 46167 25285
rect 46109 25245 46121 25279
rect 46155 25245 46167 25279
rect 46109 25239 46167 25245
rect 44284 25180 45508 25208
rect 40954 25149 40960 25152
rect 39264 25112 40724 25140
rect 40941 25143 40960 25149
rect 39264 25100 39270 25112
rect 40941 25109 40953 25143
rect 40941 25103 40960 25109
rect 40954 25100 40960 25103
rect 41012 25100 41018 25152
rect 41601 25143 41659 25149
rect 41601 25109 41613 25143
rect 41647 25140 41659 25143
rect 42886 25140 42892 25152
rect 41647 25112 42892 25140
rect 41647 25109 41659 25112
rect 41601 25103 41659 25109
rect 42886 25100 42892 25112
rect 42944 25100 42950 25152
rect 45002 25100 45008 25152
rect 45060 25100 45066 25152
rect 45480 25140 45508 25180
rect 45554 25168 45560 25220
rect 45612 25208 45618 25220
rect 46124 25208 46152 25239
rect 46290 25236 46296 25288
rect 46348 25276 46354 25288
rect 46676 25285 46704 25384
rect 49418 25372 49424 25384
rect 49476 25372 49482 25424
rect 46842 25304 46848 25356
rect 46900 25304 46906 25356
rect 46943 25353 46949 25356
rect 46937 25307 46949 25353
rect 47001 25344 47007 25356
rect 51261 25347 51319 25353
rect 47001 25316 47037 25344
rect 47136 25316 47992 25344
rect 46943 25304 46949 25307
rect 47001 25304 47007 25316
rect 46661 25279 46719 25285
rect 46661 25276 46673 25279
rect 46348 25248 46673 25276
rect 46348 25236 46354 25248
rect 46661 25245 46673 25248
rect 46707 25245 46719 25279
rect 46661 25239 46719 25245
rect 46753 25279 46811 25285
rect 46753 25245 46765 25279
rect 46799 25245 46811 25279
rect 46860 25276 46888 25304
rect 47136 25285 47164 25316
rect 47964 25285 47992 25316
rect 51261 25313 51273 25347
rect 51307 25344 51319 25347
rect 52748 25344 52776 25440
rect 54846 25412 54852 25424
rect 51307 25316 52776 25344
rect 53116 25384 54852 25412
rect 51307 25313 51319 25316
rect 51261 25307 51319 25313
rect 47121 25279 47179 25285
rect 47121 25276 47133 25279
rect 46860 25248 47133 25276
rect 46753 25239 46811 25245
rect 47121 25245 47133 25248
rect 47167 25245 47179 25279
rect 47121 25239 47179 25245
rect 47305 25279 47363 25285
rect 47305 25245 47317 25279
rect 47351 25276 47363 25279
rect 47949 25279 48007 25285
rect 47351 25248 47440 25276
rect 47351 25245 47363 25248
rect 47305 25239 47363 25245
rect 46768 25208 46796 25239
rect 47026 25208 47032 25220
rect 45612 25180 46511 25208
rect 46768 25180 47032 25208
rect 45612 25168 45618 25180
rect 46198 25140 46204 25152
rect 45480 25112 46204 25140
rect 46198 25100 46204 25112
rect 46256 25100 46262 25152
rect 46382 25100 46388 25152
rect 46440 25100 46446 25152
rect 46483 25140 46511 25180
rect 47026 25168 47032 25180
rect 47084 25168 47090 25220
rect 47412 25152 47440 25248
rect 47949 25245 47961 25279
rect 47995 25245 48007 25279
rect 47949 25239 48007 25245
rect 48866 25236 48872 25288
rect 48924 25276 48930 25288
rect 49237 25279 49295 25285
rect 49237 25276 49249 25279
rect 48924 25248 49249 25276
rect 48924 25236 48930 25248
rect 49237 25245 49249 25248
rect 49283 25245 49295 25279
rect 49237 25239 49295 25245
rect 51537 25279 51595 25285
rect 51537 25245 51549 25279
rect 51583 25276 51595 25279
rect 53116 25276 53144 25384
rect 54846 25372 54852 25384
rect 54904 25412 54910 25424
rect 58253 25415 58311 25421
rect 58253 25412 58265 25415
rect 54904 25384 58265 25412
rect 54904 25372 54910 25384
rect 58253 25381 58265 25384
rect 58299 25381 58311 25415
rect 58253 25375 58311 25381
rect 53285 25347 53343 25353
rect 53285 25313 53297 25347
rect 53331 25344 53343 25347
rect 53837 25347 53895 25353
rect 53837 25344 53849 25347
rect 53331 25316 53512 25344
rect 53331 25313 53343 25316
rect 53285 25307 53343 25313
rect 51583 25248 53144 25276
rect 53193 25279 53251 25285
rect 51583 25245 51595 25248
rect 51537 25239 51595 25245
rect 53193 25245 53205 25279
rect 53239 25245 53251 25279
rect 53193 25239 53251 25245
rect 53208 25208 53236 25239
rect 53374 25236 53380 25288
rect 53432 25236 53438 25288
rect 53484 25285 53512 25316
rect 53668 25316 53849 25344
rect 53668 25285 53696 25316
rect 53837 25313 53849 25316
rect 53883 25313 53895 25347
rect 53837 25307 53895 25313
rect 54478 25304 54484 25356
rect 54536 25344 54542 25356
rect 54938 25344 54944 25356
rect 54536 25316 54944 25344
rect 54536 25304 54542 25316
rect 53469 25279 53527 25285
rect 53469 25245 53481 25279
rect 53515 25245 53527 25279
rect 53469 25239 53527 25245
rect 53653 25279 53711 25285
rect 53653 25245 53665 25279
rect 53699 25245 53711 25279
rect 53653 25239 53711 25245
rect 53742 25236 53748 25288
rect 53800 25236 53806 25288
rect 53929 25279 53987 25285
rect 53929 25245 53941 25279
rect 53975 25245 53987 25279
rect 53929 25239 53987 25245
rect 54205 25279 54263 25285
rect 54205 25245 54217 25279
rect 54251 25276 54263 25279
rect 54294 25276 54300 25288
rect 54251 25248 54300 25276
rect 54251 25245 54263 25248
rect 54205 25239 54263 25245
rect 53834 25208 53840 25220
rect 53024 25180 53840 25208
rect 47213 25143 47271 25149
rect 47213 25140 47225 25143
rect 46483 25112 47225 25140
rect 47213 25109 47225 25112
rect 47259 25109 47271 25143
rect 47213 25103 47271 25109
rect 47394 25100 47400 25152
rect 47452 25100 47458 25152
rect 48590 25100 48596 25152
rect 48648 25140 48654 25152
rect 48685 25143 48743 25149
rect 48685 25140 48697 25143
rect 48648 25112 48697 25140
rect 48648 25100 48654 25112
rect 48685 25109 48697 25112
rect 48731 25109 48743 25143
rect 48685 25103 48743 25109
rect 49142 25100 49148 25152
rect 49200 25140 49206 25152
rect 53024 25149 53052 25180
rect 53834 25168 53840 25180
rect 53892 25168 53898 25220
rect 53944 25208 53972 25239
rect 54294 25236 54300 25248
rect 54352 25236 54358 25288
rect 54588 25285 54616 25316
rect 54938 25304 54944 25316
rect 54996 25344 55002 25356
rect 57425 25347 57483 25353
rect 54996 25316 57368 25344
rect 54996 25304 55002 25316
rect 54389 25279 54447 25285
rect 54389 25245 54401 25279
rect 54435 25245 54447 25279
rect 54389 25239 54447 25245
rect 54573 25279 54631 25285
rect 54573 25245 54585 25279
rect 54619 25245 54631 25279
rect 54573 25239 54631 25245
rect 54757 25279 54815 25285
rect 54757 25245 54769 25279
rect 54803 25245 54815 25279
rect 54757 25239 54815 25245
rect 55953 25279 56011 25285
rect 55953 25245 55965 25279
rect 55999 25276 56011 25279
rect 56226 25276 56232 25288
rect 55999 25248 56232 25276
rect 55999 25245 56011 25248
rect 55953 25239 56011 25245
rect 54404 25208 54432 25239
rect 54665 25211 54723 25217
rect 54665 25208 54677 25211
rect 53944 25180 54340 25208
rect 54404 25180 54677 25208
rect 53009 25143 53067 25149
rect 53009 25140 53021 25143
rect 49200 25112 53021 25140
rect 49200 25100 49206 25112
rect 53009 25109 53021 25112
rect 53055 25109 53067 25143
rect 53009 25103 53067 25109
rect 53466 25100 53472 25152
rect 53524 25100 53530 25152
rect 54312 25149 54340 25180
rect 54665 25177 54677 25180
rect 54711 25177 54723 25211
rect 54772 25208 54800 25239
rect 56226 25236 56232 25248
rect 56284 25236 56290 25288
rect 57146 25236 57152 25288
rect 57204 25236 57210 25288
rect 57241 25279 57299 25285
rect 57241 25245 57253 25279
rect 57287 25245 57299 25279
rect 57340 25276 57368 25316
rect 57425 25313 57437 25347
rect 57471 25344 57483 25347
rect 57701 25347 57759 25353
rect 57701 25344 57713 25347
rect 57471 25316 57713 25344
rect 57471 25313 57483 25316
rect 57425 25307 57483 25313
rect 57701 25313 57713 25316
rect 57747 25313 57759 25347
rect 57974 25344 57980 25356
rect 57701 25307 57759 25313
rect 57808 25316 57980 25344
rect 57808 25285 57836 25316
rect 57974 25304 57980 25316
rect 58032 25304 58038 25356
rect 58066 25304 58072 25356
rect 58124 25344 58130 25356
rect 58124 25316 58204 25344
rect 58124 25304 58130 25316
rect 58176 25285 58204 25316
rect 57609 25279 57667 25285
rect 57609 25276 57621 25279
rect 57340 25248 57621 25276
rect 57241 25239 57299 25245
rect 57609 25245 57621 25248
rect 57655 25276 57667 25279
rect 57793 25279 57851 25285
rect 57655 25248 57744 25276
rect 57655 25245 57667 25248
rect 57609 25239 57667 25245
rect 55030 25208 55036 25220
rect 54772 25180 55036 25208
rect 54665 25171 54723 25177
rect 55030 25168 55036 25180
rect 55088 25168 55094 25220
rect 56594 25168 56600 25220
rect 56652 25208 56658 25220
rect 57256 25208 57284 25239
rect 57716 25208 57744 25248
rect 57793 25245 57805 25279
rect 57839 25245 57851 25279
rect 57793 25239 57851 25245
rect 57885 25279 57943 25285
rect 57885 25245 57897 25279
rect 57931 25245 57943 25279
rect 57885 25239 57943 25245
rect 58161 25279 58219 25285
rect 58161 25245 58173 25279
rect 58207 25245 58219 25279
rect 58161 25239 58219 25245
rect 57900 25208 57928 25239
rect 58618 25208 58624 25220
rect 56652 25180 57652 25208
rect 57716 25180 57836 25208
rect 57900 25180 58624 25208
rect 56652 25168 56658 25180
rect 57624 25152 57652 25180
rect 57808 25152 57836 25180
rect 58618 25168 58624 25180
rect 58676 25168 58682 25220
rect 54297 25143 54355 25149
rect 54297 25109 54309 25143
rect 54343 25109 54355 25143
rect 54297 25103 54355 25109
rect 55306 25100 55312 25152
rect 55364 25100 55370 25152
rect 57422 25100 57428 25152
rect 57480 25100 57486 25152
rect 57606 25100 57612 25152
rect 57664 25100 57670 25152
rect 57790 25100 57796 25152
rect 57848 25100 57854 25152
rect 58066 25100 58072 25152
rect 58124 25100 58130 25152
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 3694 24896 3700 24948
rect 3752 24936 3758 24948
rect 4065 24939 4123 24945
rect 4065 24936 4077 24939
rect 3752 24908 4077 24936
rect 3752 24896 3758 24908
rect 4065 24905 4077 24908
rect 4111 24905 4123 24939
rect 4065 24899 4123 24905
rect 5718 24896 5724 24948
rect 5776 24936 5782 24948
rect 5905 24939 5963 24945
rect 5905 24936 5917 24939
rect 5776 24908 5917 24936
rect 5776 24896 5782 24908
rect 5905 24905 5917 24908
rect 5951 24905 5963 24939
rect 5905 24899 5963 24905
rect 11977 24939 12035 24945
rect 11977 24905 11989 24939
rect 12023 24936 12035 24939
rect 12526 24936 12532 24948
rect 12023 24908 12532 24936
rect 12023 24905 12035 24908
rect 11977 24899 12035 24905
rect 12526 24896 12532 24908
rect 12584 24896 12590 24948
rect 12618 24896 12624 24948
rect 12676 24896 12682 24948
rect 13078 24896 13084 24948
rect 13136 24936 13142 24948
rect 14553 24939 14611 24945
rect 14553 24936 14565 24939
rect 13136 24908 14565 24936
rect 13136 24896 13142 24908
rect 14553 24905 14565 24908
rect 14599 24905 14611 24939
rect 14553 24899 14611 24905
rect 38381 24939 38439 24945
rect 38381 24905 38393 24939
rect 38427 24936 38439 24939
rect 38930 24936 38936 24948
rect 38427 24908 38936 24936
rect 38427 24905 38439 24908
rect 38381 24899 38439 24905
rect 38930 24896 38936 24908
rect 38988 24896 38994 24948
rect 40034 24896 40040 24948
rect 40092 24896 40098 24948
rect 40497 24939 40555 24945
rect 40497 24905 40509 24939
rect 40543 24936 40555 24939
rect 41046 24936 41052 24948
rect 40543 24908 41052 24936
rect 40543 24905 40555 24908
rect 40497 24899 40555 24905
rect 41046 24896 41052 24908
rect 41104 24896 41110 24948
rect 41601 24939 41659 24945
rect 41601 24905 41613 24939
rect 41647 24936 41659 24939
rect 41874 24936 41880 24948
rect 41647 24908 41880 24936
rect 41647 24905 41659 24908
rect 41601 24899 41659 24905
rect 41874 24896 41880 24908
rect 41932 24896 41938 24948
rect 42702 24896 42708 24948
rect 42760 24896 42766 24948
rect 42794 24896 42800 24948
rect 42852 24896 42858 24948
rect 45002 24896 45008 24948
rect 45060 24896 45066 24948
rect 45738 24896 45744 24948
rect 45796 24896 45802 24948
rect 46753 24939 46811 24945
rect 46753 24936 46765 24939
rect 46032 24908 46765 24936
rect 5442 24828 5448 24880
rect 5500 24868 5506 24880
rect 10042 24868 10048 24880
rect 5500 24840 10048 24868
rect 5500 24828 5506 24840
rect 10042 24828 10048 24840
rect 10100 24868 10106 24880
rect 13446 24877 13452 24880
rect 12161 24871 12219 24877
rect 12161 24868 12173 24871
rect 10100 24840 12173 24868
rect 10100 24828 10106 24840
rect 12161 24837 12173 24840
rect 12207 24837 12219 24871
rect 13440 24868 13452 24877
rect 13407 24840 13452 24868
rect 12161 24831 12219 24837
rect 13440 24831 13452 24840
rect 13446 24828 13452 24831
rect 13504 24828 13510 24880
rect 38120 24840 38884 24868
rect 2682 24760 2688 24812
rect 2740 24760 2746 24812
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24800 12311 24803
rect 12529 24803 12587 24809
rect 12299 24772 12434 24800
rect 12299 24769 12311 24772
rect 12253 24763 12311 24769
rect 934 24692 940 24744
rect 992 24732 998 24744
rect 1581 24735 1639 24741
rect 1581 24732 1593 24735
rect 992 24704 1593 24732
rect 992 24692 998 24704
rect 1581 24701 1593 24704
rect 1627 24701 1639 24735
rect 1581 24695 1639 24701
rect 3694 24692 3700 24744
rect 3752 24692 3758 24744
rect 7282 24692 7288 24744
rect 7340 24732 7346 24744
rect 11330 24732 11336 24744
rect 7340 24704 11336 24732
rect 7340 24692 7346 24704
rect 11330 24692 11336 24704
rect 11388 24692 11394 24744
rect 7834 24624 7840 24676
rect 7892 24664 7898 24676
rect 7892 24636 10640 24664
rect 7892 24624 7898 24636
rect 10612 24608 10640 24636
rect 11882 24624 11888 24676
rect 11940 24664 11946 24676
rect 12406 24664 12434 24772
rect 12529 24769 12541 24803
rect 12575 24769 12587 24803
rect 12529 24763 12587 24769
rect 12544 24732 12572 24763
rect 12986 24760 12992 24812
rect 13044 24800 13050 24812
rect 13173 24803 13231 24809
rect 13173 24800 13185 24803
rect 13044 24772 13185 24800
rect 13044 24760 13050 24772
rect 13173 24769 13185 24772
rect 13219 24769 13231 24803
rect 13173 24763 13231 24769
rect 36814 24760 36820 24812
rect 36872 24760 36878 24812
rect 37366 24760 37372 24812
rect 37424 24800 37430 24812
rect 37461 24803 37519 24809
rect 37461 24800 37473 24803
rect 37424 24772 37473 24800
rect 37424 24760 37430 24772
rect 37461 24769 37473 24772
rect 37507 24769 37519 24803
rect 37461 24763 37519 24769
rect 37645 24803 37703 24809
rect 37645 24769 37657 24803
rect 37691 24800 37703 24803
rect 38120 24800 38148 24840
rect 37691 24772 38148 24800
rect 38197 24803 38255 24809
rect 37691 24769 37703 24772
rect 37645 24763 37703 24769
rect 38197 24769 38209 24803
rect 38243 24769 38255 24803
rect 38197 24763 38255 24769
rect 12710 24732 12716 24744
rect 12544 24704 12716 24732
rect 12710 24692 12716 24704
rect 12768 24692 12774 24744
rect 36832 24732 36860 24760
rect 37182 24732 37188 24744
rect 36832 24704 37188 24732
rect 37182 24692 37188 24704
rect 37240 24732 37246 24744
rect 37737 24735 37795 24741
rect 37737 24732 37749 24735
rect 37240 24704 37749 24732
rect 37240 24692 37246 24704
rect 37737 24701 37749 24704
rect 37783 24701 37795 24735
rect 38212 24732 38240 24763
rect 38470 24760 38476 24812
rect 38528 24760 38534 24812
rect 38749 24803 38807 24809
rect 38749 24769 38761 24803
rect 38795 24769 38807 24803
rect 38856 24800 38884 24840
rect 39022 24800 39028 24812
rect 38856 24772 39028 24800
rect 38749 24763 38807 24769
rect 38764 24732 38792 24763
rect 39022 24760 39028 24772
rect 39080 24760 39086 24812
rect 39758 24760 39764 24812
rect 39816 24760 39822 24812
rect 39945 24803 40003 24809
rect 39945 24769 39957 24803
rect 39991 24800 40003 24803
rect 40052 24800 40080 24896
rect 41340 24840 41644 24868
rect 39991 24772 40080 24800
rect 40405 24803 40463 24809
rect 39991 24769 40003 24772
rect 39945 24763 40003 24769
rect 40405 24769 40417 24803
rect 40451 24769 40463 24803
rect 40405 24763 40463 24769
rect 38212 24704 38792 24732
rect 37737 24695 37795 24701
rect 12526 24664 12532 24676
rect 11940 24636 12296 24664
rect 12406 24636 12532 24664
rect 11940 24624 11946 24636
rect 3050 24556 3056 24608
rect 3108 24596 3114 24608
rect 3145 24599 3203 24605
rect 3145 24596 3157 24599
rect 3108 24568 3157 24596
rect 3108 24556 3114 24568
rect 3145 24565 3157 24568
rect 3191 24565 3203 24599
rect 3145 24559 3203 24565
rect 9674 24556 9680 24608
rect 9732 24596 9738 24608
rect 10137 24599 10195 24605
rect 10137 24596 10149 24599
rect 9732 24568 10149 24596
rect 9732 24556 9738 24568
rect 10137 24565 10149 24568
rect 10183 24565 10195 24599
rect 10137 24559 10195 24565
rect 10594 24556 10600 24608
rect 10652 24556 10658 24608
rect 12268 24596 12296 24636
rect 12526 24624 12532 24636
rect 12584 24664 12590 24676
rect 12989 24667 13047 24673
rect 12989 24664 13001 24667
rect 12584 24636 13001 24664
rect 12584 24624 12590 24636
rect 12989 24633 13001 24636
rect 13035 24633 13047 24667
rect 12989 24627 13047 24633
rect 37366 24624 37372 24676
rect 37424 24664 37430 24676
rect 38657 24667 38715 24673
rect 38657 24664 38669 24667
rect 37424 24636 38669 24664
rect 37424 24624 37430 24636
rect 38657 24633 38669 24636
rect 38703 24633 38715 24667
rect 38764 24664 38792 24704
rect 39853 24735 39911 24741
rect 39853 24701 39865 24735
rect 39899 24732 39911 24735
rect 40420 24732 40448 24763
rect 40678 24760 40684 24812
rect 40736 24760 40742 24812
rect 40865 24803 40923 24809
rect 40865 24769 40877 24803
rect 40911 24800 40923 24803
rect 40954 24800 40960 24812
rect 40911 24772 40960 24800
rect 40911 24769 40923 24772
rect 40865 24763 40923 24769
rect 40954 24760 40960 24772
rect 41012 24800 41018 24812
rect 41340 24809 41368 24840
rect 41616 24812 41644 24840
rect 42886 24828 42892 24880
rect 42944 24868 42950 24880
rect 45020 24868 45048 24896
rect 42944 24840 44036 24868
rect 42944 24828 42950 24840
rect 41233 24803 41291 24809
rect 41233 24800 41245 24803
rect 41012 24772 41245 24800
rect 41012 24760 41018 24772
rect 41233 24769 41245 24772
rect 41279 24769 41291 24803
rect 41233 24763 41291 24769
rect 41325 24803 41383 24809
rect 41325 24769 41337 24803
rect 41371 24769 41383 24803
rect 41325 24763 41383 24769
rect 41506 24760 41512 24812
rect 41564 24760 41570 24812
rect 41598 24760 41604 24812
rect 41656 24760 41662 24812
rect 41693 24803 41751 24809
rect 41693 24769 41705 24803
rect 41739 24769 41751 24803
rect 41693 24763 41751 24769
rect 43717 24803 43775 24809
rect 43717 24769 43729 24803
rect 43763 24769 43775 24803
rect 43717 24763 43775 24769
rect 39899 24704 40448 24732
rect 39899 24701 39911 24704
rect 39853 24695 39911 24701
rect 40865 24667 40923 24673
rect 40865 24664 40877 24667
rect 38764 24636 40877 24664
rect 38657 24627 38715 24633
rect 40865 24633 40877 24636
rect 40911 24633 40923 24667
rect 41708 24664 41736 24763
rect 43441 24735 43499 24741
rect 43441 24701 43453 24735
rect 43487 24732 43499 24735
rect 43533 24735 43591 24741
rect 43533 24732 43545 24735
rect 43487 24704 43545 24732
rect 43487 24701 43499 24704
rect 43441 24695 43499 24701
rect 43533 24701 43545 24704
rect 43579 24701 43591 24735
rect 43732 24732 43760 24763
rect 43806 24760 43812 24812
rect 43864 24760 43870 24812
rect 44008 24809 44036 24840
rect 44100 24840 45048 24868
rect 45756 24868 45784 24896
rect 45925 24871 45983 24877
rect 45925 24868 45937 24871
rect 45756 24840 45937 24868
rect 44100 24809 44128 24840
rect 45925 24837 45937 24840
rect 45971 24837 45983 24871
rect 45925 24831 45983 24837
rect 43993 24803 44051 24809
rect 43993 24769 44005 24803
rect 44039 24769 44051 24803
rect 43993 24763 44051 24769
rect 44085 24803 44143 24809
rect 44085 24769 44097 24803
rect 44131 24769 44143 24803
rect 44085 24763 44143 24769
rect 44174 24760 44180 24812
rect 44232 24800 44238 24812
rect 44358 24800 44364 24812
rect 44232 24772 44364 24800
rect 44232 24760 44238 24772
rect 44358 24760 44364 24772
rect 44416 24760 44422 24812
rect 44450 24760 44456 24812
rect 44508 24760 44514 24812
rect 44542 24760 44548 24812
rect 44600 24760 44606 24812
rect 44637 24803 44695 24809
rect 44637 24769 44649 24803
rect 44683 24769 44695 24803
rect 44637 24763 44695 24769
rect 44652 24732 44680 24763
rect 45186 24760 45192 24812
rect 45244 24800 45250 24812
rect 45281 24803 45339 24809
rect 45281 24800 45293 24803
rect 45244 24772 45293 24800
rect 45244 24760 45250 24772
rect 45281 24769 45293 24772
rect 45327 24769 45339 24803
rect 45281 24763 45339 24769
rect 45370 24760 45376 24812
rect 45428 24800 45434 24812
rect 45465 24803 45523 24809
rect 45465 24800 45477 24803
rect 45428 24772 45477 24800
rect 45428 24760 45434 24772
rect 45465 24769 45477 24772
rect 45511 24800 45523 24803
rect 46032 24800 46060 24908
rect 46753 24905 46765 24908
rect 46799 24905 46811 24939
rect 48593 24939 48651 24945
rect 46753 24899 46811 24905
rect 46860 24908 48084 24936
rect 46198 24828 46204 24880
rect 46256 24868 46262 24880
rect 46860 24868 46888 24908
rect 46256 24840 46888 24868
rect 46921 24871 46979 24877
rect 46256 24828 46262 24840
rect 46921 24837 46933 24871
rect 46967 24868 46979 24871
rect 46967 24837 46980 24868
rect 46921 24831 46980 24837
rect 45511 24772 46060 24800
rect 46109 24803 46167 24809
rect 45511 24769 45523 24772
rect 45465 24763 45523 24769
rect 46109 24769 46121 24803
rect 46155 24800 46167 24803
rect 46216 24800 46244 24828
rect 46155 24772 46244 24800
rect 46155 24769 46167 24772
rect 46109 24763 46167 24769
rect 46382 24760 46388 24812
rect 46440 24760 46446 24812
rect 46477 24803 46535 24809
rect 46477 24769 46489 24803
rect 46523 24769 46535 24803
rect 46477 24763 46535 24769
rect 45002 24732 45008 24744
rect 43732 24704 44036 24732
rect 44652 24704 45008 24732
rect 43533 24695 43591 24701
rect 44008 24676 44036 24704
rect 45002 24692 45008 24704
rect 45060 24732 45066 24744
rect 46492 24732 46520 24763
rect 46658 24760 46664 24812
rect 46716 24760 46722 24812
rect 45060 24704 46520 24732
rect 46952 24732 46980 24831
rect 47026 24828 47032 24880
rect 47084 24868 47090 24880
rect 47121 24871 47179 24877
rect 47121 24868 47133 24871
rect 47084 24840 47133 24868
rect 47084 24828 47090 24840
rect 47121 24837 47133 24840
rect 47167 24868 47179 24871
rect 47305 24871 47363 24877
rect 47305 24868 47317 24871
rect 47167 24840 47317 24868
rect 47167 24837 47179 24840
rect 47121 24831 47179 24837
rect 47305 24837 47317 24840
rect 47351 24837 47363 24871
rect 47305 24831 47363 24837
rect 47670 24828 47676 24880
rect 47728 24868 47734 24880
rect 47728 24840 47992 24868
rect 47728 24828 47734 24840
rect 47210 24760 47216 24812
rect 47268 24760 47274 24812
rect 47394 24760 47400 24812
rect 47452 24800 47458 24812
rect 47964 24809 47992 24840
rect 48056 24809 48084 24908
rect 48593 24905 48605 24939
rect 48639 24936 48651 24939
rect 48774 24936 48780 24948
rect 48639 24908 48780 24936
rect 48639 24905 48651 24908
rect 48593 24899 48651 24905
rect 48774 24896 48780 24908
rect 48832 24896 48838 24948
rect 53098 24936 53104 24948
rect 51644 24908 53104 24936
rect 48406 24828 48412 24880
rect 48464 24868 48470 24880
rect 49234 24868 49240 24880
rect 48464 24840 49240 24868
rect 48464 24828 48470 24840
rect 49234 24828 49240 24840
rect 49292 24868 49298 24880
rect 51644 24868 51672 24908
rect 53098 24896 53104 24908
rect 53156 24896 53162 24948
rect 53466 24896 53472 24948
rect 53524 24896 53530 24948
rect 53742 24896 53748 24948
rect 53800 24896 53806 24948
rect 57422 24896 57428 24948
rect 57480 24896 57486 24948
rect 58066 24896 58072 24948
rect 58124 24896 58130 24948
rect 52454 24868 52460 24880
rect 49292 24840 49450 24868
rect 51552 24840 51672 24868
rect 51736 24840 52460 24868
rect 49292 24828 49298 24840
rect 47949 24803 48007 24809
rect 47452 24772 47900 24800
rect 47452 24760 47458 24772
rect 47486 24732 47492 24744
rect 46952 24704 47492 24732
rect 45060 24692 45066 24704
rect 41708 24636 43944 24664
rect 40865 24627 40923 24633
rect 13170 24596 13176 24608
rect 12268 24568 13176 24596
rect 13170 24556 13176 24568
rect 13228 24596 13234 24608
rect 35894 24596 35900 24608
rect 13228 24568 35900 24596
rect 13228 24556 13234 24568
rect 35894 24556 35900 24568
rect 35952 24596 35958 24608
rect 36722 24596 36728 24608
rect 35952 24568 36728 24596
rect 35952 24556 35958 24568
rect 36722 24556 36728 24568
rect 36780 24596 36786 24608
rect 37001 24599 37059 24605
rect 37001 24596 37013 24599
rect 36780 24568 37013 24596
rect 36780 24556 36786 24568
rect 37001 24565 37013 24568
rect 37047 24565 37059 24599
rect 37001 24559 37059 24565
rect 37274 24556 37280 24608
rect 37332 24556 37338 24608
rect 38010 24556 38016 24608
rect 38068 24556 38074 24608
rect 42061 24599 42119 24605
rect 42061 24565 42073 24599
rect 42107 24596 42119 24599
rect 42242 24596 42248 24608
rect 42107 24568 42248 24596
rect 42107 24565 42119 24568
rect 42061 24559 42119 24565
rect 42242 24556 42248 24568
rect 42300 24556 42306 24608
rect 43916 24596 43944 24636
rect 43990 24624 43996 24676
rect 44048 24624 44054 24676
rect 44315 24667 44373 24673
rect 44315 24633 44327 24667
rect 44361 24664 44373 24667
rect 45646 24664 45652 24676
rect 44361 24636 45652 24664
rect 44361 24633 44373 24636
rect 44315 24627 44373 24633
rect 45646 24624 45652 24636
rect 45704 24624 45710 24676
rect 45830 24624 45836 24676
rect 45888 24664 45894 24676
rect 46952 24664 46980 24704
rect 47486 24692 47492 24704
rect 47544 24692 47550 24744
rect 47872 24673 47900 24772
rect 47949 24769 47961 24803
rect 47995 24769 48007 24803
rect 47949 24763 48007 24769
rect 48041 24803 48099 24809
rect 48041 24769 48053 24803
rect 48087 24769 48099 24803
rect 48041 24763 48099 24769
rect 48222 24760 48228 24812
rect 48280 24760 48286 24812
rect 48317 24803 48375 24809
rect 48317 24769 48329 24803
rect 48363 24769 48375 24803
rect 48317 24763 48375 24769
rect 48133 24735 48191 24741
rect 48133 24701 48145 24735
rect 48179 24732 48191 24735
rect 48332 24732 48360 24763
rect 48498 24760 48504 24812
rect 48556 24800 48562 24812
rect 48685 24803 48743 24809
rect 48685 24800 48697 24803
rect 48556 24772 48697 24800
rect 48556 24760 48562 24772
rect 48685 24769 48697 24772
rect 48731 24769 48743 24803
rect 48685 24763 48743 24769
rect 50893 24803 50951 24809
rect 50893 24769 50905 24803
rect 50939 24769 50951 24803
rect 50893 24763 50951 24769
rect 51353 24803 51411 24809
rect 51353 24769 51365 24803
rect 51399 24800 51411 24803
rect 51552 24800 51580 24840
rect 51399 24772 51580 24800
rect 51399 24769 51411 24772
rect 51353 24763 51411 24769
rect 48179 24704 48360 24732
rect 48179 24701 48191 24704
rect 48133 24695 48191 24701
rect 48590 24692 48596 24744
rect 48648 24692 48654 24744
rect 48958 24692 48964 24744
rect 49016 24692 49022 24744
rect 45888 24636 46980 24664
rect 47857 24667 47915 24673
rect 45888 24624 45894 24636
rect 47857 24633 47869 24667
rect 47903 24664 47915 24667
rect 50908 24664 50936 24763
rect 51626 24760 51632 24812
rect 51684 24800 51690 24812
rect 51736 24800 51764 24840
rect 52454 24828 52460 24840
rect 52512 24868 52518 24880
rect 53484 24868 53512 24896
rect 52512 24840 52776 24868
rect 52512 24828 52518 24840
rect 51684 24772 51764 24800
rect 51684 24760 51690 24772
rect 51810 24760 51816 24812
rect 51868 24760 51874 24812
rect 51905 24803 51963 24809
rect 51905 24769 51917 24803
rect 51951 24769 51963 24803
rect 51905 24763 51963 24769
rect 51920 24732 51948 24763
rect 52086 24760 52092 24812
rect 52144 24760 52150 24812
rect 52748 24809 52776 24840
rect 52932 24840 53512 24868
rect 54941 24871 54999 24877
rect 52932 24809 52960 24840
rect 54941 24837 54953 24871
rect 54987 24868 54999 24871
rect 54987 24840 55260 24868
rect 54987 24837 54999 24840
rect 54941 24831 54999 24837
rect 52733 24803 52791 24809
rect 52733 24769 52745 24803
rect 52779 24769 52791 24803
rect 52733 24763 52791 24769
rect 52917 24803 52975 24809
rect 52917 24769 52929 24803
rect 52963 24769 52975 24803
rect 52917 24763 52975 24769
rect 53009 24803 53067 24809
rect 53009 24769 53021 24803
rect 53055 24769 53067 24803
rect 53009 24763 53067 24769
rect 53193 24803 53251 24809
rect 53193 24769 53205 24803
rect 53239 24769 53251 24803
rect 53193 24763 53251 24769
rect 53285 24803 53343 24809
rect 53285 24769 53297 24803
rect 53331 24800 53343 24803
rect 53374 24800 53380 24812
rect 53331 24772 53380 24800
rect 53331 24769 53343 24772
rect 53285 24763 53343 24769
rect 47903 24636 48636 24664
rect 47903 24633 47915 24636
rect 47857 24627 47915 24633
rect 45370 24596 45376 24608
rect 43916 24568 45376 24596
rect 45370 24556 45376 24568
rect 45428 24556 45434 24608
rect 45462 24556 45468 24608
rect 45520 24556 45526 24608
rect 46198 24556 46204 24608
rect 46256 24596 46262 24608
rect 46937 24599 46995 24605
rect 46937 24596 46949 24599
rect 46256 24568 46949 24596
rect 46256 24556 46262 24568
rect 46937 24565 46949 24568
rect 46983 24565 46995 24599
rect 46937 24559 46995 24565
rect 47118 24556 47124 24608
rect 47176 24596 47182 24608
rect 48406 24596 48412 24608
rect 47176 24568 48412 24596
rect 47176 24556 47182 24568
rect 48406 24556 48412 24568
rect 48464 24556 48470 24608
rect 48608 24596 48636 24636
rect 49988 24636 50936 24664
rect 51092 24704 51948 24732
rect 52825 24735 52883 24741
rect 49988 24596 50016 24636
rect 51092 24608 51120 24704
rect 52825 24701 52837 24735
rect 52871 24732 52883 24735
rect 53024 24732 53052 24763
rect 52871 24704 53052 24732
rect 53208 24732 53236 24763
rect 53374 24760 53380 24772
rect 53432 24760 53438 24812
rect 53469 24803 53527 24809
rect 53469 24769 53481 24803
rect 53515 24800 53527 24803
rect 53558 24800 53564 24812
rect 53515 24772 53564 24800
rect 53515 24769 53527 24772
rect 53469 24763 53527 24769
rect 53558 24760 53564 24772
rect 53616 24760 53622 24812
rect 54665 24803 54723 24809
rect 54665 24769 54677 24803
rect 54711 24800 54723 24803
rect 55033 24803 55091 24809
rect 54711 24772 54892 24800
rect 54711 24769 54723 24772
rect 54665 24763 54723 24769
rect 53208 24704 53328 24732
rect 52871 24701 52883 24704
rect 52825 24695 52883 24701
rect 51997 24667 52055 24673
rect 51997 24664 52009 24667
rect 51460 24636 52009 24664
rect 51460 24608 51488 24636
rect 51997 24633 52009 24636
rect 52043 24633 52055 24667
rect 51997 24627 52055 24633
rect 48608 24568 50016 24596
rect 50433 24599 50491 24605
rect 50433 24565 50445 24599
rect 50479 24596 50491 24599
rect 51074 24596 51080 24608
rect 50479 24568 51080 24596
rect 50479 24565 50491 24568
rect 50433 24559 50491 24565
rect 51074 24556 51080 24568
rect 51132 24556 51138 24608
rect 51442 24556 51448 24608
rect 51500 24556 51506 24608
rect 51718 24556 51724 24608
rect 51776 24556 51782 24608
rect 52362 24556 52368 24608
rect 52420 24596 52426 24608
rect 53101 24599 53159 24605
rect 53101 24596 53113 24599
rect 52420 24568 53113 24596
rect 52420 24556 52426 24568
rect 53101 24565 53113 24568
rect 53147 24565 53159 24599
rect 53300 24596 53328 24704
rect 54754 24692 54760 24744
rect 54812 24692 54818 24744
rect 54864 24608 54892 24772
rect 55033 24769 55045 24803
rect 55079 24800 55091 24803
rect 55122 24800 55128 24812
rect 55079 24772 55128 24800
rect 55079 24769 55091 24772
rect 55033 24763 55091 24769
rect 55122 24760 55128 24772
rect 55180 24760 55186 24812
rect 55232 24800 55260 24840
rect 55289 24803 55347 24809
rect 55289 24800 55301 24803
rect 55232 24772 55301 24800
rect 55289 24769 55301 24772
rect 55335 24769 55347 24803
rect 56965 24803 57023 24809
rect 56965 24800 56977 24803
rect 55289 24763 55347 24769
rect 56796 24772 56977 24800
rect 54941 24735 54999 24741
rect 54941 24701 54953 24735
rect 54987 24701 54999 24735
rect 54941 24695 54999 24701
rect 53377 24599 53435 24605
rect 53377 24596 53389 24599
rect 53300 24568 53389 24596
rect 53101 24559 53159 24565
rect 53377 24565 53389 24568
rect 53423 24565 53435 24599
rect 53377 24559 53435 24565
rect 54846 24556 54852 24608
rect 54904 24556 54910 24608
rect 54956 24596 54984 24695
rect 56042 24624 56048 24676
rect 56100 24664 56106 24676
rect 56796 24673 56824 24772
rect 56965 24769 56977 24772
rect 57011 24769 57023 24803
rect 56965 24763 57023 24769
rect 57149 24803 57207 24809
rect 57149 24769 57161 24803
rect 57195 24800 57207 24803
rect 57440 24800 57468 24896
rect 58084 24868 58112 24896
rect 58084 24840 58204 24868
rect 58176 24809 58204 24840
rect 57195 24772 57468 24800
rect 58069 24803 58127 24809
rect 57195 24769 57207 24772
rect 57149 24763 57207 24769
rect 58069 24769 58081 24803
rect 58115 24769 58127 24803
rect 58069 24763 58127 24769
rect 58161 24803 58219 24809
rect 58161 24769 58173 24803
rect 58207 24769 58219 24803
rect 58161 24763 58219 24769
rect 57974 24692 57980 24744
rect 58032 24692 58038 24744
rect 58084 24732 58112 24763
rect 58084 24704 58756 24732
rect 56781 24667 56839 24673
rect 56781 24664 56793 24667
rect 56100 24636 56793 24664
rect 56100 24624 56106 24636
rect 56781 24633 56793 24636
rect 56827 24633 56839 24667
rect 57992 24664 58020 24692
rect 58253 24667 58311 24673
rect 58253 24664 58265 24667
rect 57992 24636 58265 24664
rect 56781 24627 56839 24633
rect 58253 24633 58265 24636
rect 58299 24633 58311 24667
rect 58253 24627 58311 24633
rect 58728 24608 58756 24704
rect 55306 24596 55312 24608
rect 54956 24568 55312 24596
rect 55306 24556 55312 24568
rect 55364 24556 55370 24608
rect 55950 24556 55956 24608
rect 56008 24596 56014 24608
rect 56413 24599 56471 24605
rect 56413 24596 56425 24599
rect 56008 24568 56425 24596
rect 56008 24556 56014 24568
rect 56413 24565 56425 24568
rect 56459 24565 56471 24599
rect 56413 24559 56471 24565
rect 57054 24556 57060 24608
rect 57112 24556 57118 24608
rect 57882 24556 57888 24608
rect 57940 24556 57946 24608
rect 58710 24556 58716 24608
rect 58768 24556 58774 24608
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 3050 24352 3056 24404
rect 3108 24352 3114 24404
rect 3326 24352 3332 24404
rect 3384 24352 3390 24404
rect 3421 24395 3479 24401
rect 3421 24361 3433 24395
rect 3467 24392 3479 24395
rect 3694 24392 3700 24404
rect 3467 24364 3700 24392
rect 3467 24361 3479 24364
rect 3421 24355 3479 24361
rect 3694 24352 3700 24364
rect 3752 24352 3758 24404
rect 6730 24352 6736 24404
rect 6788 24352 6794 24404
rect 7929 24395 7987 24401
rect 7929 24392 7941 24395
rect 6932 24364 7941 24392
rect 2869 24259 2927 24265
rect 2869 24225 2881 24259
rect 2915 24256 2927 24259
rect 3068 24256 3096 24352
rect 4890 24284 4896 24336
rect 4948 24284 4954 24336
rect 2915 24228 3096 24256
rect 2915 24225 2927 24228
rect 2869 24219 2927 24225
rect 3142 24216 3148 24268
rect 3200 24216 3206 24268
rect 6748 24265 6776 24352
rect 3513 24259 3571 24265
rect 3513 24225 3525 24259
rect 3559 24256 3571 24259
rect 3789 24259 3847 24265
rect 3789 24256 3801 24259
rect 3559 24228 3801 24256
rect 3559 24225 3571 24228
rect 3513 24219 3571 24225
rect 3789 24225 3801 24228
rect 3835 24225 3847 24259
rect 3789 24219 3847 24225
rect 6733 24259 6791 24265
rect 6733 24225 6745 24259
rect 6779 24225 6791 24259
rect 6733 24219 6791 24225
rect 3234 24148 3240 24200
rect 3292 24148 3298 24200
rect 4338 24148 4344 24200
rect 4396 24148 4402 24200
rect 4617 24191 4675 24197
rect 4617 24157 4629 24191
rect 4663 24157 4675 24191
rect 4617 24151 4675 24157
rect 2406 24080 2412 24132
rect 2464 24080 2470 24132
rect 2866 24080 2872 24132
rect 2924 24120 2930 24132
rect 3326 24120 3332 24132
rect 2924 24092 3332 24120
rect 2924 24080 2930 24092
rect 3326 24080 3332 24092
rect 3384 24080 3390 24132
rect 4632 24064 4660 24151
rect 4706 24148 4712 24200
rect 4764 24148 4770 24200
rect 5718 24148 5724 24200
rect 5776 24188 5782 24200
rect 6546 24188 6552 24200
rect 5776 24160 6552 24188
rect 5776 24148 5782 24160
rect 6546 24148 6552 24160
rect 6604 24188 6610 24200
rect 6932 24197 6960 24364
rect 7929 24361 7941 24364
rect 7975 24392 7987 24395
rect 9674 24392 9680 24404
rect 7975 24364 9680 24392
rect 7975 24361 7987 24364
rect 7929 24355 7987 24361
rect 9674 24352 9680 24364
rect 9732 24352 9738 24404
rect 9950 24352 9956 24404
rect 10008 24352 10014 24404
rect 11885 24395 11943 24401
rect 11885 24392 11897 24395
rect 10152 24364 11897 24392
rect 7650 24284 7656 24336
rect 7708 24284 7714 24336
rect 8478 24284 8484 24336
rect 8536 24284 8542 24336
rect 7484 24228 8340 24256
rect 6917 24191 6975 24197
rect 6917 24188 6929 24191
rect 6604 24160 6929 24188
rect 6604 24148 6610 24160
rect 6917 24157 6929 24160
rect 6963 24157 6975 24191
rect 6917 24151 6975 24157
rect 7006 24148 7012 24200
rect 7064 24148 7070 24200
rect 7374 24148 7380 24200
rect 7432 24148 7438 24200
rect 7484 24197 7512 24228
rect 8312 24200 8340 24228
rect 7469 24191 7527 24197
rect 7469 24157 7481 24191
rect 7515 24157 7527 24191
rect 7469 24151 7527 24157
rect 7576 24160 8156 24188
rect 7576 24132 7604 24160
rect 4893 24123 4951 24129
rect 4893 24089 4905 24123
rect 4939 24120 4951 24123
rect 5258 24120 5264 24132
rect 4939 24092 5264 24120
rect 4939 24089 4951 24092
rect 4893 24083 4951 24089
rect 5258 24080 5264 24092
rect 5316 24120 5322 24132
rect 5316 24092 7512 24120
rect 5316 24080 5322 24092
rect 1397 24055 1455 24061
rect 1397 24021 1409 24055
rect 1443 24052 1455 24055
rect 2682 24052 2688 24064
rect 1443 24024 2688 24052
rect 1443 24021 1455 24024
rect 1397 24015 1455 24021
rect 2682 24012 2688 24024
rect 2740 24012 2746 24064
rect 4614 24012 4620 24064
rect 4672 24012 4678 24064
rect 6362 24012 6368 24064
rect 6420 24052 6426 24064
rect 6733 24055 6791 24061
rect 6733 24052 6745 24055
rect 6420 24024 6745 24052
rect 6420 24012 6426 24024
rect 6733 24021 6745 24024
rect 6779 24021 6791 24055
rect 7484 24052 7512 24092
rect 7558 24080 7564 24132
rect 7616 24080 7622 24132
rect 7653 24123 7711 24129
rect 7653 24089 7665 24123
rect 7699 24120 7711 24123
rect 7834 24120 7840 24132
rect 7699 24092 7840 24120
rect 7699 24089 7711 24092
rect 7653 24083 7711 24089
rect 7668 24052 7696 24083
rect 7834 24080 7840 24092
rect 7892 24080 7898 24132
rect 8128 24120 8156 24160
rect 8202 24148 8208 24200
rect 8260 24148 8266 24200
rect 8294 24148 8300 24200
rect 8352 24148 8358 24200
rect 9692 24188 9720 24352
rect 9769 24259 9827 24265
rect 9769 24225 9781 24259
rect 9815 24256 9827 24259
rect 9968 24256 9996 24352
rect 10152 24256 10180 24364
rect 11885 24361 11897 24364
rect 11931 24361 11943 24395
rect 12434 24392 12440 24404
rect 11885 24355 11943 24361
rect 11992 24364 12440 24392
rect 10413 24327 10471 24333
rect 10413 24293 10425 24327
rect 10459 24293 10471 24327
rect 10413 24287 10471 24293
rect 9815 24228 9996 24256
rect 10060 24228 10180 24256
rect 10428 24256 10456 24287
rect 10428 24228 10640 24256
rect 9815 24225 9827 24228
rect 9769 24219 9827 24225
rect 10060 24200 10088 24228
rect 9953 24191 10011 24197
rect 9953 24188 9965 24191
rect 9692 24160 9965 24188
rect 9953 24157 9965 24160
rect 9999 24157 10011 24191
rect 9953 24151 10011 24157
rect 10042 24148 10048 24200
rect 10100 24148 10106 24200
rect 10134 24148 10140 24200
rect 10192 24148 10198 24200
rect 10502 24148 10508 24200
rect 10560 24148 10566 24200
rect 10612 24188 10640 24228
rect 10761 24191 10819 24197
rect 10761 24188 10773 24191
rect 10612 24160 10773 24188
rect 10761 24157 10773 24160
rect 10807 24157 10819 24191
rect 10761 24151 10819 24157
rect 8481 24123 8539 24129
rect 8481 24120 8493 24123
rect 8128 24092 8493 24120
rect 8481 24089 8493 24092
rect 8527 24120 8539 24123
rect 10413 24123 10471 24129
rect 10413 24120 10425 24123
rect 8527 24092 10425 24120
rect 8527 24089 8539 24092
rect 8481 24083 8539 24089
rect 10413 24089 10425 24092
rect 10459 24120 10471 24123
rect 11992 24120 12020 24364
rect 12434 24352 12440 24364
rect 12492 24392 12498 24404
rect 12894 24392 12900 24404
rect 12492 24364 12900 24392
rect 12492 24352 12498 24364
rect 12894 24352 12900 24364
rect 12952 24352 12958 24404
rect 13630 24352 13636 24404
rect 13688 24392 13694 24404
rect 14277 24395 14335 24401
rect 14277 24392 14289 24395
rect 13688 24364 14289 24392
rect 13688 24352 13694 24364
rect 14277 24361 14289 24364
rect 14323 24361 14335 24395
rect 14277 24355 14335 24361
rect 37182 24352 37188 24404
rect 37240 24392 37246 24404
rect 37737 24395 37795 24401
rect 37737 24392 37749 24395
rect 37240 24364 37749 24392
rect 37240 24352 37246 24364
rect 37737 24361 37749 24364
rect 37783 24361 37795 24395
rect 37737 24355 37795 24361
rect 39022 24352 39028 24404
rect 39080 24392 39086 24404
rect 39577 24395 39635 24401
rect 39577 24392 39589 24395
rect 39080 24364 39589 24392
rect 39080 24352 39086 24364
rect 39577 24361 39589 24364
rect 39623 24361 39635 24395
rect 39577 24355 39635 24361
rect 40034 24352 40040 24404
rect 40092 24352 40098 24404
rect 43806 24352 43812 24404
rect 43864 24392 43870 24404
rect 44545 24395 44603 24401
rect 44545 24392 44557 24395
rect 43864 24364 44557 24392
rect 43864 24352 43870 24364
rect 44545 24361 44557 24364
rect 44591 24361 44603 24395
rect 44545 24355 44603 24361
rect 45002 24352 45008 24404
rect 45060 24352 45066 24404
rect 45462 24352 45468 24404
rect 45520 24352 45526 24404
rect 47118 24352 47124 24404
rect 47176 24392 47182 24404
rect 47578 24392 47584 24404
rect 47176 24364 47584 24392
rect 47176 24352 47182 24364
rect 47578 24352 47584 24364
rect 47636 24352 47642 24404
rect 48222 24352 48228 24404
rect 48280 24392 48286 24404
rect 48593 24395 48651 24401
rect 48280 24352 48314 24392
rect 48593 24361 48605 24395
rect 48639 24392 48651 24395
rect 48866 24392 48872 24404
rect 48639 24364 48872 24392
rect 48639 24361 48651 24364
rect 48593 24355 48651 24361
rect 48866 24352 48872 24364
rect 48924 24352 48930 24404
rect 48958 24352 48964 24404
rect 49016 24392 49022 24404
rect 49421 24395 49479 24401
rect 49421 24392 49433 24395
rect 49016 24364 49433 24392
rect 49016 24352 49022 24364
rect 49421 24361 49433 24364
rect 49467 24361 49479 24395
rect 49421 24355 49479 24361
rect 51718 24352 51724 24404
rect 51776 24352 51782 24404
rect 51810 24352 51816 24404
rect 51868 24352 51874 24404
rect 52086 24352 52092 24404
rect 52144 24392 52150 24404
rect 56686 24392 56692 24404
rect 52144 24364 56692 24392
rect 52144 24352 52150 24364
rect 56686 24352 56692 24364
rect 56744 24352 56750 24404
rect 57054 24352 57060 24404
rect 57112 24352 57118 24404
rect 57882 24352 57888 24404
rect 57940 24352 57946 24404
rect 13648 24256 13676 24352
rect 13814 24284 13820 24336
rect 13872 24284 13878 24336
rect 40052 24324 40080 24352
rect 43717 24327 43775 24333
rect 43717 24324 43729 24327
rect 39592 24296 40080 24324
rect 42720 24296 43729 24324
rect 12452 24228 13676 24256
rect 12452 24197 12480 24228
rect 12437 24191 12495 24197
rect 12437 24157 12449 24191
rect 12483 24157 12495 24191
rect 12437 24151 12495 24157
rect 12529 24191 12587 24197
rect 12529 24157 12541 24191
rect 12575 24157 12587 24191
rect 12529 24151 12587 24157
rect 10459 24092 12020 24120
rect 12161 24123 12219 24129
rect 10459 24089 10471 24092
rect 10413 24083 10471 24089
rect 12161 24089 12173 24123
rect 12207 24089 12219 24123
rect 12161 24083 12219 24089
rect 7484 24024 7696 24052
rect 6733 24015 6791 24021
rect 9766 24012 9772 24064
rect 9824 24012 9830 24064
rect 10229 24055 10287 24061
rect 10229 24021 10241 24055
rect 10275 24052 10287 24055
rect 10318 24052 10324 24064
rect 10275 24024 10324 24052
rect 10275 24021 10287 24024
rect 10229 24015 10287 24021
rect 10318 24012 10324 24024
rect 10376 24012 10382 24064
rect 10594 24012 10600 24064
rect 10652 24052 10658 24064
rect 11422 24052 11428 24064
rect 10652 24024 11428 24052
rect 10652 24012 10658 24024
rect 11422 24012 11428 24024
rect 11480 24052 11486 24064
rect 12176 24052 12204 24083
rect 12544 24064 12572 24151
rect 12710 24148 12716 24200
rect 12768 24148 12774 24200
rect 12894 24148 12900 24200
rect 12952 24188 12958 24200
rect 13354 24188 13360 24200
rect 12952 24160 13360 24188
rect 12952 24148 12958 24160
rect 13354 24148 13360 24160
rect 13412 24188 13418 24200
rect 13449 24191 13507 24197
rect 13449 24188 13461 24191
rect 13412 24160 13461 24188
rect 13412 24148 13418 24160
rect 13449 24157 13461 24160
rect 13495 24157 13507 24191
rect 13449 24151 13507 24157
rect 13541 24191 13599 24197
rect 13541 24157 13553 24191
rect 13587 24157 13599 24191
rect 13648 24188 13676 24228
rect 34514 24216 34520 24268
rect 34572 24256 34578 24268
rect 35069 24259 35127 24265
rect 35069 24256 35081 24259
rect 34572 24228 35081 24256
rect 34572 24216 34578 24228
rect 35069 24225 35081 24228
rect 35115 24256 35127 24259
rect 35161 24259 35219 24265
rect 35161 24256 35173 24259
rect 35115 24228 35173 24256
rect 35115 24225 35127 24228
rect 35069 24219 35127 24225
rect 35161 24225 35173 24228
rect 35207 24256 35219 24259
rect 35434 24256 35440 24268
rect 35207 24228 35440 24256
rect 35207 24225 35219 24228
rect 35161 24219 35219 24225
rect 35434 24216 35440 24228
rect 35492 24216 35498 24268
rect 36909 24259 36967 24265
rect 36909 24225 36921 24259
rect 36955 24256 36967 24259
rect 37826 24256 37832 24268
rect 36955 24228 37832 24256
rect 36955 24225 36967 24228
rect 36909 24219 36967 24225
rect 37826 24216 37832 24228
rect 37884 24256 37890 24268
rect 38289 24259 38347 24265
rect 38289 24256 38301 24259
rect 37884 24228 38301 24256
rect 37884 24216 37890 24228
rect 38289 24225 38301 24228
rect 38335 24225 38347 24259
rect 38289 24219 38347 24225
rect 13817 24191 13875 24197
rect 13817 24188 13829 24191
rect 13648 24160 13829 24188
rect 13541 24151 13599 24157
rect 13817 24157 13829 24160
rect 13863 24157 13875 24191
rect 13817 24151 13875 24157
rect 12618 24080 12624 24132
rect 12676 24120 12682 24132
rect 12986 24120 12992 24132
rect 12676 24092 12992 24120
rect 12676 24080 12682 24092
rect 12986 24080 12992 24092
rect 13044 24120 13050 24132
rect 13173 24123 13231 24129
rect 13173 24120 13185 24123
rect 13044 24092 13185 24120
rect 13044 24080 13050 24092
rect 13173 24089 13185 24092
rect 13219 24089 13231 24123
rect 13173 24083 13231 24089
rect 11480 24024 12204 24052
rect 11480 24012 11486 24024
rect 12526 24012 12532 24064
rect 12584 24012 12590 24064
rect 12710 24012 12716 24064
rect 12768 24052 12774 24064
rect 13556 24052 13584 24151
rect 37550 24148 37556 24200
rect 37608 24148 37614 24200
rect 38562 24148 38568 24200
rect 38620 24148 38626 24200
rect 39114 24148 39120 24200
rect 39172 24148 39178 24200
rect 39209 24191 39267 24197
rect 39209 24157 39221 24191
rect 39255 24157 39267 24191
rect 39209 24151 39267 24157
rect 35434 24080 35440 24132
rect 35492 24080 35498 24132
rect 35894 24080 35900 24132
rect 35952 24080 35958 24132
rect 38580 24120 38608 24148
rect 39224 24120 39252 24151
rect 39390 24148 39396 24200
rect 39448 24148 39454 24200
rect 39485 24191 39543 24197
rect 39485 24157 39497 24191
rect 39531 24157 39543 24191
rect 39592 24188 39620 24296
rect 42150 24216 42156 24268
rect 42208 24256 42214 24268
rect 42720 24256 42748 24296
rect 43717 24293 43729 24296
rect 43763 24324 43775 24327
rect 44082 24324 44088 24336
rect 43763 24296 44088 24324
rect 43763 24293 43775 24296
rect 43717 24287 43775 24293
rect 44082 24284 44088 24296
rect 44140 24284 44146 24336
rect 44361 24327 44419 24333
rect 44361 24293 44373 24327
rect 44407 24324 44419 24327
rect 45020 24324 45048 24352
rect 44407 24296 45048 24324
rect 44407 24293 44419 24296
rect 44361 24287 44419 24293
rect 42208 24228 42748 24256
rect 42208 24216 42214 24228
rect 42720 24200 42748 24228
rect 43073 24259 43131 24265
rect 43073 24225 43085 24259
rect 43119 24256 43131 24259
rect 43119 24228 43300 24256
rect 43119 24225 43131 24228
rect 43073 24219 43131 24225
rect 39669 24191 39727 24197
rect 39669 24188 39681 24191
rect 39592 24160 39681 24188
rect 39485 24151 39543 24157
rect 39669 24157 39681 24160
rect 39715 24157 39727 24191
rect 39669 24151 39727 24157
rect 38580 24092 39252 24120
rect 39500 24120 39528 24151
rect 39758 24148 39764 24200
rect 39816 24188 39822 24200
rect 39853 24191 39911 24197
rect 39853 24188 39865 24191
rect 39816 24160 39865 24188
rect 39816 24148 39822 24160
rect 39853 24157 39865 24160
rect 39899 24188 39911 24191
rect 39899 24160 40080 24188
rect 39899 24157 39911 24160
rect 39853 24151 39911 24157
rect 39945 24123 40003 24129
rect 39945 24120 39957 24123
rect 39500 24092 39957 24120
rect 39945 24089 39957 24092
rect 39991 24089 40003 24123
rect 39945 24083 40003 24089
rect 12768 24024 13584 24052
rect 12768 24012 12774 24024
rect 13630 24012 13636 24064
rect 13688 24012 13694 24064
rect 36998 24012 37004 24064
rect 37056 24012 37062 24064
rect 38378 24012 38384 24064
rect 38436 24052 38442 24064
rect 38473 24055 38531 24061
rect 38473 24052 38485 24055
rect 38436 24024 38485 24052
rect 38436 24012 38442 24024
rect 38473 24021 38485 24024
rect 38519 24021 38531 24055
rect 38473 24015 38531 24021
rect 39301 24055 39359 24061
rect 39301 24021 39313 24055
rect 39347 24052 39359 24055
rect 40052 24052 40080 24160
rect 41322 24148 41328 24200
rect 41380 24148 41386 24200
rect 42702 24148 42708 24200
rect 42760 24148 42766 24200
rect 43272 24197 43300 24228
rect 43898 24216 43904 24268
rect 43956 24256 43962 24268
rect 43956 24228 44680 24256
rect 43956 24216 43962 24228
rect 44652 24197 44680 24228
rect 45020 24197 45048 24296
rect 43257 24191 43315 24197
rect 43257 24157 43269 24191
rect 43303 24188 43315 24191
rect 44637 24191 44695 24197
rect 43303 24160 44312 24188
rect 43303 24157 43315 24160
rect 43257 24151 43315 24157
rect 41598 24080 41604 24132
rect 41656 24080 41662 24132
rect 43898 24080 43904 24132
rect 43956 24120 43962 24132
rect 43993 24123 44051 24129
rect 43993 24120 44005 24123
rect 43956 24092 44005 24120
rect 43956 24080 43962 24092
rect 43993 24089 44005 24092
rect 44039 24089 44051 24123
rect 43993 24083 44051 24089
rect 44082 24080 44088 24132
rect 44140 24120 44146 24132
rect 44177 24123 44235 24129
rect 44177 24120 44189 24123
rect 44140 24092 44189 24120
rect 44140 24080 44146 24092
rect 44177 24089 44189 24092
rect 44223 24089 44235 24123
rect 44177 24083 44235 24089
rect 44284 24064 44312 24160
rect 44637 24157 44649 24191
rect 44683 24157 44695 24191
rect 44637 24151 44695 24157
rect 45005 24191 45063 24197
rect 45005 24157 45017 24191
rect 45051 24157 45063 24191
rect 45005 24151 45063 24157
rect 39347 24024 40080 24052
rect 39347 24021 39359 24024
rect 39301 24015 39359 24021
rect 43438 24012 43444 24064
rect 43496 24012 43502 24064
rect 44266 24012 44272 24064
rect 44324 24012 44330 24064
rect 44652 24052 44680 24151
rect 45278 24148 45284 24200
rect 45336 24148 45342 24200
rect 45480 24197 45508 24352
rect 48286 24324 48314 24352
rect 49697 24327 49755 24333
rect 49697 24324 49709 24327
rect 47044 24296 48176 24324
rect 48286 24296 49709 24324
rect 47044 24265 47072 24296
rect 48148 24268 48176 24296
rect 49697 24293 49709 24296
rect 49743 24324 49755 24327
rect 51626 24324 51632 24336
rect 49743 24296 51632 24324
rect 49743 24293 49755 24296
rect 49697 24287 49755 24293
rect 51626 24284 51632 24296
rect 51684 24284 51690 24336
rect 47029 24259 47087 24265
rect 47029 24225 47041 24259
rect 47075 24225 47087 24259
rect 47305 24259 47363 24265
rect 47305 24256 47317 24259
rect 47029 24219 47087 24225
rect 47136 24228 47317 24256
rect 45465 24191 45523 24197
rect 45465 24157 45477 24191
rect 45511 24157 45523 24191
rect 45465 24151 45523 24157
rect 45646 24148 45652 24200
rect 45704 24188 45710 24200
rect 47136 24197 47164 24228
rect 47305 24225 47317 24228
rect 47351 24225 47363 24259
rect 47305 24219 47363 24225
rect 48130 24216 48136 24268
rect 48188 24216 48194 24268
rect 48774 24216 48780 24268
rect 48832 24216 48838 24268
rect 51736 24256 51764 24352
rect 51276 24228 51764 24256
rect 51828 24256 51856 24352
rect 55030 24284 55036 24336
rect 55088 24324 55094 24336
rect 56137 24327 56195 24333
rect 55088 24296 56088 24324
rect 55088 24284 55094 24296
rect 51828 24228 54432 24256
rect 47121 24191 47179 24197
rect 47121 24188 47133 24191
rect 45704 24160 47133 24188
rect 45704 24148 45710 24160
rect 47121 24157 47133 24160
rect 47167 24157 47179 24191
rect 47121 24151 47179 24157
rect 47213 24191 47271 24197
rect 47213 24157 47225 24191
rect 47259 24157 47271 24191
rect 47213 24151 47271 24157
rect 47397 24191 47455 24197
rect 47397 24157 47409 24191
rect 47443 24188 47455 24191
rect 47670 24188 47676 24200
rect 47443 24160 47676 24188
rect 47443 24157 47455 24160
rect 47397 24151 47455 24157
rect 45094 24080 45100 24132
rect 45152 24080 45158 24132
rect 47228 24064 47256 24151
rect 47670 24148 47676 24160
rect 47728 24148 47734 24200
rect 48501 24191 48559 24197
rect 48501 24157 48513 24191
rect 48547 24157 48559 24191
rect 48501 24151 48559 24157
rect 47486 24080 47492 24132
rect 47544 24120 47550 24132
rect 48516 24120 48544 24151
rect 48590 24148 48596 24200
rect 48648 24188 48654 24200
rect 48685 24191 48743 24197
rect 48685 24188 48697 24191
rect 48648 24160 48697 24188
rect 48648 24148 48654 24160
rect 48685 24157 48697 24160
rect 48731 24188 48743 24191
rect 48958 24188 48964 24200
rect 48731 24160 48964 24188
rect 48731 24157 48743 24160
rect 48685 24151 48743 24157
rect 48958 24148 48964 24160
rect 49016 24148 49022 24200
rect 49605 24191 49663 24197
rect 49605 24157 49617 24191
rect 49651 24188 49663 24191
rect 50614 24188 50620 24200
rect 49651 24160 50620 24188
rect 49651 24157 49663 24160
rect 49605 24151 49663 24157
rect 49620 24120 49648 24151
rect 50614 24148 50620 24160
rect 50672 24148 50678 24200
rect 51276 24197 51304 24228
rect 50801 24191 50859 24197
rect 50801 24157 50813 24191
rect 50847 24157 50859 24191
rect 50801 24151 50859 24157
rect 51261 24191 51319 24197
rect 51261 24157 51273 24191
rect 51307 24157 51319 24191
rect 51261 24151 51319 24157
rect 50816 24120 50844 24151
rect 51442 24148 51448 24200
rect 51500 24148 51506 24200
rect 51537 24191 51595 24197
rect 51537 24157 51549 24191
rect 51583 24157 51595 24191
rect 51537 24151 51595 24157
rect 51721 24191 51779 24197
rect 51721 24157 51733 24191
rect 51767 24188 51779 24191
rect 52270 24188 52276 24200
rect 51767 24160 52276 24188
rect 51767 24157 51779 24160
rect 51721 24151 51779 24157
rect 51074 24120 51080 24132
rect 47544 24092 48314 24120
rect 48516 24092 49648 24120
rect 49712 24092 50752 24120
rect 50816 24092 51080 24120
rect 47544 24080 47550 24092
rect 46753 24055 46811 24061
rect 46753 24052 46765 24055
rect 44652 24024 46765 24052
rect 46753 24021 46765 24024
rect 46799 24021 46811 24055
rect 46753 24015 46811 24021
rect 47210 24012 47216 24064
rect 47268 24012 47274 24064
rect 47670 24012 47676 24064
rect 47728 24052 47734 24064
rect 47765 24055 47823 24061
rect 47765 24052 47777 24055
rect 47728 24024 47777 24052
rect 47728 24012 47734 24024
rect 47765 24021 47777 24024
rect 47811 24052 47823 24055
rect 48130 24052 48136 24064
rect 47811 24024 48136 24052
rect 47811 24021 47823 24024
rect 47765 24015 47823 24021
rect 48130 24012 48136 24024
rect 48188 24012 48194 24064
rect 48286 24052 48314 24092
rect 49712 24052 49740 24092
rect 50724 24064 50752 24092
rect 51074 24080 51080 24092
rect 51132 24120 51138 24132
rect 51552 24120 51580 24151
rect 52270 24148 52276 24160
rect 52328 24148 52334 24200
rect 52825 24191 52883 24197
rect 52825 24157 52837 24191
rect 52871 24157 52883 24191
rect 52825 24151 52883 24157
rect 53009 24191 53067 24197
rect 53009 24157 53021 24191
rect 53055 24188 53067 24191
rect 53282 24188 53288 24200
rect 53055 24160 53288 24188
rect 53055 24157 53067 24160
rect 53009 24151 53067 24157
rect 52840 24120 52868 24151
rect 53282 24148 53288 24160
rect 53340 24148 53346 24200
rect 53374 24148 53380 24200
rect 53432 24148 53438 24200
rect 53392 24120 53420 24148
rect 51132 24092 53420 24120
rect 54404 24120 54432 24228
rect 55950 24216 55956 24268
rect 56008 24216 56014 24268
rect 56060 24256 56088 24296
rect 56137 24293 56149 24327
rect 56183 24324 56195 24327
rect 56226 24324 56232 24336
rect 56183 24296 56232 24324
rect 56183 24293 56195 24296
rect 56137 24287 56195 24293
rect 56226 24284 56232 24296
rect 56284 24284 56290 24336
rect 57072 24256 57100 24352
rect 56060 24228 56180 24256
rect 54849 24191 54907 24197
rect 54849 24157 54861 24191
rect 54895 24188 54907 24191
rect 56045 24191 56103 24197
rect 54895 24160 55352 24188
rect 54895 24157 54907 24160
rect 54849 24151 54907 24157
rect 55324 24129 55352 24160
rect 56045 24157 56057 24191
rect 56091 24157 56103 24191
rect 56045 24151 56103 24157
rect 55309 24123 55367 24129
rect 54404 24092 54892 24120
rect 51132 24080 51138 24092
rect 48286 24024 49740 24052
rect 50614 24012 50620 24064
rect 50672 24012 50678 24064
rect 50706 24012 50712 24064
rect 50764 24012 50770 24064
rect 51350 24012 51356 24064
rect 51408 24012 51414 24064
rect 51721 24055 51779 24061
rect 51721 24021 51733 24055
rect 51767 24052 51779 24055
rect 51902 24052 51908 24064
rect 51767 24024 51908 24052
rect 51767 24021 51779 24024
rect 51721 24015 51779 24021
rect 51902 24012 51908 24024
rect 51960 24012 51966 24064
rect 52914 24012 52920 24064
rect 52972 24012 52978 24064
rect 54202 24012 54208 24064
rect 54260 24052 54266 24064
rect 54757 24055 54815 24061
rect 54757 24052 54769 24055
rect 54260 24024 54769 24052
rect 54260 24012 54266 24024
rect 54757 24021 54769 24024
rect 54803 24021 54815 24055
rect 54864 24052 54892 24092
rect 55309 24089 55321 24123
rect 55355 24120 55367 24123
rect 56060 24120 56088 24151
rect 55355 24092 56088 24120
rect 56152 24120 56180 24228
rect 56888 24228 57100 24256
rect 56229 24191 56287 24197
rect 56229 24157 56241 24191
rect 56275 24188 56287 24191
rect 56502 24188 56508 24200
rect 56275 24160 56508 24188
rect 56275 24157 56287 24160
rect 56229 24151 56287 24157
rect 56502 24148 56508 24160
rect 56560 24148 56566 24200
rect 56888 24197 56916 24228
rect 56873 24191 56931 24197
rect 56873 24157 56885 24191
rect 56919 24157 56931 24191
rect 56873 24151 56931 24157
rect 57057 24191 57115 24197
rect 57057 24157 57069 24191
rect 57103 24188 57115 24191
rect 57422 24188 57428 24200
rect 57103 24160 57428 24188
rect 57103 24157 57115 24160
rect 57057 24151 57115 24157
rect 57422 24148 57428 24160
rect 57480 24148 57486 24200
rect 57900 24197 57928 24352
rect 57885 24191 57943 24197
rect 57885 24157 57897 24191
rect 57931 24157 57943 24191
rect 57885 24151 57943 24157
rect 58158 24148 58164 24200
rect 58216 24148 58222 24200
rect 58253 24123 58311 24129
rect 58253 24120 58265 24123
rect 56152 24092 58265 24120
rect 55355 24089 55367 24092
rect 55309 24083 55367 24089
rect 58253 24089 58265 24092
rect 58299 24089 58311 24123
rect 58253 24083 58311 24089
rect 56873 24055 56931 24061
rect 56873 24052 56885 24055
rect 54864 24024 56885 24052
rect 54757 24015 54815 24021
rect 56873 24021 56885 24024
rect 56919 24021 56931 24055
rect 56873 24015 56931 24021
rect 57974 24012 57980 24064
rect 58032 24012 58038 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 2682 23808 2688 23860
rect 2740 23808 2746 23860
rect 3234 23808 3240 23860
rect 3292 23808 3298 23860
rect 3973 23851 4031 23857
rect 3973 23817 3985 23851
rect 4019 23848 4031 23851
rect 4338 23848 4344 23860
rect 4019 23820 4344 23848
rect 4019 23817 4031 23820
rect 3973 23811 4031 23817
rect 4338 23808 4344 23820
rect 4396 23808 4402 23860
rect 4890 23808 4896 23860
rect 4948 23808 4954 23860
rect 7282 23808 7288 23860
rect 7340 23808 7346 23860
rect 7650 23808 7656 23860
rect 7708 23808 7714 23860
rect 7926 23808 7932 23860
rect 7984 23808 7990 23860
rect 8021 23851 8079 23857
rect 8021 23817 8033 23851
rect 8067 23848 8079 23851
rect 8202 23848 8208 23860
rect 8067 23820 8208 23848
rect 8067 23817 8079 23820
rect 8021 23811 8079 23817
rect 8202 23808 8208 23820
rect 8260 23808 8266 23860
rect 8478 23808 8484 23860
rect 8536 23808 8542 23860
rect 10042 23808 10048 23860
rect 10100 23808 10106 23860
rect 10134 23808 10140 23860
rect 10192 23808 10198 23860
rect 10502 23808 10508 23860
rect 10560 23808 10566 23860
rect 11330 23808 11336 23860
rect 11388 23848 11394 23860
rect 12250 23848 12256 23860
rect 11388 23820 12256 23848
rect 11388 23808 11394 23820
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 12897 23851 12955 23857
rect 12897 23817 12909 23851
rect 12943 23848 12955 23851
rect 13630 23848 13636 23860
rect 12943 23820 13636 23848
rect 12943 23817 12955 23820
rect 12897 23811 12955 23817
rect 13630 23808 13636 23820
rect 13688 23808 13694 23860
rect 13814 23808 13820 23860
rect 13872 23808 13878 23860
rect 35434 23808 35440 23860
rect 35492 23848 35498 23860
rect 35713 23851 35771 23857
rect 35713 23848 35725 23851
rect 35492 23820 35725 23848
rect 35492 23808 35498 23820
rect 35713 23817 35725 23820
rect 35759 23817 35771 23851
rect 36998 23848 37004 23860
rect 35713 23811 35771 23817
rect 36556 23820 37004 23848
rect 2700 23721 2728 23808
rect 3252 23780 3280 23808
rect 4157 23783 4215 23789
rect 4157 23780 4169 23783
rect 3252 23752 4169 23780
rect 4157 23749 4169 23752
rect 4203 23749 4215 23783
rect 4908 23780 4936 23808
rect 5454 23783 5512 23789
rect 5454 23780 5466 23783
rect 4908 23752 5466 23780
rect 4157 23743 4215 23749
rect 5454 23749 5466 23752
rect 5500 23749 5512 23783
rect 5454 23743 5512 23749
rect 2685 23715 2743 23721
rect 2685 23681 2697 23715
rect 2731 23681 2743 23715
rect 2685 23675 2743 23681
rect 3329 23715 3387 23721
rect 3329 23681 3341 23715
rect 3375 23712 3387 23715
rect 3789 23715 3847 23721
rect 3789 23712 3801 23715
rect 3375 23684 3801 23712
rect 3375 23681 3387 23684
rect 3329 23675 3387 23681
rect 3789 23681 3801 23684
rect 3835 23681 3847 23715
rect 3789 23675 3847 23681
rect 3970 23672 3976 23724
rect 4028 23672 4034 23724
rect 4062 23672 4068 23724
rect 4120 23672 4126 23724
rect 4249 23715 4307 23721
rect 4249 23681 4261 23715
rect 4295 23681 4307 23715
rect 4249 23675 4307 23681
rect 5721 23715 5779 23721
rect 5721 23681 5733 23715
rect 5767 23712 5779 23715
rect 7300 23712 7328 23808
rect 7500 23783 7558 23789
rect 7500 23749 7512 23783
rect 7546 23780 7558 23783
rect 7668 23780 7696 23808
rect 7546 23752 7696 23780
rect 7944 23780 7972 23808
rect 8380 23783 8438 23789
rect 7944 23752 8064 23780
rect 7546 23749 7558 23752
rect 7500 23743 7558 23749
rect 8036 23721 8064 23752
rect 8380 23749 8392 23783
rect 8426 23780 8438 23783
rect 8496 23780 8524 23808
rect 8426 23752 8524 23780
rect 10060 23780 10088 23808
rect 12158 23780 12164 23792
rect 10060 23752 10364 23780
rect 8426 23749 8438 23752
rect 8380 23743 8438 23749
rect 7745 23715 7803 23721
rect 7745 23712 7757 23715
rect 5767 23684 7757 23712
rect 5767 23681 5779 23684
rect 5721 23675 5779 23681
rect 7745 23681 7757 23684
rect 7791 23681 7803 23715
rect 7745 23675 7803 23681
rect 7837 23715 7895 23721
rect 7837 23681 7849 23715
rect 7883 23712 7895 23715
rect 8021 23715 8079 23721
rect 7883 23684 7972 23712
rect 7883 23681 7895 23684
rect 7837 23675 7895 23681
rect 3878 23604 3884 23656
rect 3936 23644 3942 23656
rect 4080 23644 4108 23672
rect 3936 23616 4108 23644
rect 3936 23604 3942 23616
rect 4264 23576 4292 23675
rect 4264 23548 4844 23576
rect 4816 23520 4844 23548
rect 7944 23520 7972 23684
rect 8021 23681 8033 23715
rect 8067 23712 8079 23715
rect 10134 23712 10140 23724
rect 8067 23684 10140 23712
rect 8067 23681 8079 23684
rect 8021 23675 8079 23681
rect 10134 23672 10140 23684
rect 10192 23672 10198 23724
rect 10336 23721 10364 23752
rect 11900 23752 12164 23780
rect 10321 23715 10379 23721
rect 10321 23681 10333 23715
rect 10367 23681 10379 23715
rect 10321 23675 10379 23681
rect 10413 23715 10471 23721
rect 10413 23681 10425 23715
rect 10459 23712 10471 23715
rect 10962 23712 10968 23724
rect 10459 23684 10968 23712
rect 10459 23681 10471 23684
rect 10413 23675 10471 23681
rect 10962 23672 10968 23684
rect 11020 23672 11026 23724
rect 8110 23604 8116 23656
rect 8168 23604 8174 23656
rect 10152 23644 10180 23672
rect 11900 23644 11928 23752
rect 12158 23740 12164 23752
rect 12216 23780 12222 23792
rect 13832 23780 13860 23808
rect 14102 23783 14160 23789
rect 14102 23780 14114 23783
rect 12216 23752 12848 23780
rect 13832 23752 14114 23780
rect 12216 23740 12222 23752
rect 12820 23724 12848 23752
rect 14102 23749 14114 23752
rect 14148 23749 14160 23783
rect 14102 23743 14160 23749
rect 36449 23783 36507 23789
rect 36449 23749 36461 23783
rect 36495 23749 36507 23783
rect 36449 23743 36507 23749
rect 12253 23715 12311 23721
rect 12253 23681 12265 23715
rect 12299 23712 12311 23715
rect 12713 23715 12771 23721
rect 12713 23712 12725 23715
rect 12299 23684 12725 23712
rect 12299 23681 12311 23684
rect 12253 23675 12311 23681
rect 12713 23681 12725 23684
rect 12759 23681 12771 23715
rect 12713 23675 12771 23681
rect 10152 23616 11928 23644
rect 11974 23604 11980 23656
rect 12032 23604 12038 23656
rect 12728 23644 12756 23675
rect 12802 23672 12808 23724
rect 12860 23712 12866 23724
rect 12897 23715 12955 23721
rect 12897 23712 12909 23715
rect 12860 23684 12909 23712
rect 12860 23672 12866 23684
rect 12897 23681 12909 23684
rect 12943 23681 12955 23715
rect 12897 23675 12955 23681
rect 12986 23672 12992 23724
rect 13044 23712 13050 23724
rect 14369 23715 14427 23721
rect 14369 23712 14381 23715
rect 13044 23684 14381 23712
rect 13044 23672 13050 23684
rect 14369 23681 14381 23684
rect 14415 23681 14427 23715
rect 14369 23675 14427 23681
rect 36357 23715 36415 23721
rect 36357 23681 36369 23715
rect 36403 23712 36415 23715
rect 36464 23712 36492 23743
rect 36403 23684 36492 23712
rect 36403 23681 36415 23684
rect 36357 23675 36415 23681
rect 36449 23647 36507 23653
rect 12728 23616 13032 23644
rect 12161 23579 12219 23585
rect 12161 23576 12173 23579
rect 11900 23548 12173 23576
rect 11900 23520 11928 23548
rect 12161 23545 12173 23548
rect 12207 23545 12219 23579
rect 12161 23539 12219 23545
rect 12250 23536 12256 23588
rect 12308 23576 12314 23588
rect 12618 23576 12624 23588
rect 12308 23548 12624 23576
rect 12308 23536 12314 23548
rect 12618 23536 12624 23548
rect 12676 23536 12682 23588
rect 13004 23585 13032 23616
rect 36449 23613 36461 23647
rect 36495 23644 36507 23647
rect 36556 23644 36584 23820
rect 36998 23808 37004 23820
rect 37056 23808 37062 23860
rect 37274 23808 37280 23860
rect 37332 23808 37338 23860
rect 38010 23848 38016 23860
rect 37384 23820 38016 23848
rect 37292 23780 37320 23808
rect 36740 23752 37320 23780
rect 36740 23721 36768 23752
rect 36725 23715 36783 23721
rect 36725 23681 36737 23715
rect 36771 23681 36783 23715
rect 36725 23675 36783 23681
rect 36814 23672 36820 23724
rect 36872 23672 36878 23724
rect 37001 23715 37059 23721
rect 37001 23681 37013 23715
rect 37047 23712 37059 23715
rect 37090 23712 37096 23724
rect 37047 23684 37096 23712
rect 37047 23681 37059 23684
rect 37001 23675 37059 23681
rect 36495 23616 36584 23644
rect 36495 23613 36507 23616
rect 36449 23607 36507 23613
rect 12989 23579 13047 23585
rect 12989 23545 13001 23579
rect 13035 23545 13047 23579
rect 12989 23539 13047 23545
rect 36633 23579 36691 23585
rect 36633 23545 36645 23579
rect 36679 23576 36691 23579
rect 37016 23576 37044 23675
rect 37090 23672 37096 23684
rect 37148 23672 37154 23724
rect 37384 23721 37412 23820
rect 38010 23808 38016 23820
rect 38068 23808 38074 23860
rect 38378 23808 38384 23860
rect 38436 23808 38442 23860
rect 38470 23808 38476 23860
rect 38528 23808 38534 23860
rect 38562 23808 38568 23860
rect 38620 23808 38626 23860
rect 39114 23808 39120 23860
rect 39172 23848 39178 23860
rect 39577 23851 39635 23857
rect 39577 23848 39589 23851
rect 39172 23820 39589 23848
rect 39172 23808 39178 23820
rect 39577 23817 39589 23820
rect 39623 23817 39635 23851
rect 39577 23811 39635 23817
rect 41598 23808 41604 23860
rect 41656 23848 41662 23860
rect 42429 23851 42487 23857
rect 42429 23848 42441 23851
rect 41656 23820 42441 23848
rect 41656 23808 41662 23820
rect 42429 23817 42441 23820
rect 42475 23817 42487 23851
rect 42429 23811 42487 23817
rect 43806 23808 43812 23860
rect 43864 23848 43870 23860
rect 44085 23851 44143 23857
rect 44085 23848 44097 23851
rect 43864 23820 44097 23848
rect 43864 23808 43870 23820
rect 44085 23817 44097 23820
rect 44131 23817 44143 23851
rect 44085 23811 44143 23817
rect 49786 23808 49792 23860
rect 49844 23848 49850 23860
rect 50522 23848 50528 23860
rect 49844 23820 50528 23848
rect 49844 23808 49850 23820
rect 50522 23808 50528 23820
rect 50580 23808 50586 23860
rect 50614 23808 50620 23860
rect 50672 23808 50678 23860
rect 53834 23808 53840 23860
rect 53892 23808 53898 23860
rect 54846 23808 54852 23860
rect 54904 23848 54910 23860
rect 54904 23820 55168 23848
rect 54904 23808 54910 23820
rect 37645 23783 37703 23789
rect 37645 23749 37657 23783
rect 37691 23780 37703 23783
rect 37691 23752 38332 23780
rect 37691 23749 37703 23752
rect 37645 23743 37703 23749
rect 38304 23721 38332 23752
rect 37369 23715 37427 23721
rect 37369 23681 37381 23715
rect 37415 23681 37427 23715
rect 37369 23675 37427 23681
rect 38289 23715 38347 23721
rect 38289 23681 38301 23715
rect 38335 23681 38347 23715
rect 38289 23675 38347 23681
rect 37645 23647 37703 23653
rect 37645 23613 37657 23647
rect 37691 23644 37703 23647
rect 38396 23644 38424 23808
rect 38473 23715 38531 23721
rect 38473 23681 38485 23715
rect 38519 23712 38531 23715
rect 38580 23712 38608 23808
rect 38841 23783 38899 23789
rect 38841 23780 38853 23783
rect 38672 23752 38853 23780
rect 38672 23721 38700 23752
rect 38841 23749 38853 23752
rect 38887 23780 38899 23783
rect 39390 23780 39396 23792
rect 38887 23752 39396 23780
rect 38887 23749 38899 23752
rect 38841 23743 38899 23749
rect 39390 23740 39396 23752
rect 39448 23780 39454 23792
rect 39448 23752 39804 23780
rect 39448 23740 39454 23752
rect 39776 23721 39804 23752
rect 43438 23740 43444 23792
rect 43496 23780 43502 23792
rect 50632 23780 50660 23808
rect 43496 23752 44312 23780
rect 43496 23740 43502 23752
rect 43916 23721 43944 23752
rect 38519 23684 38608 23712
rect 38657 23715 38715 23721
rect 38519 23681 38531 23684
rect 38473 23675 38531 23681
rect 38657 23681 38669 23715
rect 38703 23681 38715 23715
rect 38657 23675 38715 23681
rect 39577 23715 39635 23721
rect 39577 23681 39589 23715
rect 39623 23681 39635 23715
rect 39577 23675 39635 23681
rect 39761 23715 39819 23721
rect 39761 23681 39773 23715
rect 39807 23681 39819 23715
rect 39761 23675 39819 23681
rect 43349 23715 43407 23721
rect 43349 23681 43361 23715
rect 43395 23712 43407 23715
rect 43717 23715 43775 23721
rect 43717 23712 43729 23715
rect 43395 23684 43729 23712
rect 43395 23681 43407 23684
rect 43349 23675 43407 23681
rect 43717 23681 43729 23684
rect 43763 23681 43775 23715
rect 43717 23675 43775 23681
rect 43901 23715 43959 23721
rect 43901 23681 43913 23715
rect 43947 23681 43959 23715
rect 43901 23675 43959 23681
rect 37691 23616 38424 23644
rect 37691 23613 37703 23616
rect 37645 23607 37703 23613
rect 39390 23604 39396 23656
rect 39448 23604 39454 23656
rect 37461 23579 37519 23585
rect 37461 23576 37473 23579
rect 36679 23548 37473 23576
rect 36679 23545 36691 23548
rect 36633 23539 36691 23545
rect 37461 23545 37473 23548
rect 37507 23576 37519 23579
rect 39592 23576 39620 23675
rect 43990 23672 43996 23724
rect 44048 23712 44054 23724
rect 44284 23721 44312 23752
rect 48148 23752 50660 23780
rect 48148 23721 48176 23752
rect 44177 23715 44235 23721
rect 44177 23712 44189 23715
rect 44048 23684 44189 23712
rect 44048 23672 44054 23684
rect 44177 23681 44189 23684
rect 44223 23681 44235 23715
rect 44177 23675 44235 23681
rect 44269 23715 44327 23721
rect 44269 23681 44281 23715
rect 44315 23681 44327 23715
rect 44269 23675 44327 23681
rect 47949 23715 48007 23721
rect 47949 23681 47961 23715
rect 47995 23681 48007 23715
rect 47949 23675 48007 23681
rect 48133 23715 48191 23721
rect 48133 23681 48145 23715
rect 48179 23681 48191 23715
rect 48133 23675 48191 23681
rect 41325 23647 41383 23653
rect 41325 23613 41337 23647
rect 41371 23644 41383 23647
rect 41509 23647 41567 23653
rect 41509 23644 41521 23647
rect 41371 23616 41521 23644
rect 41371 23613 41383 23616
rect 41325 23607 41383 23613
rect 41509 23613 41521 23616
rect 41555 23613 41567 23647
rect 41509 23607 41567 23613
rect 42153 23647 42211 23653
rect 42153 23613 42165 23647
rect 42199 23644 42211 23647
rect 42242 23644 42248 23656
rect 42199 23616 42248 23644
rect 42199 23613 42211 23616
rect 42153 23607 42211 23613
rect 42242 23604 42248 23616
rect 42300 23604 42306 23656
rect 43073 23647 43131 23653
rect 43073 23613 43085 23647
rect 43119 23644 43131 23647
rect 43165 23647 43223 23653
rect 43165 23644 43177 23647
rect 43119 23616 43177 23644
rect 43119 23613 43131 23616
rect 43073 23607 43131 23613
rect 43165 23613 43177 23616
rect 43211 23613 43223 23647
rect 43165 23607 43223 23613
rect 43625 23647 43683 23653
rect 43625 23613 43637 23647
rect 43671 23644 43683 23647
rect 44361 23647 44419 23653
rect 44361 23644 44373 23647
rect 43671 23616 44373 23644
rect 43671 23613 43683 23616
rect 43625 23607 43683 23613
rect 44361 23613 44373 23616
rect 44407 23613 44419 23647
rect 44361 23607 44419 23613
rect 46566 23604 46572 23656
rect 46624 23604 46630 23656
rect 47964 23644 47992 23675
rect 48958 23672 48964 23724
rect 49016 23712 49022 23724
rect 50264 23721 50292 23752
rect 52822 23740 52828 23792
rect 52880 23780 52886 23792
rect 53852 23780 53880 23808
rect 54757 23783 54815 23789
rect 54757 23780 54769 23783
rect 52880 23752 53328 23780
rect 53852 23752 54432 23780
rect 52880 23740 52886 23752
rect 49973 23715 50031 23721
rect 49973 23712 49985 23715
rect 49016 23684 49985 23712
rect 49016 23672 49022 23684
rect 49973 23681 49985 23684
rect 50019 23681 50031 23715
rect 49973 23675 50031 23681
rect 50157 23715 50215 23721
rect 50157 23681 50169 23715
rect 50203 23681 50215 23715
rect 50157 23675 50215 23681
rect 50249 23715 50307 23721
rect 50249 23681 50261 23715
rect 50295 23681 50307 23715
rect 50427 23715 50485 23721
rect 50427 23712 50439 23715
rect 50249 23675 50307 23681
rect 50356 23684 50439 23712
rect 49605 23647 49663 23653
rect 49605 23644 49617 23647
rect 47964 23616 49617 23644
rect 49605 23613 49617 23616
rect 49651 23613 49663 23647
rect 49605 23607 49663 23613
rect 37507 23548 39620 23576
rect 41049 23579 41107 23585
rect 37507 23545 37519 23548
rect 37461 23539 37519 23545
rect 41049 23545 41061 23579
rect 41095 23576 41107 23579
rect 44634 23576 44640 23588
rect 41095 23548 44640 23576
rect 41095 23545 41107 23548
rect 41049 23539 41107 23545
rect 44634 23536 44640 23548
rect 44692 23536 44698 23588
rect 49620 23576 49648 23607
rect 49786 23604 49792 23656
rect 49844 23644 49850 23656
rect 49881 23647 49939 23653
rect 49881 23644 49893 23647
rect 49844 23616 49893 23644
rect 49844 23604 49850 23616
rect 49881 23613 49893 23616
rect 49927 23613 49939 23647
rect 49881 23607 49939 23613
rect 50062 23604 50068 23656
rect 50120 23604 50126 23656
rect 50172 23644 50200 23675
rect 50356 23644 50384 23684
rect 50427 23681 50439 23684
rect 50473 23681 50485 23715
rect 50427 23675 50485 23681
rect 50522 23672 50528 23724
rect 50580 23672 50586 23724
rect 50709 23715 50767 23721
rect 50709 23681 50721 23715
rect 50755 23712 50767 23715
rect 50755 23684 51074 23712
rect 50755 23681 50767 23684
rect 50709 23675 50767 23681
rect 50172 23616 50384 23644
rect 51046 23644 51074 23684
rect 52730 23672 52736 23724
rect 52788 23672 52794 23724
rect 52914 23672 52920 23724
rect 52972 23672 52978 23724
rect 53300 23712 53328 23752
rect 54404 23724 54432 23752
rect 54588 23752 54769 23780
rect 53926 23712 53932 23724
rect 53300 23684 53932 23712
rect 53926 23672 53932 23684
rect 53984 23712 53990 23724
rect 54021 23715 54079 23721
rect 54021 23712 54033 23715
rect 53984 23684 54033 23712
rect 53984 23672 53990 23684
rect 54021 23681 54033 23684
rect 54067 23681 54079 23715
rect 54021 23675 54079 23681
rect 54202 23672 54208 23724
rect 54260 23672 54266 23724
rect 54294 23672 54300 23724
rect 54352 23672 54358 23724
rect 54386 23672 54392 23724
rect 54444 23672 54450 23724
rect 54588 23721 54616 23752
rect 54757 23749 54769 23752
rect 54803 23749 54815 23783
rect 54757 23743 54815 23749
rect 55140 23780 55168 23820
rect 57974 23808 57980 23860
rect 58032 23808 58038 23860
rect 57992 23780 58020 23808
rect 55140 23752 58020 23780
rect 54573 23715 54631 23721
rect 54573 23681 54585 23715
rect 54619 23681 54631 23715
rect 54573 23675 54631 23681
rect 54665 23715 54723 23721
rect 54665 23681 54677 23715
rect 54711 23681 54723 23715
rect 54665 23675 54723 23681
rect 54849 23715 54907 23721
rect 54849 23681 54861 23715
rect 54895 23681 54907 23715
rect 54849 23675 54907 23681
rect 52825 23647 52883 23653
rect 52825 23644 52837 23647
rect 51046 23616 52837 23644
rect 50172 23576 50200 23616
rect 52825 23613 52837 23616
rect 52871 23613 52883 23647
rect 54680 23644 54708 23675
rect 52825 23607 52883 23613
rect 54312 23616 54708 23644
rect 54864 23644 54892 23675
rect 54938 23672 54944 23724
rect 54996 23672 55002 23724
rect 55140 23721 55168 23752
rect 56502 23721 56508 23724
rect 55125 23715 55183 23721
rect 55125 23681 55137 23715
rect 55171 23681 55183 23715
rect 55125 23675 55183 23681
rect 56496 23675 56508 23721
rect 56502 23672 56508 23675
rect 56560 23672 56566 23724
rect 55033 23647 55091 23653
rect 55033 23644 55045 23647
rect 54864 23616 55045 23644
rect 50338 23576 50344 23588
rect 49620 23548 50344 23576
rect 50338 23536 50344 23548
rect 50396 23536 50402 23588
rect 50706 23536 50712 23588
rect 50764 23576 50770 23588
rect 54312 23585 54340 23616
rect 55033 23613 55045 23616
rect 55079 23613 55091 23647
rect 55033 23607 55091 23613
rect 56226 23604 56232 23656
rect 56284 23604 56290 23656
rect 58437 23647 58495 23653
rect 58437 23613 58449 23647
rect 58483 23613 58495 23647
rect 58437 23607 58495 23613
rect 54297 23579 54355 23585
rect 50764 23548 53972 23576
rect 50764 23536 50770 23548
rect 4341 23511 4399 23517
rect 4341 23477 4353 23511
rect 4387 23508 4399 23511
rect 4706 23508 4712 23520
rect 4387 23480 4712 23508
rect 4387 23477 4399 23480
rect 4341 23471 4399 23477
rect 4706 23468 4712 23480
rect 4764 23468 4770 23520
rect 4798 23468 4804 23520
rect 4856 23468 4862 23520
rect 6365 23511 6423 23517
rect 6365 23477 6377 23511
rect 6411 23508 6423 23511
rect 7006 23508 7012 23520
rect 6411 23480 7012 23508
rect 6411 23477 6423 23480
rect 6365 23471 6423 23477
rect 7006 23468 7012 23480
rect 7064 23468 7070 23520
rect 7926 23468 7932 23520
rect 7984 23508 7990 23520
rect 9493 23511 9551 23517
rect 9493 23508 9505 23511
rect 7984 23480 9505 23508
rect 7984 23468 7990 23480
rect 9493 23477 9505 23480
rect 9539 23477 9551 23511
rect 9493 23471 9551 23477
rect 10962 23468 10968 23520
rect 11020 23468 11026 23520
rect 11882 23468 11888 23520
rect 11940 23468 11946 23520
rect 12066 23468 12072 23520
rect 12124 23468 12130 23520
rect 12526 23468 12532 23520
rect 12584 23468 12590 23520
rect 36909 23511 36967 23517
rect 36909 23477 36921 23511
rect 36955 23508 36967 23511
rect 37550 23508 37556 23520
rect 36955 23480 37556 23508
rect 36955 23477 36967 23480
rect 36909 23471 36967 23477
rect 37550 23468 37556 23480
rect 37608 23468 37614 23520
rect 37734 23468 37740 23520
rect 37792 23468 37798 23520
rect 40862 23468 40868 23520
rect 40920 23468 40926 23520
rect 43533 23511 43591 23517
rect 43533 23477 43545 23511
rect 43579 23508 43591 23511
rect 44358 23508 44364 23520
rect 43579 23480 44364 23508
rect 43579 23477 43591 23480
rect 43533 23471 43591 23477
rect 44358 23468 44364 23480
rect 44416 23508 44422 23520
rect 45094 23508 45100 23520
rect 44416 23480 45100 23508
rect 44416 23468 44422 23480
rect 45094 23468 45100 23480
rect 45152 23468 45158 23520
rect 45922 23468 45928 23520
rect 45980 23468 45986 23520
rect 48038 23468 48044 23520
rect 48096 23468 48102 23520
rect 48590 23468 48596 23520
rect 48648 23508 48654 23520
rect 49326 23508 49332 23520
rect 48648 23480 49332 23508
rect 48648 23468 48654 23480
rect 49326 23468 49332 23480
rect 49384 23508 49390 23520
rect 50249 23511 50307 23517
rect 50249 23508 50261 23511
rect 49384 23480 50261 23508
rect 49384 23468 49390 23480
rect 50249 23477 50261 23480
rect 50295 23477 50307 23511
rect 50249 23471 50307 23477
rect 50614 23468 50620 23520
rect 50672 23468 50678 23520
rect 53944 23508 53972 23548
rect 54297 23545 54309 23579
rect 54343 23545 54355 23579
rect 57609 23579 57667 23585
rect 54297 23539 54355 23545
rect 54404 23548 54616 23576
rect 54404 23508 54432 23548
rect 53944 23480 54432 23508
rect 54478 23468 54484 23520
rect 54536 23468 54542 23520
rect 54588 23508 54616 23548
rect 57609 23545 57621 23579
rect 57655 23576 57667 23579
rect 58452 23576 58480 23607
rect 57655 23548 58480 23576
rect 57655 23545 57667 23548
rect 57609 23539 57667 23545
rect 56594 23508 56600 23520
rect 54588 23480 56600 23508
rect 56594 23468 56600 23480
rect 56652 23468 56658 23520
rect 57882 23468 57888 23520
rect 57940 23468 57946 23520
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 4614 23264 4620 23316
rect 4672 23304 4678 23316
rect 4709 23307 4767 23313
rect 4709 23304 4721 23307
rect 4672 23276 4721 23304
rect 4672 23264 4678 23276
rect 4709 23273 4721 23276
rect 4755 23273 4767 23307
rect 4709 23267 4767 23273
rect 6822 23264 6828 23316
rect 6880 23264 6886 23316
rect 7285 23307 7343 23313
rect 7285 23273 7297 23307
rect 7331 23304 7343 23307
rect 7374 23304 7380 23316
rect 7331 23276 7380 23304
rect 7331 23273 7343 23276
rect 7285 23267 7343 23273
rect 7374 23264 7380 23276
rect 7432 23264 7438 23316
rect 7926 23264 7932 23316
rect 7984 23264 7990 23316
rect 8110 23264 8116 23316
rect 8168 23304 8174 23316
rect 8205 23307 8263 23313
rect 8205 23304 8217 23307
rect 8168 23276 8217 23304
rect 8168 23264 8174 23276
rect 8205 23273 8217 23276
rect 8251 23273 8263 23307
rect 8205 23267 8263 23273
rect 11882 23264 11888 23316
rect 11940 23304 11946 23316
rect 12345 23307 12403 23313
rect 12345 23304 12357 23307
rect 11940 23276 12357 23304
rect 11940 23264 11946 23276
rect 12345 23273 12357 23276
rect 12391 23273 12403 23307
rect 12345 23267 12403 23273
rect 39209 23307 39267 23313
rect 39209 23273 39221 23307
rect 39255 23304 39267 23307
rect 39390 23304 39396 23316
rect 39255 23276 39396 23304
rect 39255 23273 39267 23276
rect 39209 23267 39267 23273
rect 39390 23264 39396 23276
rect 39448 23264 39454 23316
rect 40218 23304 40224 23316
rect 39592 23276 40224 23304
rect 3510 23196 3516 23248
rect 3568 23236 3574 23248
rect 3881 23239 3939 23245
rect 3881 23236 3893 23239
rect 3568 23208 3893 23236
rect 3568 23196 3574 23208
rect 3881 23205 3893 23208
rect 3927 23205 3939 23239
rect 3881 23199 3939 23205
rect 4706 23128 4712 23180
rect 4764 23128 4770 23180
rect 6641 23171 6699 23177
rect 6641 23137 6653 23171
rect 6687 23168 6699 23171
rect 6840 23168 6868 23264
rect 7944 23168 7972 23264
rect 6687 23140 6868 23168
rect 6932 23140 7972 23168
rect 37369 23171 37427 23177
rect 6687 23137 6699 23140
rect 6641 23131 6699 23137
rect 2593 23103 2651 23109
rect 2593 23100 2605 23103
rect 2332 23072 2605 23100
rect 934 22992 940 23044
rect 992 23032 998 23044
rect 1581 23035 1639 23041
rect 1581 23032 1593 23035
rect 992 23004 1593 23032
rect 992 22992 998 23004
rect 1581 23001 1593 23004
rect 1627 23001 1639 23035
rect 1581 22995 1639 23001
rect 1394 22924 1400 22976
rect 1452 22964 1458 22976
rect 2332 22964 2360 23072
rect 2593 23069 2605 23072
rect 2639 23100 2651 23103
rect 2869 23103 2927 23109
rect 2869 23100 2881 23103
rect 2639 23072 2881 23100
rect 2639 23069 2651 23072
rect 2593 23063 2651 23069
rect 2869 23069 2881 23072
rect 2915 23069 2927 23103
rect 2869 23063 2927 23069
rect 3789 23103 3847 23109
rect 3789 23069 3801 23103
rect 3835 23100 3847 23103
rect 3878 23100 3884 23112
rect 3835 23072 3884 23100
rect 3835 23069 3847 23072
rect 3789 23063 3847 23069
rect 3878 23060 3884 23072
rect 3936 23060 3942 23112
rect 3973 23103 4031 23109
rect 3973 23069 3985 23103
rect 4019 23100 4031 23103
rect 4617 23103 4675 23109
rect 4617 23100 4629 23103
rect 4019 23072 4629 23100
rect 4019 23069 4031 23072
rect 3973 23063 4031 23069
rect 4617 23069 4629 23072
rect 4663 23100 4675 23103
rect 4724 23100 4752 23128
rect 4663 23072 4752 23100
rect 4801 23103 4859 23109
rect 4663 23069 4675 23072
rect 4617 23063 4675 23069
rect 4801 23069 4813 23103
rect 4847 23069 4859 23103
rect 4801 23063 4859 23069
rect 4816 23032 4844 23063
rect 6546 23060 6552 23112
rect 6604 23100 6610 23112
rect 6932 23109 6960 23140
rect 37369 23137 37381 23171
rect 37415 23168 37427 23171
rect 37461 23171 37519 23177
rect 37461 23168 37473 23171
rect 37415 23140 37473 23168
rect 37415 23137 37427 23140
rect 37369 23131 37427 23137
rect 37461 23137 37473 23140
rect 37507 23168 37519 23171
rect 39592 23168 39620 23276
rect 40218 23264 40224 23276
rect 40276 23264 40282 23316
rect 42702 23264 42708 23316
rect 42760 23264 42766 23316
rect 47302 23264 47308 23316
rect 47360 23264 47366 23316
rect 47872 23276 48268 23304
rect 37507 23140 39620 23168
rect 37507 23137 37519 23140
rect 37461 23131 37519 23137
rect 6825 23103 6883 23109
rect 6825 23100 6837 23103
rect 6604 23072 6837 23100
rect 6604 23060 6610 23072
rect 6825 23069 6837 23072
rect 6871 23069 6883 23103
rect 6825 23063 6883 23069
rect 6917 23103 6975 23109
rect 6917 23069 6929 23103
rect 6963 23069 6975 23103
rect 6917 23063 6975 23069
rect 4724 23004 4844 23032
rect 6840 23032 6868 23063
rect 7006 23060 7012 23112
rect 7064 23100 7070 23112
rect 7193 23103 7251 23109
rect 7193 23100 7205 23103
rect 7064 23072 7205 23100
rect 7064 23060 7070 23072
rect 7193 23069 7205 23072
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 7377 23103 7435 23109
rect 7377 23069 7389 23103
rect 7423 23100 7435 23103
rect 7834 23100 7840 23112
rect 7423 23072 7840 23100
rect 7423 23069 7435 23072
rect 7377 23063 7435 23069
rect 7834 23060 7840 23072
rect 7892 23060 7898 23112
rect 8297 23103 8355 23109
rect 8297 23069 8309 23103
rect 8343 23100 8355 23103
rect 8386 23100 8392 23112
rect 8343 23072 8392 23100
rect 8343 23069 8355 23072
rect 8297 23063 8355 23069
rect 8386 23060 8392 23072
rect 8444 23100 8450 23112
rect 8573 23103 8631 23109
rect 8573 23100 8585 23103
rect 8444 23072 8585 23100
rect 8444 23060 8450 23072
rect 8573 23069 8585 23072
rect 8619 23069 8631 23103
rect 8573 23063 8631 23069
rect 9950 23060 9956 23112
rect 10008 23060 10014 23112
rect 10134 23060 10140 23112
rect 10192 23060 10198 23112
rect 39390 23060 39396 23112
rect 39448 23100 39454 23112
rect 39500 23109 39528 23140
rect 39485 23103 39543 23109
rect 39485 23100 39497 23103
rect 39448 23072 39497 23100
rect 39448 23060 39454 23072
rect 39485 23069 39497 23072
rect 39531 23069 39543 23103
rect 39485 23063 39543 23069
rect 39577 23103 39635 23109
rect 39577 23069 39589 23103
rect 39623 23100 39635 23103
rect 39853 23103 39911 23109
rect 39853 23100 39865 23103
rect 39623 23072 39865 23100
rect 39623 23069 39635 23072
rect 39577 23063 39635 23069
rect 39853 23069 39865 23072
rect 39899 23069 39911 23103
rect 39853 23063 39911 23069
rect 41230 23060 41236 23112
rect 41288 23100 41294 23112
rect 42720 23100 42748 23264
rect 46658 23236 46664 23248
rect 46400 23208 46664 23236
rect 41288 23072 42748 23100
rect 41288 23060 41294 23072
rect 44174 23060 44180 23112
rect 44232 23100 44238 23112
rect 45005 23103 45063 23109
rect 45005 23100 45017 23103
rect 44232 23072 45017 23100
rect 44232 23060 44238 23072
rect 45005 23069 45017 23072
rect 45051 23069 45063 23103
rect 46400 23086 46428 23208
rect 46658 23196 46664 23208
rect 46716 23236 46722 23248
rect 47320 23236 47348 23264
rect 46716 23208 47348 23236
rect 46716 23196 46722 23208
rect 46753 23171 46811 23177
rect 46753 23137 46765 23171
rect 46799 23168 46811 23171
rect 47872 23168 47900 23276
rect 48240 23248 48268 23276
rect 48590 23264 48596 23316
rect 48648 23264 48654 23316
rect 49970 23304 49976 23316
rect 48700 23276 49976 23304
rect 48038 23196 48044 23248
rect 48096 23196 48102 23248
rect 48222 23196 48228 23248
rect 48280 23236 48286 23248
rect 48700 23236 48728 23276
rect 49970 23264 49976 23276
rect 50028 23264 50034 23316
rect 52730 23264 52736 23316
rect 52788 23304 52794 23316
rect 52825 23307 52883 23313
rect 52825 23304 52837 23307
rect 52788 23276 52837 23304
rect 52788 23264 52794 23276
rect 52825 23273 52837 23276
rect 52871 23273 52883 23307
rect 52825 23267 52883 23273
rect 56502 23264 56508 23316
rect 56560 23264 56566 23316
rect 56597 23307 56655 23313
rect 56597 23273 56609 23307
rect 56643 23304 56655 23307
rect 56778 23304 56784 23316
rect 56643 23276 56784 23304
rect 56643 23273 56655 23276
rect 56597 23267 56655 23273
rect 56778 23264 56784 23276
rect 56836 23264 56842 23316
rect 58345 23307 58403 23313
rect 58345 23304 58357 23307
rect 57256 23276 58357 23304
rect 48280 23208 48728 23236
rect 48777 23239 48835 23245
rect 48280 23196 48286 23208
rect 46799 23140 46888 23168
rect 46799 23137 46811 23140
rect 46753 23131 46811 23137
rect 46860 23109 46888 23140
rect 47780 23140 47900 23168
rect 48056 23168 48084 23196
rect 48516 23177 48544 23208
rect 48777 23205 48789 23239
rect 48823 23205 48835 23239
rect 48777 23199 48835 23205
rect 48501 23171 48559 23177
rect 48056 23140 48268 23168
rect 47780 23109 47808 23140
rect 46845 23103 46903 23109
rect 45005 23063 45063 23069
rect 46845 23069 46857 23103
rect 46891 23069 46903 23103
rect 46845 23063 46903 23069
rect 47765 23103 47823 23109
rect 47765 23069 47777 23103
rect 47811 23069 47823 23103
rect 47765 23063 47823 23069
rect 47854 23060 47860 23112
rect 47912 23100 47918 23112
rect 48240 23109 48268 23140
rect 48501 23137 48513 23171
rect 48547 23137 48559 23171
rect 48501 23131 48559 23137
rect 48041 23103 48099 23109
rect 48041 23100 48053 23103
rect 47912 23072 48053 23100
rect 47912 23060 47918 23072
rect 48041 23069 48053 23072
rect 48087 23069 48099 23103
rect 48041 23063 48099 23069
rect 48225 23103 48283 23109
rect 48225 23069 48237 23103
rect 48271 23069 48283 23103
rect 48792 23100 48820 23199
rect 48958 23196 48964 23248
rect 49016 23196 49022 23248
rect 49602 23196 49608 23248
rect 49660 23236 49666 23248
rect 51166 23236 51172 23248
rect 49660 23208 51172 23236
rect 49660 23196 49666 23208
rect 51166 23196 51172 23208
rect 51224 23196 51230 23248
rect 52454 23236 52460 23248
rect 51276 23208 52460 23236
rect 49145 23171 49203 23177
rect 49145 23137 49157 23171
rect 49191 23168 49203 23171
rect 49237 23171 49295 23177
rect 49237 23168 49249 23171
rect 49191 23140 49249 23168
rect 49191 23137 49203 23140
rect 49145 23131 49203 23137
rect 49237 23137 49249 23140
rect 49283 23137 49295 23171
rect 49237 23131 49295 23137
rect 49881 23171 49939 23177
rect 49881 23137 49893 23171
rect 49927 23168 49939 23171
rect 50062 23168 50068 23180
rect 49927 23140 50068 23168
rect 49927 23137 49939 23140
rect 49881 23131 49939 23137
rect 50062 23128 50068 23140
rect 50120 23128 50126 23180
rect 48869 23103 48927 23109
rect 48869 23100 48881 23103
rect 48792 23072 48881 23100
rect 48225 23063 48283 23069
rect 48869 23069 48881 23072
rect 48915 23069 48927 23103
rect 48869 23063 48927 23069
rect 50157 23103 50215 23109
rect 50157 23069 50169 23103
rect 50203 23069 50215 23103
rect 50157 23063 50215 23069
rect 7653 23035 7711 23041
rect 7653 23032 7665 23035
rect 6840 23004 7665 23032
rect 4724 22976 4752 23004
rect 7653 23001 7665 23004
rect 7699 23001 7711 23035
rect 7653 22995 7711 23001
rect 37734 22992 37740 23044
rect 37792 22992 37798 23044
rect 39758 23032 39764 23044
rect 38962 23004 39764 23032
rect 39758 22992 39764 23004
rect 39816 22992 39822 23044
rect 40126 22992 40132 23044
rect 40184 22992 40190 23044
rect 41877 23035 41935 23041
rect 41877 23001 41889 23035
rect 41923 23001 41935 23035
rect 41877 22995 41935 23001
rect 1452 22936 2360 22964
rect 1452 22924 1458 22936
rect 3510 22924 3516 22976
rect 3568 22924 3574 22976
rect 4706 22924 4712 22976
rect 4764 22924 4770 22976
rect 6638 22924 6644 22976
rect 6696 22924 6702 22976
rect 10134 22924 10140 22976
rect 10192 22924 10198 22976
rect 12894 22924 12900 22976
rect 12952 22924 12958 22976
rect 41892 22964 41920 22995
rect 45278 22992 45284 23044
rect 45336 22992 45342 23044
rect 46934 22992 46940 23044
rect 46992 23032 46998 23044
rect 47581 23035 47639 23041
rect 47581 23032 47593 23035
rect 46992 23004 47593 23032
rect 46992 22992 46998 23004
rect 47581 23001 47593 23004
rect 47627 23001 47639 23035
rect 47581 22995 47639 23001
rect 49145 23035 49203 23041
rect 49145 23001 49157 23035
rect 49191 23032 49203 23035
rect 50172 23032 50200 23063
rect 50338 23060 50344 23112
rect 50396 23100 50402 23112
rect 50893 23103 50951 23109
rect 50893 23100 50905 23103
rect 50396 23072 50905 23100
rect 50396 23060 50402 23072
rect 50893 23069 50905 23072
rect 50939 23069 50951 23103
rect 50893 23063 50951 23069
rect 51169 23103 51227 23109
rect 51169 23069 51181 23103
rect 51215 23100 51227 23103
rect 51276 23100 51304 23208
rect 52454 23196 52460 23208
rect 52512 23236 52518 23248
rect 52512 23208 52776 23236
rect 52512 23196 52518 23208
rect 52549 23171 52607 23177
rect 52549 23168 52561 23171
rect 52104 23140 52561 23168
rect 51215 23072 51304 23100
rect 51215 23069 51227 23072
rect 51169 23063 51227 23069
rect 51350 23060 51356 23112
rect 51408 23060 51414 23112
rect 51537 23103 51595 23109
rect 51537 23069 51549 23103
rect 51583 23100 51595 23103
rect 51629 23103 51687 23109
rect 51629 23100 51641 23103
rect 51583 23072 51641 23100
rect 51583 23069 51595 23072
rect 51537 23063 51595 23069
rect 51629 23069 51641 23072
rect 51675 23069 51687 23103
rect 51629 23063 51687 23069
rect 51813 23103 51871 23109
rect 51813 23069 51825 23103
rect 51859 23069 51871 23103
rect 51813 23063 51871 23069
rect 49191 23004 50200 23032
rect 49191 23001 49203 23004
rect 49145 22995 49203 23001
rect 50522 22992 50528 23044
rect 50580 23032 50586 23044
rect 51552 23032 51580 23063
rect 50580 23004 51580 23032
rect 50580 22992 50586 23004
rect 42242 22964 42248 22976
rect 41892 22936 42248 22964
rect 42242 22924 42248 22936
rect 42300 22924 42306 22976
rect 47026 22924 47032 22976
rect 47084 22924 47090 22976
rect 47946 22924 47952 22976
rect 48004 22924 48010 22976
rect 50798 22924 50804 22976
rect 50856 22924 50862 22976
rect 51442 22924 51448 22976
rect 51500 22924 51506 22976
rect 51552 22964 51580 23004
rect 51718 22992 51724 23044
rect 51776 22992 51782 23044
rect 51828 23032 51856 23063
rect 51902 23060 51908 23112
rect 51960 23060 51966 23112
rect 52104 23109 52132 23140
rect 52549 23137 52561 23140
rect 52595 23137 52607 23171
rect 52549 23131 52607 23137
rect 52089 23103 52147 23109
rect 52089 23069 52101 23103
rect 52135 23069 52147 23103
rect 52089 23063 52147 23069
rect 52181 23103 52239 23109
rect 52181 23069 52193 23103
rect 52227 23069 52239 23103
rect 52181 23063 52239 23069
rect 51997 23035 52055 23041
rect 51997 23032 52009 23035
rect 51828 23004 52009 23032
rect 51997 23001 52009 23004
rect 52043 23001 52055 23035
rect 51997 22995 52055 23001
rect 52196 22964 52224 23063
rect 52362 23060 52368 23112
rect 52420 23060 52426 23112
rect 52454 23060 52460 23112
rect 52512 23060 52518 23112
rect 52748 23109 52776 23208
rect 55677 23171 55735 23177
rect 55677 23168 55689 23171
rect 55508 23140 55689 23168
rect 52641 23103 52699 23109
rect 52641 23102 52653 23103
rect 52564 23074 52653 23102
rect 51552 22936 52224 22964
rect 52270 22924 52276 22976
rect 52328 22924 52334 22976
rect 52564 22964 52592 23074
rect 52641 23069 52653 23074
rect 52687 23069 52699 23103
rect 52641 23063 52699 23069
rect 52733 23103 52791 23109
rect 52733 23069 52745 23103
rect 52779 23069 52791 23103
rect 52733 23063 52791 23069
rect 52917 23103 52975 23109
rect 52917 23069 52929 23103
rect 52963 23069 52975 23103
rect 52917 23063 52975 23069
rect 52932 23032 52960 23063
rect 53466 23060 53472 23112
rect 53524 23060 53530 23112
rect 53653 23103 53711 23109
rect 53653 23069 53665 23103
rect 53699 23100 53711 23103
rect 54478 23100 54484 23112
rect 53699 23072 54484 23100
rect 53699 23069 53711 23072
rect 53653 23063 53711 23069
rect 54478 23060 54484 23072
rect 54536 23060 54542 23112
rect 55306 23060 55312 23112
rect 55364 23060 55370 23112
rect 55508 23109 55536 23140
rect 55677 23137 55689 23140
rect 55723 23137 55735 23171
rect 55677 23131 55735 23137
rect 56413 23171 56471 23177
rect 56413 23137 56425 23171
rect 56459 23168 56471 23171
rect 56781 23171 56839 23177
rect 56781 23168 56793 23171
rect 56459 23140 56793 23168
rect 56459 23137 56471 23140
rect 56413 23131 56471 23137
rect 56781 23137 56793 23140
rect 56827 23137 56839 23171
rect 56781 23131 56839 23137
rect 55493 23103 55551 23109
rect 55493 23069 55505 23103
rect 55539 23069 55551 23103
rect 55493 23063 55551 23069
rect 55585 23103 55643 23109
rect 55585 23069 55597 23103
rect 55631 23069 55643 23103
rect 55585 23063 55643 23069
rect 55769 23103 55827 23109
rect 55769 23069 55781 23103
rect 55815 23069 55827 23103
rect 55769 23063 55827 23069
rect 56689 23103 56747 23109
rect 56689 23069 56701 23103
rect 56735 23100 56747 23103
rect 57256 23100 57284 23276
rect 57882 23236 57888 23248
rect 57532 23208 57888 23236
rect 57532 23112 57560 23208
rect 57882 23196 57888 23208
rect 57940 23196 57946 23248
rect 57793 23171 57851 23177
rect 57793 23137 57805 23171
rect 57839 23168 57851 23171
rect 58069 23171 58127 23177
rect 58069 23168 58081 23171
rect 57839 23140 58081 23168
rect 57839 23137 57851 23140
rect 57793 23131 57851 23137
rect 58069 23137 58081 23140
rect 58115 23137 58127 23171
rect 58069 23131 58127 23137
rect 56735 23072 57284 23100
rect 56735 23069 56747 23072
rect 56689 23063 56747 23069
rect 55401 23035 55459 23041
rect 55401 23032 55413 23035
rect 52932 23004 55413 23032
rect 55401 23001 55413 23004
rect 55447 23001 55459 23035
rect 55401 22995 55459 23001
rect 53561 22967 53619 22973
rect 53561 22964 53573 22967
rect 52564 22936 53573 22964
rect 53561 22933 53573 22936
rect 53607 22933 53619 22967
rect 53561 22927 53619 22933
rect 54386 22924 54392 22976
rect 54444 22964 54450 22976
rect 55600 22964 55628 23063
rect 55784 23032 55812 23063
rect 57330 23060 57336 23112
rect 57388 23060 57394 23112
rect 57514 23060 57520 23112
rect 57572 23060 57578 23112
rect 57606 23060 57612 23112
rect 57664 23060 57670 23112
rect 57974 23060 57980 23112
rect 58032 23060 58038 23112
rect 58176 23109 58204 23276
rect 58345 23273 58357 23276
rect 58391 23273 58403 23307
rect 58345 23267 58403 23273
rect 58161 23103 58219 23109
rect 58161 23069 58173 23103
rect 58207 23069 58219 23103
rect 58161 23063 58219 23069
rect 58250 23060 58256 23112
rect 58308 23060 58314 23112
rect 57793 23035 57851 23041
rect 57793 23032 57805 23035
rect 55784 23004 57805 23032
rect 57793 23001 57805 23004
rect 57839 23001 57851 23035
rect 57793 22995 57851 23001
rect 56042 22964 56048 22976
rect 54444 22936 56048 22964
rect 54444 22924 54450 22936
rect 56042 22924 56048 22936
rect 56100 22924 56106 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 1394 22720 1400 22772
rect 1452 22720 1458 22772
rect 3510 22720 3516 22772
rect 3568 22720 3574 22772
rect 3970 22720 3976 22772
rect 4028 22760 4034 22772
rect 4154 22760 4160 22772
rect 4028 22732 4160 22760
rect 4028 22720 4034 22732
rect 4154 22720 4160 22732
rect 4212 22720 4218 22772
rect 8018 22720 8024 22772
rect 8076 22720 8082 22772
rect 8386 22720 8392 22772
rect 8444 22760 8450 22772
rect 8665 22763 8723 22769
rect 8665 22760 8677 22763
rect 8444 22732 8677 22760
rect 8444 22720 8450 22732
rect 8665 22729 8677 22732
rect 8711 22729 8723 22763
rect 8665 22723 8723 22729
rect 9950 22720 9956 22772
rect 10008 22720 10014 22772
rect 11882 22720 11888 22772
rect 11940 22760 11946 22772
rect 11940 22732 26234 22760
rect 11940 22720 11946 22732
rect 2406 22652 2412 22704
rect 2464 22652 2470 22704
rect 3142 22584 3148 22636
rect 3200 22584 3206 22636
rect 3528 22624 3556 22720
rect 4172 22633 4200 22720
rect 3973 22627 4031 22633
rect 3973 22624 3985 22627
rect 3528 22596 3985 22624
rect 3973 22593 3985 22596
rect 4019 22593 4031 22627
rect 3973 22587 4031 22593
rect 4157 22627 4215 22633
rect 4157 22593 4169 22627
rect 4203 22593 4215 22627
rect 4157 22587 4215 22593
rect 4525 22627 4583 22633
rect 4525 22593 4537 22627
rect 4571 22593 4583 22627
rect 4525 22587 4583 22593
rect 2869 22559 2927 22565
rect 2869 22525 2881 22559
rect 2915 22556 2927 22559
rect 3326 22556 3332 22568
rect 2915 22528 3332 22556
rect 2915 22525 2927 22528
rect 2869 22519 2927 22525
rect 3326 22516 3332 22528
rect 3384 22516 3390 22568
rect 3881 22559 3939 22565
rect 3881 22525 3893 22559
rect 3927 22556 3939 22559
rect 4065 22559 4123 22565
rect 4065 22556 4077 22559
rect 3927 22528 4077 22556
rect 3927 22525 3939 22528
rect 3881 22519 3939 22525
rect 4065 22525 4077 22528
rect 4111 22525 4123 22559
rect 4065 22519 4123 22525
rect 4540 22488 4568 22587
rect 4706 22584 4712 22636
rect 4764 22584 4770 22636
rect 7374 22584 7380 22636
rect 7432 22624 7438 22636
rect 7929 22627 7987 22633
rect 7929 22624 7941 22627
rect 7432 22596 7941 22624
rect 7432 22584 7438 22596
rect 7929 22593 7941 22596
rect 7975 22593 7987 22627
rect 8036 22624 8064 22720
rect 8113 22627 8171 22633
rect 8113 22624 8125 22627
rect 8036 22596 8125 22624
rect 7929 22587 7987 22593
rect 8113 22593 8125 22596
rect 8159 22593 8171 22627
rect 8113 22587 8171 22593
rect 8205 22627 8263 22633
rect 8205 22593 8217 22627
rect 8251 22624 8263 22627
rect 8404 22624 8432 22720
rect 9306 22652 9312 22704
rect 9364 22652 9370 22704
rect 8251 22596 8432 22624
rect 9125 22627 9183 22633
rect 8251 22593 8263 22596
rect 8205 22587 8263 22593
rect 9125 22593 9137 22627
rect 9171 22624 9183 22627
rect 9214 22624 9220 22636
rect 9171 22596 9220 22624
rect 9171 22593 9183 22596
rect 9125 22587 9183 22593
rect 4724 22556 4752 22584
rect 5350 22556 5356 22568
rect 4724 22528 5356 22556
rect 5350 22516 5356 22528
rect 5408 22516 5414 22568
rect 7006 22516 7012 22568
rect 7064 22556 7070 22568
rect 8220 22556 8248 22587
rect 9214 22584 9220 22596
rect 9272 22584 9278 22636
rect 9674 22584 9680 22636
rect 9732 22624 9738 22636
rect 9769 22627 9827 22633
rect 9769 22624 9781 22627
rect 9732 22596 9781 22624
rect 9732 22584 9738 22596
rect 9769 22593 9781 22596
rect 9815 22593 9827 22627
rect 9769 22587 9827 22593
rect 9861 22627 9919 22633
rect 9861 22593 9873 22627
rect 9907 22624 9919 22627
rect 9968 22624 9996 22720
rect 12621 22695 12679 22701
rect 12621 22661 12633 22695
rect 12667 22692 12679 22695
rect 12897 22695 12955 22701
rect 12897 22692 12909 22695
rect 12667 22664 12909 22692
rect 12667 22661 12679 22664
rect 12621 22655 12679 22661
rect 12897 22661 12909 22664
rect 12943 22661 12955 22695
rect 12897 22655 12955 22661
rect 9907 22596 9996 22624
rect 9907 22593 9919 22596
rect 9861 22587 9919 22593
rect 7064 22528 8248 22556
rect 7064 22516 7070 22528
rect 4798 22488 4804 22500
rect 4540 22460 4804 22488
rect 4798 22448 4804 22460
rect 4856 22448 4862 22500
rect 8220 22488 8248 22528
rect 9493 22559 9551 22565
rect 9493 22525 9505 22559
rect 9539 22556 9551 22559
rect 9585 22559 9643 22565
rect 9585 22556 9597 22559
rect 9539 22528 9597 22556
rect 9539 22525 9551 22528
rect 9493 22519 9551 22525
rect 9585 22525 9597 22528
rect 9631 22525 9643 22559
rect 9784 22556 9812 22587
rect 10778 22584 10784 22636
rect 10836 22624 10842 22636
rect 11066 22627 11124 22633
rect 11066 22624 11078 22627
rect 10836 22596 11078 22624
rect 10836 22584 10842 22596
rect 11066 22593 11078 22596
rect 11112 22593 11124 22627
rect 11066 22587 11124 22593
rect 12434 22584 12440 22636
rect 12492 22584 12498 22636
rect 12710 22584 12716 22636
rect 12768 22584 12774 22636
rect 12802 22584 12808 22636
rect 12860 22584 12866 22636
rect 12986 22584 12992 22636
rect 13044 22584 13050 22636
rect 9950 22556 9956 22568
rect 9784 22528 9956 22556
rect 9585 22519 9643 22525
rect 9950 22516 9956 22528
rect 10008 22516 10014 22568
rect 11330 22516 11336 22568
rect 11388 22516 11394 22568
rect 26206 22488 26234 22732
rect 39390 22720 39396 22772
rect 39448 22720 39454 22772
rect 40126 22720 40132 22772
rect 40184 22760 40190 22772
rect 40313 22763 40371 22769
rect 40313 22760 40325 22763
rect 40184 22732 40325 22760
rect 40184 22720 40190 22732
rect 40313 22729 40325 22732
rect 40359 22729 40371 22763
rect 40313 22723 40371 22729
rect 40862 22720 40868 22772
rect 40920 22720 40926 22772
rect 43254 22720 43260 22772
rect 43312 22720 43318 22772
rect 43901 22763 43959 22769
rect 43901 22729 43913 22763
rect 43947 22760 43959 22763
rect 43990 22760 43996 22772
rect 43947 22732 43996 22760
rect 43947 22729 43959 22732
rect 43901 22723 43959 22729
rect 43990 22720 43996 22732
rect 44048 22720 44054 22772
rect 45278 22720 45284 22772
rect 45336 22760 45342 22772
rect 45557 22763 45615 22769
rect 45557 22760 45569 22763
rect 45336 22732 45569 22760
rect 45336 22720 45342 22732
rect 45557 22729 45569 22732
rect 45603 22729 45615 22763
rect 45557 22723 45615 22729
rect 46566 22720 46572 22772
rect 46624 22760 46630 22772
rect 46661 22763 46719 22769
rect 46661 22760 46673 22763
rect 46624 22732 46673 22760
rect 46624 22720 46630 22732
rect 46661 22729 46673 22732
rect 46707 22729 46719 22763
rect 46661 22723 46719 22729
rect 46934 22720 46940 22772
rect 46992 22720 46998 22772
rect 47026 22720 47032 22772
rect 47084 22720 47090 22772
rect 47397 22763 47455 22769
rect 47397 22729 47409 22763
rect 47443 22760 47455 22763
rect 47854 22760 47860 22772
rect 47443 22732 47860 22760
rect 47443 22729 47455 22732
rect 47397 22723 47455 22729
rect 47854 22720 47860 22732
rect 47912 22720 47918 22772
rect 47946 22720 47952 22772
rect 48004 22720 48010 22772
rect 48038 22720 48044 22772
rect 48096 22720 48102 22772
rect 49053 22763 49111 22769
rect 49053 22729 49065 22763
rect 49099 22760 49111 22763
rect 49786 22760 49792 22772
rect 49099 22732 49792 22760
rect 49099 22729 49111 22732
rect 49053 22723 49111 22729
rect 49786 22720 49792 22732
rect 49844 22720 49850 22772
rect 50798 22760 50804 22772
rect 50540 22732 50804 22760
rect 40497 22627 40555 22633
rect 40497 22593 40509 22627
rect 40543 22624 40555 22627
rect 40880 22624 40908 22720
rect 43272 22692 43300 22720
rect 46293 22695 46351 22701
rect 43272 22664 45876 22692
rect 40543 22596 40908 22624
rect 40543 22593 40555 22596
rect 40497 22587 40555 22593
rect 43162 22584 43168 22636
rect 43220 22624 43226 22636
rect 43349 22627 43407 22633
rect 43349 22624 43361 22627
rect 43220 22596 43361 22624
rect 43220 22584 43226 22596
rect 43349 22593 43361 22596
rect 43395 22624 43407 22627
rect 43993 22627 44051 22633
rect 43993 22624 44005 22627
rect 43395 22596 44005 22624
rect 43395 22593 43407 22596
rect 43349 22587 43407 22593
rect 43993 22593 44005 22596
rect 44039 22593 44051 22627
rect 43993 22587 44051 22593
rect 44177 22627 44235 22633
rect 44177 22593 44189 22627
rect 44223 22624 44235 22627
rect 44266 22624 44272 22636
rect 44223 22596 44272 22624
rect 44223 22593 44235 22596
rect 44177 22587 44235 22593
rect 44266 22584 44272 22596
rect 44324 22584 44330 22636
rect 39758 22516 39764 22568
rect 39816 22556 39822 22568
rect 41230 22556 41236 22568
rect 39816 22528 41236 22556
rect 39816 22516 39822 22528
rect 41230 22516 41236 22528
rect 41288 22516 41294 22568
rect 42978 22516 42984 22568
rect 43036 22516 43042 22568
rect 43438 22516 43444 22568
rect 43496 22556 43502 22568
rect 43625 22559 43683 22565
rect 43625 22556 43637 22559
rect 43496 22528 43637 22556
rect 43496 22516 43502 22528
rect 43625 22525 43637 22528
rect 43671 22525 43683 22559
rect 43625 22519 43683 22525
rect 44818 22488 44824 22500
rect 8220 22460 9812 22488
rect 26206 22460 44824 22488
rect 3234 22380 3240 22432
rect 3292 22380 3298 22432
rect 4614 22380 4620 22432
rect 4672 22380 4678 22432
rect 8018 22380 8024 22432
rect 8076 22380 8082 22432
rect 8297 22423 8355 22429
rect 8297 22389 8309 22423
rect 8343 22420 8355 22423
rect 8570 22420 8576 22432
rect 8343 22392 8576 22420
rect 8343 22389 8355 22392
rect 8297 22383 8355 22389
rect 8570 22380 8576 22392
rect 8628 22380 8634 22432
rect 9674 22380 9680 22432
rect 9732 22380 9738 22432
rect 9784 22420 9812 22460
rect 44818 22448 44824 22460
rect 44876 22448 44882 22500
rect 45848 22488 45876 22664
rect 46293 22661 46305 22695
rect 46339 22661 46351 22695
rect 46952 22692 46980 22720
rect 46293 22655 46351 22661
rect 46584 22664 46980 22692
rect 47044 22692 47072 22720
rect 48056 22692 48084 22720
rect 47044 22664 47624 22692
rect 46201 22627 46259 22633
rect 46201 22593 46213 22627
rect 46247 22624 46259 22627
rect 46308 22624 46336 22655
rect 46584 22633 46612 22664
rect 46247 22596 46336 22624
rect 46569 22627 46627 22633
rect 46247 22593 46259 22596
rect 46201 22587 46259 22593
rect 46569 22593 46581 22627
rect 46615 22593 46627 22627
rect 46569 22587 46627 22593
rect 46661 22627 46719 22633
rect 46661 22593 46673 22627
rect 46707 22624 46719 22627
rect 46750 22624 46756 22636
rect 46707 22596 46756 22624
rect 46707 22593 46719 22596
rect 46661 22587 46719 22593
rect 45922 22516 45928 22568
rect 45980 22556 45986 22568
rect 46293 22559 46351 22565
rect 46293 22556 46305 22559
rect 45980 22528 46305 22556
rect 45980 22516 45986 22528
rect 46293 22525 46305 22528
rect 46339 22525 46351 22559
rect 46293 22519 46351 22525
rect 46477 22559 46535 22565
rect 46477 22525 46489 22559
rect 46523 22556 46535 22559
rect 46676 22556 46704 22587
rect 46750 22584 46756 22596
rect 46808 22584 46814 22636
rect 46845 22627 46903 22633
rect 46845 22593 46857 22627
rect 46891 22624 46903 22627
rect 47044 22624 47072 22664
rect 47596 22633 47624 22664
rect 47780 22664 48084 22692
rect 48961 22695 49019 22701
rect 47780 22633 47808 22664
rect 48961 22661 48973 22695
rect 49007 22692 49019 22695
rect 49234 22692 49240 22704
rect 49007 22664 49240 22692
rect 49007 22661 49019 22664
rect 48961 22655 49019 22661
rect 49234 22652 49240 22664
rect 49292 22692 49298 22704
rect 50540 22701 50568 22732
rect 50798 22720 50804 22732
rect 50856 22720 50862 22772
rect 52822 22720 52828 22772
rect 52880 22760 52886 22772
rect 53098 22760 53104 22772
rect 52880 22732 53104 22760
rect 52880 22720 52886 22732
rect 53098 22720 53104 22732
rect 53156 22760 53162 22772
rect 53285 22763 53343 22769
rect 53285 22760 53297 22763
rect 53156 22732 53297 22760
rect 53156 22720 53162 22732
rect 53285 22729 53297 22732
rect 53331 22729 53343 22763
rect 53285 22723 53343 22729
rect 50525 22695 50583 22701
rect 49292 22664 49358 22692
rect 49292 22652 49298 22664
rect 50525 22661 50537 22695
rect 50571 22661 50583 22695
rect 53300 22692 53328 22723
rect 53466 22720 53472 22772
rect 53524 22760 53530 22772
rect 53561 22763 53619 22769
rect 53561 22760 53573 22763
rect 53524 22732 53573 22760
rect 53524 22720 53530 22732
rect 53561 22729 53573 22732
rect 53607 22729 53619 22763
rect 53561 22723 53619 22729
rect 55306 22720 55312 22772
rect 55364 22720 55370 22772
rect 57057 22763 57115 22769
rect 57057 22729 57069 22763
rect 57103 22760 57115 22763
rect 57330 22760 57336 22772
rect 57103 22732 57336 22760
rect 57103 22729 57115 22732
rect 57057 22723 57115 22729
rect 57330 22720 57336 22732
rect 57388 22720 57394 22772
rect 57422 22720 57428 22772
rect 57480 22720 57486 22772
rect 57514 22720 57520 22772
rect 57572 22720 57578 22772
rect 58069 22763 58127 22769
rect 58069 22729 58081 22763
rect 58115 22760 58127 22763
rect 58158 22760 58164 22772
rect 58115 22732 58164 22760
rect 58115 22729 58127 22732
rect 58069 22723 58127 22729
rect 58158 22720 58164 22732
rect 58216 22720 58222 22772
rect 58250 22720 58256 22772
rect 58308 22760 58314 22772
rect 58345 22763 58403 22769
rect 58345 22760 58357 22763
rect 58308 22732 58357 22760
rect 58308 22720 58314 22732
rect 58345 22729 58357 22732
rect 58391 22729 58403 22763
rect 58345 22723 58403 22729
rect 58894 22720 58900 22772
rect 58952 22720 58958 22772
rect 54941 22695 54999 22701
rect 54941 22692 54953 22695
rect 53300 22664 54953 22692
rect 50525 22655 50583 22661
rect 47121 22627 47179 22633
rect 47121 22624 47133 22627
rect 46891 22596 47133 22624
rect 46891 22593 46903 22596
rect 46845 22587 46903 22593
rect 47121 22593 47133 22596
rect 47167 22624 47179 22627
rect 47213 22627 47271 22633
rect 47213 22624 47225 22627
rect 47167 22596 47225 22624
rect 47167 22593 47179 22596
rect 47121 22587 47179 22593
rect 47213 22593 47225 22596
rect 47259 22593 47271 22627
rect 47213 22587 47271 22593
rect 47397 22627 47455 22633
rect 47397 22593 47409 22627
rect 47443 22593 47455 22627
rect 47397 22587 47455 22593
rect 47581 22627 47639 22633
rect 47581 22593 47593 22627
rect 47627 22593 47639 22627
rect 47581 22587 47639 22593
rect 47765 22627 47823 22633
rect 47765 22593 47777 22627
rect 47811 22593 47823 22627
rect 47765 22587 47823 22593
rect 47857 22627 47915 22633
rect 47857 22593 47869 22627
rect 47903 22593 47915 22627
rect 47857 22587 47915 22593
rect 46523 22528 46704 22556
rect 47412 22556 47440 22587
rect 47780 22556 47808 22587
rect 47412 22528 47808 22556
rect 46523 22525 46535 22528
rect 46477 22519 46535 22525
rect 47029 22491 47087 22497
rect 47029 22488 47041 22491
rect 45848 22460 47041 22488
rect 47029 22457 47041 22460
rect 47075 22457 47087 22491
rect 47029 22451 47087 22457
rect 10962 22420 10968 22432
rect 9784 22392 10968 22420
rect 10962 22380 10968 22392
rect 11020 22380 11026 22432
rect 11882 22380 11888 22432
rect 11940 22380 11946 22432
rect 12434 22380 12440 22432
rect 12492 22380 12498 22432
rect 42426 22380 42432 22432
rect 42484 22380 42490 22432
rect 43438 22380 43444 22432
rect 43496 22380 43502 22432
rect 43806 22380 43812 22432
rect 43864 22420 43870 22432
rect 43993 22423 44051 22429
rect 43993 22420 44005 22423
rect 43864 22392 44005 22420
rect 43864 22380 43870 22392
rect 43993 22389 44005 22392
rect 44039 22389 44051 22423
rect 47044 22420 47072 22451
rect 47210 22448 47216 22500
rect 47268 22488 47274 22500
rect 47765 22491 47823 22497
rect 47765 22488 47777 22491
rect 47268 22460 47777 22488
rect 47268 22448 47274 22460
rect 47765 22457 47777 22460
rect 47811 22488 47823 22491
rect 47872 22488 47900 22587
rect 48038 22584 48044 22636
rect 48096 22584 48102 22636
rect 53484 22633 53512 22664
rect 54941 22661 54953 22664
rect 54987 22692 54999 22695
rect 56781 22695 56839 22701
rect 56781 22692 56793 22695
rect 54987 22664 56793 22692
rect 54987 22661 54999 22664
rect 54941 22655 54999 22661
rect 53469 22627 53527 22633
rect 53469 22593 53481 22627
rect 53515 22624 53527 22627
rect 53653 22627 53711 22633
rect 53515 22596 53549 22624
rect 53515 22593 53527 22596
rect 53469 22587 53527 22593
rect 53653 22593 53665 22627
rect 53699 22624 53711 22627
rect 54754 22624 54760 22636
rect 53699 22596 54760 22624
rect 53699 22593 53711 22596
rect 53653 22587 53711 22593
rect 54754 22584 54760 22596
rect 54812 22584 54818 22636
rect 55140 22633 55168 22664
rect 56781 22661 56793 22664
rect 56827 22692 56839 22695
rect 57532 22692 57560 22720
rect 58912 22692 58940 22720
rect 56827 22664 57100 22692
rect 56827 22661 56839 22664
rect 56781 22655 56839 22661
rect 55125 22627 55183 22633
rect 55125 22593 55137 22627
rect 55171 22624 55183 22627
rect 55171 22596 55205 22624
rect 55171 22593 55183 22596
rect 55125 22587 55183 22593
rect 55306 22584 55312 22636
rect 55364 22584 55370 22636
rect 56965 22627 57023 22633
rect 56965 22593 56977 22627
rect 57011 22593 57023 22627
rect 56965 22587 57023 22593
rect 50798 22516 50804 22568
rect 50856 22516 50862 22568
rect 47811 22460 47900 22488
rect 47811 22457 47823 22460
rect 47765 22451 47823 22457
rect 56980 22432 57008 22587
rect 57072 22556 57100 22664
rect 57164 22664 57560 22692
rect 58544 22664 58940 22692
rect 57164 22633 57192 22664
rect 57149 22627 57207 22633
rect 57149 22593 57161 22627
rect 57195 22593 57207 22627
rect 57149 22587 57207 22593
rect 57241 22627 57299 22633
rect 57241 22593 57253 22627
rect 57287 22593 57299 22627
rect 57241 22587 57299 22593
rect 57256 22556 57284 22587
rect 57422 22584 57428 22636
rect 57480 22584 57486 22636
rect 58544 22633 58572 22664
rect 58253 22627 58311 22633
rect 58253 22593 58265 22627
rect 58299 22593 58311 22627
rect 58253 22587 58311 22593
rect 58529 22627 58587 22633
rect 58529 22593 58541 22627
rect 58575 22593 58587 22627
rect 58529 22587 58587 22593
rect 57072 22528 57284 22556
rect 58268 22556 58296 22587
rect 58802 22584 58808 22636
rect 58860 22584 58866 22636
rect 58820 22556 58848 22584
rect 58268 22528 58848 22556
rect 48866 22420 48872 22432
rect 47044 22392 48872 22420
rect 43993 22383 44051 22389
rect 48866 22380 48872 22392
rect 48924 22380 48930 22432
rect 52454 22380 52460 22432
rect 52512 22420 52518 22432
rect 53190 22420 53196 22432
rect 52512 22392 53196 22420
rect 52512 22380 52518 22392
rect 53190 22380 53196 22392
rect 53248 22420 53254 22432
rect 56686 22420 56692 22432
rect 53248 22392 56692 22420
rect 53248 22380 53254 22392
rect 56686 22380 56692 22392
rect 56744 22420 56750 22432
rect 56962 22420 56968 22432
rect 56744 22392 56968 22420
rect 56744 22380 56750 22392
rect 56962 22380 56968 22392
rect 57020 22380 57026 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 3234 22176 3240 22228
rect 3292 22176 3298 22228
rect 3326 22176 3332 22228
rect 3384 22176 3390 22228
rect 4798 22176 4804 22228
rect 4856 22216 4862 22228
rect 5537 22219 5595 22225
rect 5537 22216 5549 22219
rect 4856 22188 5549 22216
rect 4856 22176 4862 22188
rect 5537 22185 5549 22188
rect 5583 22185 5595 22219
rect 5537 22179 5595 22185
rect 7374 22176 7380 22228
rect 7432 22176 7438 22228
rect 8570 22176 8576 22228
rect 8628 22216 8634 22228
rect 8628 22188 8800 22216
rect 8628 22176 8634 22188
rect 2317 22151 2375 22157
rect 2317 22117 2329 22151
rect 2363 22148 2375 22151
rect 2866 22148 2872 22160
rect 2363 22120 2872 22148
rect 2363 22117 2375 22120
rect 2317 22111 2375 22117
rect 2866 22108 2872 22120
rect 2924 22108 2930 22160
rect 2501 22083 2559 22089
rect 2501 22049 2513 22083
rect 2547 22080 2559 22083
rect 3252 22080 3280 22176
rect 4062 22148 4068 22160
rect 2547 22052 3280 22080
rect 3436 22120 4068 22148
rect 2547 22049 2559 22052
rect 2501 22043 2559 22049
rect 3436 22021 3464 22120
rect 4062 22108 4068 22120
rect 4120 22108 4126 22160
rect 5718 22108 5724 22160
rect 5776 22108 5782 22160
rect 5905 22151 5963 22157
rect 5905 22117 5917 22151
rect 5951 22117 5963 22151
rect 5905 22111 5963 22117
rect 5920 22080 5948 22111
rect 3620 22052 4292 22080
rect 3620 22021 3648 22052
rect 2225 22015 2283 22021
rect 2225 21981 2237 22015
rect 2271 21981 2283 22015
rect 2685 22015 2743 22021
rect 2685 22012 2697 22015
rect 2225 21975 2283 21981
rect 2516 21984 2697 22012
rect 2240 21876 2268 21975
rect 2516 21953 2544 21984
rect 2685 21981 2697 21984
rect 2731 21981 2743 22015
rect 2685 21975 2743 21981
rect 3421 22015 3479 22021
rect 3421 21981 3433 22015
rect 3467 21981 3479 22015
rect 3421 21975 3479 21981
rect 3605 22015 3663 22021
rect 3605 21981 3617 22015
rect 3651 21981 3663 22015
rect 3605 21975 3663 21981
rect 3786 21972 3792 22024
rect 3844 22012 3850 22024
rect 3881 22015 3939 22021
rect 3881 22012 3893 22015
rect 3844 21984 3893 22012
rect 3844 21972 3850 21984
rect 3881 21981 3893 21984
rect 3927 21981 3939 22015
rect 3881 21975 3939 21981
rect 3973 22015 4031 22021
rect 3973 21981 3985 22015
rect 4019 22012 4031 22015
rect 4157 22015 4215 22021
rect 4157 22012 4169 22015
rect 4019 21984 4169 22012
rect 4019 21981 4031 21984
rect 3973 21975 4031 21981
rect 4157 21981 4169 21984
rect 4203 21981 4215 22015
rect 4157 21975 4215 21981
rect 2501 21947 2559 21953
rect 2501 21913 2513 21947
rect 2547 21913 2559 21947
rect 2501 21907 2559 21913
rect 3421 21879 3479 21885
rect 3421 21876 3433 21879
rect 2240 21848 3433 21876
rect 3421 21845 3433 21848
rect 3467 21845 3479 21879
rect 4264 21876 4292 22052
rect 5736 22052 5948 22080
rect 5350 21972 5356 22024
rect 5408 21972 5414 22024
rect 5626 21972 5632 22024
rect 5684 22012 5690 22024
rect 5736 22012 5764 22052
rect 5684 21984 5764 22012
rect 5813 22015 5871 22021
rect 5684 21972 5690 21984
rect 5813 21981 5825 22015
rect 5859 21981 5871 22015
rect 5813 21975 5871 21981
rect 4430 21953 4436 21956
rect 4424 21907 4436 21953
rect 4430 21904 4436 21907
rect 4488 21904 4494 21956
rect 5368 21944 5396 21972
rect 5828 21944 5856 21975
rect 5994 21972 6000 22024
rect 6052 22012 6058 22024
rect 7285 22015 7343 22021
rect 7285 22012 7297 22015
rect 6052 21984 7297 22012
rect 6052 21972 6058 21984
rect 7285 21981 7297 21984
rect 7331 21981 7343 22015
rect 7285 21975 7343 21981
rect 5368 21916 5856 21944
rect 6638 21904 6644 21956
rect 6696 21944 6702 21956
rect 7018 21947 7076 21953
rect 7018 21944 7030 21947
rect 6696 21916 7030 21944
rect 6696 21904 6702 21916
rect 7018 21913 7030 21916
rect 7064 21913 7076 21947
rect 7392 21944 7420 22176
rect 8772 22089 8800 22188
rect 9214 22176 9220 22228
rect 9272 22216 9278 22228
rect 9585 22219 9643 22225
rect 9585 22216 9597 22219
rect 9272 22188 9597 22216
rect 9272 22176 9278 22188
rect 9585 22185 9597 22188
rect 9631 22185 9643 22219
rect 9585 22179 9643 22185
rect 9950 22176 9956 22228
rect 10008 22216 10014 22228
rect 11701 22219 11759 22225
rect 11701 22216 11713 22219
rect 10008 22188 11713 22216
rect 10008 22176 10014 22188
rect 11701 22185 11713 22188
rect 11747 22216 11759 22219
rect 11882 22216 11888 22228
rect 11747 22188 11888 22216
rect 11747 22185 11759 22188
rect 11701 22179 11759 22185
rect 11882 22176 11888 22188
rect 11940 22176 11946 22228
rect 41220 22219 41278 22225
rect 41220 22185 41232 22219
rect 41266 22216 41278 22219
rect 42426 22216 42432 22228
rect 41266 22188 42432 22216
rect 41266 22185 41278 22188
rect 41220 22179 41278 22185
rect 42426 22176 42432 22188
rect 42484 22176 42490 22228
rect 42702 22176 42708 22228
rect 42760 22216 42766 22228
rect 43257 22219 43315 22225
rect 43257 22216 43269 22219
rect 42760 22188 43269 22216
rect 42760 22176 42766 22188
rect 43257 22185 43269 22188
rect 43303 22185 43315 22219
rect 43257 22179 43315 22185
rect 54754 22176 54760 22228
rect 54812 22176 54818 22228
rect 55306 22176 55312 22228
rect 55364 22216 55370 22228
rect 55401 22219 55459 22225
rect 55401 22216 55413 22219
rect 55364 22188 55413 22216
rect 55364 22176 55370 22188
rect 55401 22185 55413 22188
rect 55447 22185 55459 22219
rect 55401 22179 55459 22185
rect 57422 22176 57428 22228
rect 57480 22216 57486 22228
rect 57517 22219 57575 22225
rect 57517 22216 57529 22219
rect 57480 22188 57529 22216
rect 57480 22176 57486 22188
rect 57517 22185 57529 22188
rect 57563 22185 57575 22219
rect 57517 22179 57575 22185
rect 10412 22151 10470 22157
rect 10412 22117 10424 22151
rect 10458 22148 10470 22151
rect 10778 22148 10784 22160
rect 10458 22120 10784 22148
rect 10458 22117 10470 22120
rect 10412 22111 10470 22117
rect 10778 22108 10784 22120
rect 10836 22108 10842 22160
rect 10962 22108 10968 22160
rect 11020 22148 11026 22160
rect 54294 22148 54300 22160
rect 11020 22120 12112 22148
rect 11020 22108 11026 22120
rect 8757 22083 8815 22089
rect 8757 22049 8769 22083
rect 8803 22049 8815 22083
rect 8757 22043 8815 22049
rect 11514 22040 11520 22092
rect 11572 22040 11578 22092
rect 12084 22089 12112 22120
rect 54036 22120 54300 22148
rect 12069 22083 12127 22089
rect 12069 22049 12081 22083
rect 12115 22080 12127 22083
rect 40957 22083 41015 22089
rect 12115 22052 12296 22080
rect 12115 22049 12127 22052
rect 12069 22043 12127 22049
rect 10134 21972 10140 22024
rect 10192 21972 10198 22024
rect 10229 22015 10287 22021
rect 10229 21981 10241 22015
rect 10275 22012 10287 22015
rect 10318 22012 10324 22024
rect 10275 21984 10324 22012
rect 10275 21981 10287 21984
rect 10229 21975 10287 21981
rect 10318 21972 10324 21984
rect 10376 21972 10382 22024
rect 12268 22021 12296 22052
rect 40957 22049 40969 22083
rect 41003 22080 41015 22083
rect 41322 22080 41328 22092
rect 41003 22052 41328 22080
rect 41003 22049 41015 22052
rect 40957 22043 41015 22049
rect 41322 22040 41328 22052
rect 41380 22080 41386 22092
rect 44174 22080 44180 22092
rect 41380 22052 44180 22080
rect 41380 22040 41386 22052
rect 44174 22040 44180 22052
rect 44232 22040 44238 22092
rect 47397 22083 47455 22089
rect 47397 22049 47409 22083
rect 47443 22080 47455 22083
rect 47946 22080 47952 22092
rect 47443 22052 47952 22080
rect 47443 22049 47455 22052
rect 47397 22043 47455 22049
rect 47946 22040 47952 22052
rect 48004 22040 48010 22092
rect 48130 22040 48136 22092
rect 48188 22080 48194 22092
rect 49605 22083 49663 22089
rect 49605 22080 49617 22083
rect 48188 22052 49617 22080
rect 48188 22040 48194 22052
rect 11793 22015 11851 22021
rect 11793 21981 11805 22015
rect 11839 21981 11851 22015
rect 11793 21975 11851 21981
rect 12253 22015 12311 22021
rect 12253 21981 12265 22015
rect 12299 21981 12311 22015
rect 12253 21975 12311 21981
rect 12345 22015 12403 22021
rect 12345 21981 12357 22015
rect 12391 22012 12403 22015
rect 12529 22015 12587 22021
rect 12529 22012 12541 22015
rect 12391 21984 12541 22012
rect 12391 21981 12403 21984
rect 12345 21975 12403 21981
rect 12529 21981 12541 21984
rect 12575 21981 12587 22015
rect 42610 22012 42616 22024
rect 42366 21984 42616 22012
rect 12529 21975 12587 21981
rect 7018 21907 7076 21913
rect 7300 21916 7420 21944
rect 7300 21876 7328 21916
rect 8202 21904 8208 21956
rect 8260 21944 8266 21956
rect 8490 21947 8548 21953
rect 8490 21944 8502 21947
rect 8260 21916 8502 21944
rect 8260 21904 8266 21916
rect 8490 21913 8502 21916
rect 8536 21913 8548 21947
rect 8490 21907 8548 21913
rect 10413 21947 10471 21953
rect 10413 21913 10425 21947
rect 10459 21944 10471 21947
rect 10594 21944 10600 21956
rect 10459 21916 10600 21944
rect 10459 21913 10471 21916
rect 10413 21907 10471 21913
rect 10594 21904 10600 21916
rect 10652 21904 10658 21956
rect 4264 21848 7328 21876
rect 3421 21839 3479 21845
rect 9950 21836 9956 21888
rect 10008 21876 10014 21888
rect 11517 21879 11575 21885
rect 11517 21876 11529 21879
rect 10008 21848 11529 21876
rect 10008 21836 10014 21848
rect 11517 21845 11529 21848
rect 11563 21845 11575 21879
rect 11808 21876 11836 21975
rect 42610 21972 42616 21984
rect 42668 21972 42674 22024
rect 42797 22015 42855 22021
rect 42797 22012 42809 22015
rect 42720 21984 42809 22012
rect 12434 21904 12440 21956
rect 12492 21944 12498 21956
rect 12774 21947 12832 21953
rect 12774 21944 12786 21947
rect 12492 21916 12786 21944
rect 12492 21904 12498 21916
rect 12774 21913 12786 21916
rect 12820 21913 12832 21947
rect 12774 21907 12832 21913
rect 13078 21876 13084 21888
rect 11808 21848 13084 21876
rect 11517 21839 11575 21845
rect 13078 21836 13084 21848
rect 13136 21876 13142 21888
rect 42720 21885 42748 21984
rect 42797 21981 42809 21984
rect 42843 21981 42855 22015
rect 42797 21975 42855 21981
rect 42886 21972 42892 22024
rect 42944 22012 42950 22024
rect 44085 22015 44143 22021
rect 44085 22012 44097 22015
rect 42944 21984 44097 22012
rect 42944 21972 42950 21984
rect 44085 21981 44097 21984
rect 44131 21981 44143 22015
rect 44085 21975 44143 21981
rect 44266 21972 44272 22024
rect 44324 21972 44330 22024
rect 44453 22015 44511 22021
rect 44453 21981 44465 22015
rect 44499 21981 44511 22015
rect 44453 21975 44511 21981
rect 43162 21944 43168 21956
rect 42996 21916 43168 21944
rect 42996 21885 43024 21916
rect 43162 21904 43168 21916
rect 43220 21944 43226 21956
rect 44468 21944 44496 21975
rect 45646 21972 45652 22024
rect 45704 21972 45710 22024
rect 45741 22015 45799 22021
rect 45741 21981 45753 22015
rect 45787 21981 45799 22015
rect 45741 21975 45799 21981
rect 43220 21916 44496 21944
rect 43220 21904 43226 21916
rect 44542 21904 44548 21956
rect 44600 21944 44606 21956
rect 45756 21944 45784 21975
rect 47118 21972 47124 22024
rect 47176 21972 47182 22024
rect 48332 22021 48360 22052
rect 49605 22049 49617 22052
rect 49651 22080 49663 22083
rect 50154 22080 50160 22092
rect 49651 22052 50160 22080
rect 49651 22049 49663 22052
rect 49605 22043 49663 22049
rect 50154 22040 50160 22052
rect 50212 22080 50218 22092
rect 52549 22083 52607 22089
rect 50212 22052 51074 22080
rect 50212 22040 50218 22052
rect 48317 22015 48375 22021
rect 48317 21981 48329 22015
rect 48363 21981 48375 22015
rect 48317 21975 48375 21981
rect 49326 21972 49332 22024
rect 49384 21972 49390 22024
rect 44600 21916 45784 21944
rect 48593 21947 48651 21953
rect 44600 21904 44606 21916
rect 48593 21913 48605 21947
rect 48639 21944 48651 21947
rect 48682 21944 48688 21956
rect 48639 21916 48688 21944
rect 48639 21913 48651 21916
rect 48593 21907 48651 21913
rect 48682 21904 48688 21916
rect 48740 21944 48746 21956
rect 49142 21944 49148 21956
rect 48740 21916 49148 21944
rect 48740 21904 48746 21916
rect 49142 21904 49148 21916
rect 49200 21904 49206 21956
rect 13909 21879 13967 21885
rect 13909 21876 13921 21879
rect 13136 21848 13921 21876
rect 13136 21836 13142 21848
rect 13909 21845 13921 21848
rect 13955 21845 13967 21879
rect 13909 21839 13967 21845
rect 42705 21879 42763 21885
rect 42705 21845 42717 21879
rect 42751 21845 42763 21879
rect 42705 21839 42763 21845
rect 42981 21879 43039 21885
rect 42981 21845 42993 21879
rect 43027 21845 43039 21879
rect 42981 21839 43039 21845
rect 43530 21836 43536 21888
rect 43588 21836 43594 21888
rect 43990 21836 43996 21888
rect 44048 21876 44054 21888
rect 44269 21879 44327 21885
rect 44269 21876 44281 21879
rect 44048 21848 44281 21876
rect 44048 21836 44054 21848
rect 44269 21845 44281 21848
rect 44315 21845 44327 21879
rect 44269 21839 44327 21845
rect 44726 21836 44732 21888
rect 44784 21876 44790 21888
rect 45005 21879 45063 21885
rect 45005 21876 45017 21879
rect 44784 21848 45017 21876
rect 44784 21836 44790 21848
rect 45005 21845 45017 21848
rect 45051 21845 45063 21879
rect 45005 21839 45063 21845
rect 46198 21836 46204 21888
rect 46256 21876 46262 21888
rect 46385 21879 46443 21885
rect 46385 21876 46397 21879
rect 46256 21848 46397 21876
rect 46256 21836 46262 21848
rect 46385 21845 46397 21848
rect 46431 21845 46443 21879
rect 46385 21839 46443 21845
rect 49234 21836 49240 21888
rect 49292 21836 49298 21888
rect 51046 21876 51074 22052
rect 52549 22049 52561 22083
rect 52595 22080 52607 22083
rect 53285 22083 53343 22089
rect 53285 22080 53297 22083
rect 52595 22052 53297 22080
rect 52595 22049 52607 22052
rect 52549 22043 52607 22049
rect 53285 22049 53297 22052
rect 53331 22049 53343 22083
rect 53285 22043 53343 22049
rect 54036 22024 54064 22120
rect 54294 22108 54300 22120
rect 54352 22148 54358 22160
rect 54352 22120 54616 22148
rect 54352 22108 54358 22120
rect 54478 22080 54484 22092
rect 54220 22052 54484 22080
rect 51166 21972 51172 22024
rect 51224 22012 51230 22024
rect 51721 22015 51779 22021
rect 51721 22012 51733 22015
rect 51224 21984 51733 22012
rect 51224 21972 51230 21984
rect 51721 21981 51733 21984
rect 51767 21981 51779 22015
rect 51721 21975 51779 21981
rect 51997 22015 52055 22021
rect 51997 21981 52009 22015
rect 52043 22012 52055 22015
rect 52454 22012 52460 22024
rect 52043 21984 52460 22012
rect 52043 21981 52055 21984
rect 51997 21975 52055 21981
rect 52454 21972 52460 21984
rect 52512 21972 52518 22024
rect 52641 22015 52699 22021
rect 52641 21981 52653 22015
rect 52687 22012 52699 22015
rect 53558 22012 53564 22024
rect 52687 21984 53564 22012
rect 52687 21981 52699 21984
rect 52641 21975 52699 21981
rect 53558 21972 53564 21984
rect 53616 21972 53622 22024
rect 54018 21972 54024 22024
rect 54076 21972 54082 22024
rect 54110 21972 54116 22024
rect 54168 21972 54174 22024
rect 51445 21947 51503 21953
rect 51445 21913 51457 21947
rect 51491 21944 51503 21947
rect 52178 21944 52184 21956
rect 51491 21916 52184 21944
rect 51491 21913 51503 21916
rect 51445 21907 51503 21913
rect 52178 21904 52184 21916
rect 52236 21944 52242 21956
rect 54220 21944 54248 22052
rect 54478 22040 54484 22052
rect 54536 22040 54542 22092
rect 54588 22021 54616 22120
rect 55122 22108 55128 22160
rect 55180 22148 55186 22160
rect 55493 22151 55551 22157
rect 55493 22148 55505 22151
rect 55180 22120 55505 22148
rect 55180 22108 55186 22120
rect 55493 22117 55505 22120
rect 55539 22148 55551 22151
rect 57606 22148 57612 22160
rect 55539 22120 57612 22148
rect 55539 22117 55551 22120
rect 55493 22111 55551 22117
rect 57606 22108 57612 22120
rect 57664 22108 57670 22160
rect 55033 22083 55091 22089
rect 55033 22080 55045 22083
rect 54864 22052 55045 22080
rect 54864 22021 54892 22052
rect 55033 22049 55045 22052
rect 55079 22049 55091 22083
rect 55033 22043 55091 22049
rect 55309 22083 55367 22089
rect 55309 22049 55321 22083
rect 55355 22080 55367 22083
rect 57057 22083 57115 22089
rect 57057 22080 57069 22083
rect 55355 22052 57069 22080
rect 55355 22049 55367 22052
rect 55309 22043 55367 22049
rect 57057 22049 57069 22052
rect 57103 22049 57115 22083
rect 57057 22043 57115 22049
rect 57422 22040 57428 22092
rect 57480 22040 57486 22092
rect 57716 22052 58020 22080
rect 54573 22015 54631 22021
rect 54573 21981 54585 22015
rect 54619 21981 54631 22015
rect 54573 21975 54631 21981
rect 54665 22015 54723 22021
rect 54665 21981 54677 22015
rect 54711 21981 54723 22015
rect 54665 21975 54723 21981
rect 54849 22015 54907 22021
rect 54849 21981 54861 22015
rect 54895 21981 54907 22015
rect 54849 21975 54907 21981
rect 52236 21916 54248 21944
rect 54297 21947 54355 21953
rect 52236 21904 52242 21916
rect 54297 21913 54309 21947
rect 54343 21913 54355 21947
rect 54297 21907 54355 21913
rect 52362 21876 52368 21888
rect 51046 21848 52368 21876
rect 52362 21836 52368 21848
rect 52420 21836 52426 21888
rect 52730 21836 52736 21888
rect 52788 21836 52794 21888
rect 53926 21836 53932 21888
rect 53984 21876 53990 21888
rect 54202 21876 54208 21888
rect 53984 21848 54208 21876
rect 53984 21836 53990 21848
rect 54202 21836 54208 21848
rect 54260 21876 54266 21888
rect 54312 21876 54340 21907
rect 54478 21904 54484 21956
rect 54536 21904 54542 21956
rect 54260 21848 54340 21876
rect 54573 21879 54631 21885
rect 54260 21836 54266 21848
rect 54573 21845 54585 21879
rect 54619 21876 54631 21879
rect 54680 21876 54708 21975
rect 54938 21972 54944 22024
rect 54996 21972 55002 22024
rect 55125 22015 55183 22021
rect 55125 21981 55137 22015
rect 55171 22012 55183 22015
rect 55585 22015 55643 22021
rect 55171 21984 55260 22012
rect 55171 21981 55183 21984
rect 55125 21975 55183 21981
rect 54619 21848 54708 21876
rect 54956 21876 54984 21972
rect 55232 21956 55260 21984
rect 55585 21981 55597 22015
rect 55631 21981 55643 22015
rect 55585 21975 55643 21981
rect 55214 21904 55220 21956
rect 55272 21904 55278 21956
rect 55600 21944 55628 21975
rect 55950 21972 55956 22024
rect 56008 21972 56014 22024
rect 56689 22015 56747 22021
rect 56689 21981 56701 22015
rect 56735 21981 56747 22015
rect 56689 21975 56747 21981
rect 56597 21947 56655 21953
rect 56597 21944 56609 21947
rect 55600 21916 56609 21944
rect 56597 21913 56609 21916
rect 56643 21944 56655 21947
rect 56704 21944 56732 21975
rect 56870 21972 56876 22024
rect 56928 21972 56934 22024
rect 56965 22015 57023 22021
rect 56965 21981 56977 22015
rect 57011 21981 57023 22015
rect 56965 21975 57023 21981
rect 56643 21916 56732 21944
rect 56643 21913 56655 21916
rect 56597 21907 56655 21913
rect 56778 21904 56784 21956
rect 56836 21904 56842 21956
rect 56980 21876 57008 21975
rect 57146 21972 57152 22024
rect 57204 21972 57210 22024
rect 57716 22021 57744 22052
rect 57992 22021 58020 22052
rect 57701 22015 57759 22021
rect 57701 21981 57713 22015
rect 57747 21981 57759 22015
rect 57701 21975 57759 21981
rect 57793 22015 57851 22021
rect 57793 21981 57805 22015
rect 57839 21981 57851 22015
rect 57793 21975 57851 21981
rect 57977 22015 58035 22021
rect 57977 21981 57989 22015
rect 58023 21981 58035 22015
rect 57977 21975 58035 21981
rect 58069 22015 58127 22021
rect 58069 21981 58081 22015
rect 58115 22012 58127 22015
rect 58529 22015 58587 22021
rect 58115 21984 58480 22012
rect 58115 21981 58127 21984
rect 58069 21975 58127 21981
rect 57054 21904 57060 21956
rect 57112 21944 57118 21956
rect 57808 21944 57836 21975
rect 57112 21916 57836 21944
rect 57112 21904 57118 21916
rect 57882 21904 57888 21956
rect 57940 21904 57946 21956
rect 57992 21944 58020 21975
rect 57992 21916 58112 21944
rect 58084 21888 58112 21916
rect 57974 21876 57980 21888
rect 54956 21848 57980 21876
rect 54619 21845 54631 21848
rect 54573 21839 54631 21845
rect 57974 21836 57980 21848
rect 58032 21836 58038 21888
rect 58066 21836 58072 21888
rect 58124 21836 58130 21888
rect 58250 21836 58256 21888
rect 58308 21836 58314 21888
rect 58342 21836 58348 21888
rect 58400 21836 58406 21888
rect 58452 21876 58480 21984
rect 58529 21981 58541 22015
rect 58575 21981 58587 22015
rect 58529 21975 58587 21981
rect 58544 21944 58572 21975
rect 58894 21944 58900 21956
rect 58544 21916 58900 21944
rect 58894 21904 58900 21916
rect 58952 21904 58958 21956
rect 58710 21876 58716 21888
rect 58452 21848 58716 21876
rect 58710 21836 58716 21848
rect 58768 21836 58774 21888
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 3786 21632 3792 21684
rect 3844 21672 3850 21684
rect 4157 21675 4215 21681
rect 4157 21672 4169 21675
rect 3844 21644 4169 21672
rect 3844 21632 3850 21644
rect 4157 21641 4169 21644
rect 4203 21641 4215 21675
rect 6542 21675 6600 21681
rect 4157 21635 4215 21641
rect 4540 21644 6500 21672
rect 4540 21613 4568 21644
rect 4525 21607 4583 21613
rect 4525 21573 4537 21607
rect 4571 21573 4583 21607
rect 4525 21567 4583 21573
rect 5718 21564 5724 21616
rect 5776 21604 5782 21616
rect 6472 21604 6500 21644
rect 6542 21641 6554 21675
rect 6588 21672 6600 21675
rect 6638 21672 6644 21684
rect 6588 21644 6644 21672
rect 6588 21641 6600 21644
rect 6542 21635 6600 21641
rect 6638 21632 6644 21644
rect 6696 21632 6702 21684
rect 7006 21632 7012 21684
rect 7064 21632 7070 21684
rect 8027 21675 8085 21681
rect 8027 21641 8039 21675
rect 8073 21672 8085 21675
rect 8202 21672 8208 21684
rect 8073 21644 8208 21672
rect 8073 21641 8085 21644
rect 8027 21635 8085 21641
rect 8202 21632 8208 21644
rect 8260 21632 8266 21684
rect 42705 21675 42763 21681
rect 42705 21641 42717 21675
rect 42751 21672 42763 21675
rect 42886 21672 42892 21684
rect 42751 21644 42892 21672
rect 42751 21641 42763 21644
rect 42705 21635 42763 21641
rect 42886 21632 42892 21644
rect 42944 21632 42950 21684
rect 42978 21632 42984 21684
rect 43036 21672 43042 21684
rect 43073 21675 43131 21681
rect 43073 21672 43085 21675
rect 43036 21644 43085 21672
rect 43036 21632 43042 21644
rect 43073 21641 43085 21644
rect 43119 21641 43131 21675
rect 43073 21635 43131 21641
rect 43162 21632 43168 21684
rect 43220 21632 43226 21684
rect 43349 21675 43407 21681
rect 43349 21641 43361 21675
rect 43395 21641 43407 21675
rect 43349 21635 43407 21641
rect 7558 21604 7564 21616
rect 5776 21576 6408 21604
rect 6472 21576 7564 21604
rect 5776 21564 5782 21576
rect 2682 21496 2688 21548
rect 2740 21496 2746 21548
rect 4706 21496 4712 21548
rect 4764 21496 4770 21548
rect 4798 21496 4804 21548
rect 4856 21496 4862 21548
rect 5905 21539 5963 21545
rect 5905 21505 5917 21539
rect 5951 21505 5963 21539
rect 5905 21499 5963 21505
rect 934 21428 940 21480
rect 992 21468 998 21480
rect 1581 21471 1639 21477
rect 1581 21468 1593 21471
rect 992 21440 1593 21468
rect 992 21428 998 21440
rect 1581 21437 1593 21440
rect 1627 21437 1639 21471
rect 1581 21431 1639 21437
rect 3694 21428 3700 21480
rect 3752 21428 3758 21480
rect 4430 21428 4436 21480
rect 4488 21428 4494 21480
rect 5920 21468 5948 21499
rect 5994 21496 6000 21548
rect 6052 21496 6058 21548
rect 6380 21545 6408 21576
rect 6365 21539 6423 21545
rect 6365 21505 6377 21539
rect 6411 21505 6423 21539
rect 6365 21499 6423 21505
rect 6454 21496 6460 21548
rect 6512 21496 6518 21548
rect 6656 21545 6684 21576
rect 7558 21564 7564 21576
rect 7616 21604 7622 21616
rect 7929 21607 7987 21613
rect 7929 21604 7941 21607
rect 7616 21576 7941 21604
rect 7616 21564 7622 21576
rect 7929 21573 7941 21576
rect 7975 21573 7987 21607
rect 43180 21604 43208 21632
rect 7929 21567 7987 21573
rect 42536 21576 43208 21604
rect 6641 21539 6699 21545
rect 6641 21505 6653 21539
rect 6687 21505 6699 21539
rect 6641 21499 6699 21505
rect 7006 21496 7012 21548
rect 7064 21496 7070 21548
rect 8113 21539 8171 21545
rect 8113 21505 8125 21539
rect 8159 21505 8171 21539
rect 8113 21499 8171 21505
rect 7024 21468 7052 21496
rect 5920 21440 7052 21468
rect 4448 21400 4476 21428
rect 8128 21412 8156 21499
rect 8202 21496 8208 21548
rect 8260 21496 8266 21548
rect 42536 21545 42564 21576
rect 42521 21539 42579 21545
rect 42521 21505 42533 21539
rect 42567 21505 42579 21539
rect 42521 21499 42579 21505
rect 42705 21539 42763 21545
rect 42705 21505 42717 21539
rect 42751 21505 42763 21539
rect 42705 21499 42763 21505
rect 42797 21539 42855 21545
rect 42797 21505 42809 21539
rect 42843 21536 42855 21539
rect 43364 21536 43392 21635
rect 43530 21632 43536 21684
rect 43588 21632 43594 21684
rect 44174 21632 44180 21684
rect 44232 21672 44238 21684
rect 45462 21672 45468 21684
rect 44232 21644 45468 21672
rect 44232 21632 44238 21644
rect 45462 21632 45468 21644
rect 45520 21672 45526 21684
rect 45520 21644 46428 21672
rect 45520 21632 45526 21644
rect 42843 21508 43392 21536
rect 42843 21505 42855 21508
rect 42797 21499 42855 21505
rect 10686 21428 10692 21480
rect 10744 21428 10750 21480
rect 11517 21471 11575 21477
rect 11517 21437 11529 21471
rect 11563 21437 11575 21471
rect 42720 21468 42748 21499
rect 43073 21471 43131 21477
rect 42720 21440 42932 21468
rect 11517 21431 11575 21437
rect 4525 21403 4583 21409
rect 4525 21400 4537 21403
rect 4448 21372 4537 21400
rect 4525 21369 4537 21372
rect 4571 21369 4583 21403
rect 4525 21363 4583 21369
rect 8110 21360 8116 21412
rect 8168 21360 8174 21412
rect 9858 21360 9864 21412
rect 9916 21400 9922 21412
rect 11532 21400 11560 21431
rect 9916 21372 11560 21400
rect 9916 21360 9922 21372
rect 11974 21360 11980 21412
rect 12032 21400 12038 21412
rect 12529 21403 12587 21409
rect 12529 21400 12541 21403
rect 12032 21372 12541 21400
rect 12032 21360 12038 21372
rect 12529 21369 12541 21372
rect 12575 21400 12587 21403
rect 19978 21400 19984 21412
rect 12575 21372 19984 21400
rect 12575 21369 12587 21372
rect 12529 21363 12587 21369
rect 19978 21360 19984 21372
rect 20036 21400 20042 21412
rect 34514 21400 34520 21412
rect 20036 21372 34520 21400
rect 20036 21360 20042 21372
rect 34514 21360 34520 21372
rect 34572 21360 34578 21412
rect 42904 21344 42932 21440
rect 43073 21437 43085 21471
rect 43119 21468 43131 21471
rect 43548 21468 43576 21632
rect 44542 21564 44548 21616
rect 44600 21564 44606 21616
rect 44726 21564 44732 21616
rect 44784 21564 44790 21616
rect 46109 21607 46167 21613
rect 46109 21573 46121 21607
rect 46155 21604 46167 21607
rect 46198 21604 46204 21616
rect 46155 21576 46204 21604
rect 46155 21573 46167 21576
rect 46109 21567 46167 21573
rect 46198 21564 46204 21576
rect 46256 21564 46262 21616
rect 43901 21539 43959 21545
rect 43901 21505 43913 21539
rect 43947 21536 43959 21539
rect 43990 21536 43996 21548
rect 43947 21508 43996 21536
rect 43947 21505 43959 21508
rect 43901 21499 43959 21505
rect 43990 21496 43996 21508
rect 44048 21496 44054 21548
rect 44082 21496 44088 21548
rect 44140 21496 44146 21548
rect 44269 21539 44327 21545
rect 44269 21505 44281 21539
rect 44315 21505 44327 21539
rect 44269 21499 44327 21505
rect 43119 21440 43576 21468
rect 43625 21471 43683 21477
rect 43119 21437 43131 21440
rect 43073 21431 43131 21437
rect 43625 21437 43637 21471
rect 43671 21468 43683 21471
rect 44100 21468 44128 21496
rect 43671 21440 44128 21468
rect 43671 21437 43683 21440
rect 43625 21431 43683 21437
rect 44284 21400 44312 21499
rect 44358 21496 44364 21548
rect 44416 21496 44422 21548
rect 44545 21471 44603 21477
rect 44545 21437 44557 21471
rect 44591 21468 44603 21471
rect 44744 21468 44772 21564
rect 46400 21545 46428 21644
rect 46658 21632 46664 21684
rect 46716 21632 46722 21684
rect 49418 21632 49424 21684
rect 49476 21672 49482 21684
rect 49476 21644 50844 21672
rect 49476 21632 49482 21644
rect 46385 21539 46443 21545
rect 44591 21440 44772 21468
rect 45020 21468 45048 21522
rect 46385 21505 46397 21539
rect 46431 21505 46443 21539
rect 46385 21499 46443 21505
rect 46676 21468 46704 21632
rect 49436 21604 49464 21632
rect 50249 21607 50307 21613
rect 50249 21604 50261 21607
rect 49436 21576 49648 21604
rect 49145 21539 49203 21545
rect 49145 21505 49157 21539
rect 49191 21536 49203 21539
rect 49237 21539 49295 21545
rect 49237 21536 49249 21539
rect 49191 21508 49249 21536
rect 49191 21505 49203 21508
rect 49145 21499 49203 21505
rect 49237 21505 49249 21508
rect 49283 21505 49295 21539
rect 49237 21499 49295 21505
rect 49418 21496 49424 21548
rect 49476 21496 49482 21548
rect 49510 21496 49516 21548
rect 49568 21496 49574 21548
rect 49620 21545 49648 21576
rect 49804 21576 50261 21604
rect 49804 21545 49832 21576
rect 50249 21573 50261 21576
rect 50295 21573 50307 21607
rect 50249 21567 50307 21573
rect 50816 21604 50844 21644
rect 52178 21632 52184 21684
rect 52236 21632 52242 21684
rect 52730 21672 52736 21684
rect 52472 21644 52736 21672
rect 51074 21604 51080 21616
rect 50816 21576 51080 21604
rect 49605 21539 49663 21545
rect 49605 21505 49617 21539
rect 49651 21505 49663 21539
rect 49605 21499 49663 21505
rect 49789 21539 49847 21545
rect 49789 21505 49801 21539
rect 49835 21505 49847 21539
rect 49789 21499 49847 21505
rect 49878 21496 49884 21548
rect 49936 21496 49942 21548
rect 50065 21539 50123 21545
rect 50065 21505 50077 21539
rect 50111 21505 50123 21539
rect 50065 21499 50123 21505
rect 45020 21440 46704 21468
rect 48409 21471 48467 21477
rect 44591 21437 44603 21440
rect 44545 21431 44603 21437
rect 48409 21437 48421 21471
rect 48455 21437 48467 21471
rect 48409 21431 48467 21437
rect 48593 21471 48651 21477
rect 48593 21437 48605 21471
rect 48639 21468 48651 21471
rect 48774 21468 48780 21480
rect 48639 21440 48780 21468
rect 48639 21437 48651 21440
rect 48593 21431 48651 21437
rect 44726 21400 44732 21412
rect 44284 21372 44732 21400
rect 44726 21360 44732 21372
rect 44784 21360 44790 21412
rect 48424 21400 48452 21431
rect 48774 21428 48780 21440
rect 48832 21428 48838 21480
rect 50080 21468 50108 21499
rect 50154 21496 50160 21548
rect 50212 21496 50218 21548
rect 50341 21539 50399 21545
rect 50341 21505 50353 21539
rect 50387 21505 50399 21539
rect 50341 21499 50399 21505
rect 50080 21440 50200 21468
rect 49237 21403 49295 21409
rect 49237 21400 49249 21403
rect 48424 21372 49249 21400
rect 49237 21369 49249 21372
rect 49283 21369 49295 21403
rect 49237 21363 49295 21369
rect 49602 21360 49608 21412
rect 49660 21400 49666 21412
rect 49973 21403 50031 21409
rect 49973 21400 49985 21403
rect 49660 21372 49985 21400
rect 49660 21360 49666 21372
rect 49973 21369 49985 21372
rect 50019 21369 50031 21403
rect 49973 21363 50031 21369
rect 3050 21292 3056 21344
rect 3108 21332 3114 21344
rect 3145 21335 3203 21341
rect 3145 21332 3157 21335
rect 3108 21304 3157 21332
rect 3108 21292 3114 21304
rect 3145 21301 3157 21304
rect 3191 21301 3203 21335
rect 3145 21295 3203 21301
rect 10042 21292 10048 21344
rect 10100 21292 10106 21344
rect 12158 21292 12164 21344
rect 12216 21292 12222 21344
rect 42886 21292 42892 21344
rect 42944 21292 42950 21344
rect 43806 21292 43812 21344
rect 43864 21292 43870 21344
rect 44634 21292 44640 21344
rect 44692 21292 44698 21344
rect 47762 21292 47768 21344
rect 47820 21292 47826 21344
rect 49694 21292 49700 21344
rect 49752 21292 49758 21344
rect 50172 21332 50200 21440
rect 50356 21400 50384 21499
rect 50522 21496 50528 21548
rect 50580 21496 50586 21548
rect 50816 21545 50844 21576
rect 51074 21564 51080 21576
rect 51132 21604 51138 21616
rect 51261 21607 51319 21613
rect 51261 21604 51273 21607
rect 51132 21576 51273 21604
rect 51132 21564 51138 21576
rect 51261 21573 51273 21576
rect 51307 21573 51319 21607
rect 52196 21604 52224 21632
rect 52196 21576 52316 21604
rect 51261 21567 51319 21573
rect 50709 21539 50767 21545
rect 50709 21505 50721 21539
rect 50755 21505 50767 21539
rect 50709 21499 50767 21505
rect 50801 21539 50859 21545
rect 50801 21505 50813 21539
rect 50847 21505 50859 21539
rect 50801 21499 50859 21505
rect 50724 21468 50752 21499
rect 50982 21496 50988 21548
rect 51040 21496 51046 21548
rect 52288 21545 52316 21576
rect 52181 21539 52239 21545
rect 52181 21505 52193 21539
rect 52227 21505 52239 21539
rect 52181 21499 52239 21505
rect 52273 21539 52331 21545
rect 52273 21505 52285 21539
rect 52319 21505 52331 21539
rect 52273 21499 52331 21505
rect 50893 21471 50951 21477
rect 50893 21468 50905 21471
rect 50724 21440 50905 21468
rect 50893 21437 50905 21440
rect 50939 21437 50951 21471
rect 52196 21468 52224 21499
rect 52472 21477 52500 21644
rect 52730 21632 52736 21644
rect 52788 21632 52794 21684
rect 54110 21632 54116 21684
rect 54168 21632 54174 21684
rect 54297 21675 54355 21681
rect 54297 21641 54309 21675
rect 54343 21672 54355 21675
rect 54478 21672 54484 21684
rect 54343 21644 54484 21672
rect 54343 21641 54355 21644
rect 54297 21635 54355 21641
rect 54478 21632 54484 21644
rect 54536 21632 54542 21684
rect 55861 21675 55919 21681
rect 55861 21641 55873 21675
rect 55907 21672 55919 21675
rect 55950 21672 55956 21684
rect 55907 21644 55956 21672
rect 55907 21641 55919 21644
rect 55861 21635 55919 21641
rect 55950 21632 55956 21644
rect 56008 21632 56014 21684
rect 56778 21632 56784 21684
rect 56836 21632 56842 21684
rect 57882 21632 57888 21684
rect 57940 21632 57946 21684
rect 58066 21632 58072 21684
rect 58124 21672 58130 21684
rect 58529 21675 58587 21681
rect 58529 21672 58541 21675
rect 58124 21644 58541 21672
rect 58124 21632 58130 21644
rect 58529 21641 58541 21644
rect 58575 21641 58587 21675
rect 58529 21635 58587 21641
rect 52748 21576 56456 21604
rect 52748 21545 52776 21576
rect 52733 21539 52791 21545
rect 52733 21505 52745 21539
rect 52779 21505 52791 21539
rect 52989 21539 53047 21545
rect 52989 21536 53001 21539
rect 52733 21499 52791 21505
rect 52840 21508 53001 21536
rect 52457 21471 52515 21477
rect 52196 21440 52316 21468
rect 50893 21431 50951 21437
rect 51442 21400 51448 21412
rect 50356 21372 51448 21400
rect 51442 21360 51448 21372
rect 51500 21360 51506 21412
rect 50617 21335 50675 21341
rect 50617 21332 50629 21335
rect 50172 21304 50629 21332
rect 50617 21301 50629 21304
rect 50663 21301 50675 21335
rect 52288 21332 52316 21440
rect 52457 21437 52469 21471
rect 52503 21437 52515 21471
rect 52840 21468 52868 21508
rect 52989 21505 53001 21508
rect 53035 21505 53047 21539
rect 52989 21499 53047 21505
rect 53558 21496 53564 21548
rect 53616 21536 53622 21548
rect 54496 21545 54524 21576
rect 54754 21545 54760 21548
rect 54205 21539 54263 21545
rect 54205 21536 54217 21539
rect 53616 21508 54217 21536
rect 53616 21496 53622 21508
rect 54205 21505 54217 21508
rect 54251 21505 54263 21539
rect 54205 21499 54263 21505
rect 54481 21539 54539 21545
rect 54481 21505 54493 21539
rect 54527 21505 54539 21539
rect 54481 21499 54539 21505
rect 54748 21499 54760 21545
rect 54754 21496 54760 21499
rect 54812 21496 54818 21548
rect 56428 21480 56456 21576
rect 56597 21539 56655 21545
rect 56597 21505 56609 21539
rect 56643 21536 56655 21539
rect 56796 21536 56824 21632
rect 56643 21508 56824 21536
rect 57517 21539 57575 21545
rect 56643 21505 56655 21508
rect 56597 21499 56655 21505
rect 57517 21505 57529 21539
rect 57563 21536 57575 21539
rect 57900 21536 57928 21632
rect 57563 21508 57928 21536
rect 57563 21505 57575 21508
rect 57517 21499 57575 21505
rect 52457 21431 52515 21437
rect 52748 21440 52868 21468
rect 52365 21403 52423 21409
rect 52365 21369 52377 21403
rect 52411 21400 52423 21403
rect 52748 21400 52776 21440
rect 56410 21428 56416 21480
rect 56468 21428 56474 21480
rect 57882 21428 57888 21480
rect 57940 21428 57946 21480
rect 52411 21372 52776 21400
rect 52411 21369 52423 21372
rect 52365 21363 52423 21369
rect 55214 21332 55220 21344
rect 52288 21304 55220 21332
rect 50617 21295 50675 21301
rect 55214 21292 55220 21304
rect 55272 21292 55278 21344
rect 55398 21292 55404 21344
rect 55456 21332 55462 21344
rect 55953 21335 56011 21341
rect 55953 21332 55965 21335
rect 55456 21304 55965 21332
rect 55456 21292 55462 21304
rect 55953 21301 55965 21304
rect 55999 21301 56011 21335
rect 55953 21295 56011 21301
rect 56594 21292 56600 21344
rect 56652 21332 56658 21344
rect 56873 21335 56931 21341
rect 56873 21332 56885 21335
rect 56652 21304 56885 21332
rect 56652 21292 56658 21304
rect 56873 21301 56885 21304
rect 56919 21301 56931 21335
rect 56873 21295 56931 21301
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 3050 21088 3056 21140
rect 3108 21088 3114 21140
rect 3329 21131 3387 21137
rect 3329 21097 3341 21131
rect 3375 21128 3387 21131
rect 3694 21128 3700 21140
rect 3375 21100 3700 21128
rect 3375 21097 3387 21100
rect 3329 21091 3387 21097
rect 3694 21088 3700 21100
rect 3752 21088 3758 21140
rect 4617 21131 4675 21137
rect 4617 21097 4629 21131
rect 4663 21128 4675 21131
rect 4706 21128 4712 21140
rect 4663 21100 4712 21128
rect 4663 21097 4675 21100
rect 4617 21091 4675 21097
rect 4706 21088 4712 21100
rect 4764 21088 4770 21140
rect 6365 21131 6423 21137
rect 6365 21097 6377 21131
rect 6411 21128 6423 21131
rect 6454 21128 6460 21140
rect 6411 21100 6460 21128
rect 6411 21097 6423 21100
rect 6365 21091 6423 21097
rect 6454 21088 6460 21100
rect 6512 21088 6518 21140
rect 8110 21088 8116 21140
rect 8168 21128 8174 21140
rect 8297 21131 8355 21137
rect 8297 21128 8309 21131
rect 8168 21100 8309 21128
rect 8168 21088 8174 21100
rect 8297 21097 8309 21100
rect 8343 21097 8355 21131
rect 8297 21091 8355 21097
rect 9769 21131 9827 21137
rect 9769 21097 9781 21131
rect 9815 21128 9827 21131
rect 9858 21128 9864 21140
rect 9815 21100 9864 21128
rect 9815 21097 9827 21100
rect 9769 21091 9827 21097
rect 9858 21088 9864 21100
rect 9916 21088 9922 21140
rect 9950 21088 9956 21140
rect 10008 21088 10014 21140
rect 10042 21088 10048 21140
rect 10100 21088 10106 21140
rect 10410 21088 10416 21140
rect 10468 21088 10474 21140
rect 12158 21088 12164 21140
rect 12216 21088 12222 21140
rect 42886 21088 42892 21140
rect 42944 21128 42950 21140
rect 44358 21128 44364 21140
rect 42944 21100 44364 21128
rect 42944 21088 42950 21100
rect 44358 21088 44364 21100
rect 44416 21088 44422 21140
rect 44726 21088 44732 21140
rect 44784 21088 44790 21140
rect 45646 21088 45652 21140
rect 45704 21128 45710 21140
rect 45833 21131 45891 21137
rect 45833 21128 45845 21131
rect 45704 21100 45845 21128
rect 45704 21088 45710 21100
rect 45833 21097 45845 21100
rect 45879 21097 45891 21131
rect 45833 21091 45891 21097
rect 47762 21088 47768 21140
rect 47820 21088 47826 21140
rect 49418 21088 49424 21140
rect 49476 21088 49482 21140
rect 49602 21088 49608 21140
rect 49660 21088 49666 21140
rect 49694 21088 49700 21140
rect 49752 21088 49758 21140
rect 50433 21131 50491 21137
rect 50433 21097 50445 21131
rect 50479 21128 50491 21131
rect 50522 21128 50528 21140
rect 50479 21100 50528 21128
rect 50479 21097 50491 21100
rect 50433 21091 50491 21097
rect 50522 21088 50528 21100
rect 50580 21088 50586 21140
rect 50982 21088 50988 21140
rect 51040 21128 51046 21140
rect 51537 21131 51595 21137
rect 51537 21128 51549 21131
rect 51040 21100 51549 21128
rect 51040 21088 51046 21100
rect 51537 21097 51549 21100
rect 51583 21097 51595 21131
rect 51537 21091 51595 21097
rect 54570 21088 54576 21140
rect 54628 21088 54634 21140
rect 54754 21088 54760 21140
rect 54812 21128 54818 21140
rect 54849 21131 54907 21137
rect 54849 21128 54861 21131
rect 54812 21100 54861 21128
rect 54812 21088 54818 21100
rect 54849 21097 54861 21100
rect 54895 21097 54907 21131
rect 56594 21128 56600 21140
rect 54849 21091 54907 21097
rect 56336 21100 56600 21128
rect 2869 20995 2927 21001
rect 2869 20961 2881 20995
rect 2915 20992 2927 20995
rect 3068 20992 3096 21088
rect 9968 21060 9996 21088
rect 9600 21032 9996 21060
rect 2915 20964 3096 20992
rect 3237 20995 3295 21001
rect 2915 20961 2927 20964
rect 2869 20955 2927 20961
rect 3237 20961 3249 20995
rect 3283 20992 3295 20995
rect 3789 20995 3847 21001
rect 3789 20992 3801 20995
rect 3283 20964 3801 20992
rect 3283 20961 3295 20964
rect 3237 20955 3295 20961
rect 3789 20961 3801 20964
rect 3835 20961 3847 20995
rect 3789 20955 3847 20961
rect 3142 20884 3148 20936
rect 3200 20884 3206 20936
rect 3421 20927 3479 20933
rect 3421 20893 3433 20927
rect 3467 20893 3479 20927
rect 3421 20887 3479 20893
rect 2406 20816 2412 20868
rect 2464 20816 2470 20868
rect 2866 20816 2872 20868
rect 2924 20856 2930 20868
rect 3436 20856 3464 20887
rect 3510 20884 3516 20936
rect 3568 20884 3574 20936
rect 4338 20884 4344 20936
rect 4396 20884 4402 20936
rect 4985 20927 5043 20933
rect 4985 20924 4997 20927
rect 4632 20896 4997 20924
rect 4632 20868 4660 20896
rect 4985 20893 4997 20896
rect 5031 20924 5043 20927
rect 5350 20924 5356 20936
rect 5031 20896 5356 20924
rect 5031 20893 5043 20896
rect 4985 20887 5043 20893
rect 5350 20884 5356 20896
rect 5408 20884 5414 20936
rect 9600 20933 9628 21032
rect 9861 20995 9919 21001
rect 9861 20961 9873 20995
rect 9907 20992 9919 20995
rect 10060 20992 10088 21088
rect 9907 20964 10088 20992
rect 9907 20961 9919 20964
rect 9861 20955 9919 20961
rect 6549 20927 6607 20933
rect 6549 20893 6561 20927
rect 6595 20924 6607 20927
rect 9585 20927 9643 20933
rect 6595 20896 8892 20924
rect 6595 20893 6607 20896
rect 6549 20887 6607 20893
rect 2924 20828 3464 20856
rect 2924 20816 2930 20828
rect 4614 20816 4620 20868
rect 4672 20816 4678 20868
rect 4801 20859 4859 20865
rect 4801 20825 4813 20859
rect 4847 20825 4859 20859
rect 5368 20856 5396 20884
rect 8864 20868 8892 20896
rect 9585 20893 9597 20927
rect 9631 20893 9643 20927
rect 9585 20887 9643 20893
rect 9677 20927 9735 20933
rect 9677 20893 9689 20927
rect 9723 20924 9735 20927
rect 9950 20924 9956 20936
rect 9723 20896 9956 20924
rect 9723 20893 9735 20896
rect 9677 20887 9735 20893
rect 9950 20884 9956 20896
rect 10008 20924 10014 20936
rect 10428 20924 10456 21088
rect 12176 21060 12204 21088
rect 11808 21032 12204 21060
rect 43548 21032 44036 21060
rect 11609 20995 11667 21001
rect 11609 20961 11621 20995
rect 11655 20992 11667 20995
rect 11808 20992 11836 21032
rect 11655 20964 11836 20992
rect 11885 20995 11943 21001
rect 11655 20961 11667 20964
rect 11609 20955 11667 20961
rect 11885 20961 11897 20995
rect 11931 20992 11943 20995
rect 11974 20992 11980 21004
rect 11931 20964 11980 20992
rect 11931 20961 11943 20964
rect 11885 20955 11943 20961
rect 11974 20952 11980 20964
rect 12032 20952 12038 21004
rect 43548 21001 43576 21032
rect 44008 21004 44036 21032
rect 43533 20995 43591 21001
rect 43533 20961 43545 20995
rect 43579 20961 43591 20995
rect 43533 20955 43591 20961
rect 43809 20995 43867 21001
rect 43809 20961 43821 20995
rect 43855 20961 43867 20995
rect 43809 20955 43867 20961
rect 10008 20896 10456 20924
rect 10008 20884 10014 20896
rect 13722 20884 13728 20936
rect 13780 20924 13786 20936
rect 14277 20927 14335 20933
rect 14277 20924 14289 20927
rect 13780 20896 14289 20924
rect 13780 20884 13786 20896
rect 14277 20893 14289 20896
rect 14323 20924 14335 20927
rect 18230 20924 18236 20936
rect 14323 20896 18236 20924
rect 14323 20893 14335 20896
rect 14277 20887 14335 20893
rect 18230 20884 18236 20896
rect 18288 20884 18294 20936
rect 43438 20884 43444 20936
rect 43496 20884 43502 20936
rect 43824 20924 43852 20955
rect 43990 20952 43996 21004
rect 44048 20952 44054 21004
rect 44376 20992 44404 21088
rect 44376 20964 45140 20992
rect 44361 20927 44419 20933
rect 44361 20924 44373 20927
rect 43824 20896 44373 20924
rect 44361 20893 44373 20896
rect 44407 20893 44419 20927
rect 44361 20887 44419 20893
rect 44634 20884 44640 20936
rect 44692 20924 44698 20936
rect 45005 20927 45063 20933
rect 45005 20924 45017 20927
rect 44692 20896 45017 20924
rect 44692 20884 44698 20896
rect 45005 20893 45017 20896
rect 45051 20893 45063 20927
rect 45112 20924 45140 20964
rect 45462 20952 45468 21004
rect 45520 20992 45526 21004
rect 46201 20995 46259 21001
rect 46201 20992 46213 20995
rect 45520 20964 46213 20992
rect 45520 20952 45526 20964
rect 46201 20961 46213 20964
rect 46247 20961 46259 20995
rect 46201 20955 46259 20961
rect 45741 20927 45799 20933
rect 45741 20924 45753 20927
rect 45112 20896 45753 20924
rect 45005 20887 45063 20893
rect 45741 20893 45753 20896
rect 45787 20893 45799 20927
rect 45741 20887 45799 20893
rect 45925 20927 45983 20933
rect 45925 20893 45937 20927
rect 45971 20893 45983 20927
rect 46216 20924 46244 20955
rect 47026 20924 47032 20936
rect 46216 20896 47032 20924
rect 45925 20887 45983 20893
rect 6733 20859 6791 20865
rect 6733 20856 6745 20859
rect 5368 20828 6745 20856
rect 4801 20819 4859 20825
rect 6733 20825 6745 20828
rect 6779 20856 6791 20859
rect 6914 20856 6920 20868
rect 6779 20828 6920 20856
rect 6779 20825 6791 20828
rect 6733 20819 6791 20825
rect 1397 20791 1455 20797
rect 1397 20757 1409 20791
rect 1443 20788 1455 20791
rect 2682 20788 2688 20800
rect 1443 20760 2688 20788
rect 1443 20757 1455 20760
rect 1397 20751 1455 20757
rect 2682 20748 2688 20760
rect 2740 20748 2746 20800
rect 4816 20788 4844 20819
rect 6914 20816 6920 20828
rect 6972 20816 6978 20868
rect 8018 20816 8024 20868
rect 8076 20816 8082 20868
rect 8481 20859 8539 20865
rect 8481 20825 8493 20859
rect 8527 20825 8539 20859
rect 8481 20819 8539 20825
rect 8036 20788 8064 20816
rect 4816 20760 8064 20788
rect 8496 20788 8524 20819
rect 8570 20816 8576 20868
rect 8628 20856 8634 20868
rect 8665 20859 8723 20865
rect 8665 20856 8677 20859
rect 8628 20828 8677 20856
rect 8628 20816 8634 20828
rect 8665 20825 8677 20828
rect 8711 20825 8723 20859
rect 8665 20819 8723 20825
rect 8846 20816 8852 20868
rect 8904 20816 8910 20868
rect 9766 20816 9772 20868
rect 9824 20856 9830 20868
rect 9824 20828 10272 20856
rect 9824 20816 9830 20828
rect 10042 20788 10048 20800
rect 8496 20760 10048 20788
rect 10042 20748 10048 20760
rect 10100 20748 10106 20800
rect 10134 20748 10140 20800
rect 10192 20748 10198 20800
rect 10244 20788 10272 20828
rect 10962 20816 10968 20868
rect 11020 20816 11026 20868
rect 11977 20859 12035 20865
rect 11977 20825 11989 20859
rect 12023 20825 12035 20859
rect 11977 20819 12035 20825
rect 11992 20788 12020 20819
rect 10244 20760 12020 20788
rect 43456 20788 43484 20884
rect 44082 20816 44088 20868
rect 44140 20856 44146 20868
rect 44545 20859 44603 20865
rect 44545 20856 44557 20859
rect 44140 20828 44557 20856
rect 44140 20816 44146 20828
rect 44545 20825 44557 20828
rect 44591 20825 44603 20859
rect 45940 20856 45968 20887
rect 47026 20884 47032 20896
rect 47084 20884 47090 20936
rect 44545 20819 44603 20825
rect 45204 20828 45968 20856
rect 46468 20859 46526 20865
rect 45204 20797 45232 20828
rect 46468 20825 46480 20859
rect 46514 20856 46526 20859
rect 47780 20856 47808 21088
rect 49050 21020 49056 21072
rect 49108 21060 49114 21072
rect 49108 21032 49372 21060
rect 49108 21020 49114 21032
rect 47946 20952 47952 21004
rect 48004 20992 48010 21004
rect 48004 20964 49280 20992
rect 48004 20952 48010 20964
rect 47857 20927 47915 20933
rect 47857 20893 47869 20927
rect 47903 20893 47915 20927
rect 47857 20887 47915 20893
rect 46514 20828 47808 20856
rect 46514 20825 46526 20828
rect 46468 20819 46526 20825
rect 45189 20791 45247 20797
rect 45189 20788 45201 20791
rect 43456 20760 45201 20788
rect 45189 20757 45201 20760
rect 45235 20757 45247 20791
rect 45189 20751 45247 20757
rect 47118 20748 47124 20800
rect 47176 20788 47182 20800
rect 47581 20791 47639 20797
rect 47581 20788 47593 20791
rect 47176 20760 47593 20788
rect 47176 20748 47182 20760
rect 47581 20757 47593 20760
rect 47627 20788 47639 20791
rect 47872 20788 47900 20887
rect 48314 20884 48320 20936
rect 48372 20924 48378 20936
rect 49145 20927 49203 20933
rect 49145 20924 49157 20927
rect 48372 20896 49157 20924
rect 48372 20884 48378 20896
rect 49145 20893 49157 20896
rect 49191 20893 49203 20927
rect 49145 20887 49203 20893
rect 48406 20816 48412 20868
rect 48464 20856 48470 20868
rect 48593 20859 48651 20865
rect 48593 20856 48605 20859
rect 48464 20828 48605 20856
rect 48464 20816 48470 20828
rect 48593 20825 48605 20828
rect 48639 20825 48651 20859
rect 48593 20819 48651 20825
rect 47627 20760 47900 20788
rect 47627 20757 47639 20760
rect 47581 20751 47639 20757
rect 48498 20748 48504 20800
rect 48556 20748 48562 20800
rect 49252 20788 49280 20964
rect 49344 20933 49372 21032
rect 49329 20927 49387 20933
rect 49329 20893 49341 20927
rect 49375 20893 49387 20927
rect 49329 20887 49387 20893
rect 49436 20856 49464 21088
rect 49620 20992 49648 21088
rect 49528 20964 49648 20992
rect 49528 20933 49556 20964
rect 49513 20927 49571 20933
rect 49513 20893 49525 20927
rect 49559 20893 49571 20927
rect 49513 20887 49571 20893
rect 49605 20927 49663 20933
rect 49605 20893 49617 20927
rect 49651 20924 49663 20927
rect 49712 20924 49740 21088
rect 54588 21060 54616 21088
rect 54941 21063 54999 21069
rect 54941 21060 54953 21063
rect 54588 21032 54953 21060
rect 54941 21029 54953 21032
rect 54987 21060 54999 21063
rect 56137 21063 56195 21069
rect 56137 21060 56149 21063
rect 54987 21032 56149 21060
rect 54987 21029 54999 21032
rect 54941 21023 54999 21029
rect 56137 21029 56149 21032
rect 56183 21029 56195 21063
rect 56137 21023 56195 21029
rect 50062 20952 50068 21004
rect 50120 20992 50126 21004
rect 54757 20995 54815 21001
rect 50120 20964 50660 20992
rect 50120 20952 50126 20964
rect 49651 20896 49740 20924
rect 49789 20927 49847 20933
rect 49651 20893 49663 20896
rect 49605 20887 49663 20893
rect 49789 20893 49801 20927
rect 49835 20893 49847 20927
rect 49789 20887 49847 20893
rect 49697 20859 49755 20865
rect 49697 20856 49709 20859
rect 49436 20828 49709 20856
rect 49697 20825 49709 20828
rect 49743 20825 49755 20859
rect 49804 20856 49832 20887
rect 49970 20884 49976 20936
rect 50028 20924 50034 20936
rect 50356 20933 50384 20964
rect 50632 20933 50660 20964
rect 54757 20961 54769 20995
rect 54803 20992 54815 20995
rect 55398 20992 55404 21004
rect 54803 20964 55404 20992
rect 54803 20961 54815 20964
rect 54757 20955 54815 20961
rect 55398 20952 55404 20964
rect 55456 20952 55462 21004
rect 56336 21001 56364 21100
rect 56594 21088 56600 21100
rect 56652 21088 56658 21140
rect 57422 21088 57428 21140
rect 57480 21088 57486 21140
rect 57793 21131 57851 21137
rect 57793 21097 57805 21131
rect 57839 21128 57851 21131
rect 57882 21128 57888 21140
rect 57839 21100 57888 21128
rect 57839 21097 57851 21100
rect 57793 21091 57851 21097
rect 57882 21088 57888 21100
rect 57940 21088 57946 21140
rect 57440 21060 57468 21088
rect 58069 21063 58127 21069
rect 58069 21060 58081 21063
rect 57440 21032 58081 21060
rect 58069 21029 58081 21032
rect 58115 21029 58127 21063
rect 58069 21023 58127 21029
rect 56321 20995 56379 21001
rect 56321 20961 56333 20995
rect 56367 20961 56379 20995
rect 56321 20955 56379 20961
rect 50157 20927 50215 20933
rect 50157 20924 50169 20927
rect 50028 20896 50169 20924
rect 50028 20884 50034 20896
rect 50157 20893 50169 20896
rect 50203 20893 50215 20927
rect 50157 20887 50215 20893
rect 50341 20927 50399 20933
rect 50341 20893 50353 20927
rect 50387 20893 50399 20927
rect 50341 20887 50399 20893
rect 50433 20927 50491 20933
rect 50433 20893 50445 20927
rect 50479 20893 50491 20927
rect 50433 20887 50491 20893
rect 50617 20927 50675 20933
rect 50617 20893 50629 20927
rect 50663 20924 50675 20927
rect 50982 20924 50988 20936
rect 50663 20896 50988 20924
rect 50663 20893 50675 20896
rect 50617 20887 50675 20893
rect 50249 20859 50307 20865
rect 50249 20856 50261 20859
rect 49804 20828 50261 20856
rect 49697 20819 49755 20825
rect 50249 20825 50261 20828
rect 50295 20825 50307 20859
rect 50448 20856 50476 20887
rect 50982 20884 50988 20896
rect 51040 20884 51046 20936
rect 51442 20884 51448 20936
rect 51500 20884 51506 20936
rect 51629 20927 51687 20933
rect 51629 20893 51641 20927
rect 51675 20924 51687 20927
rect 52270 20924 52276 20936
rect 51675 20896 52276 20924
rect 51675 20893 51687 20896
rect 51629 20887 51687 20893
rect 52270 20884 52276 20896
rect 52328 20884 52334 20936
rect 55033 20927 55091 20933
rect 55033 20893 55045 20927
rect 55079 20924 55091 20927
rect 55858 20924 55864 20936
rect 55079 20896 55864 20924
rect 55079 20893 55091 20896
rect 55033 20887 55091 20893
rect 55858 20884 55864 20896
rect 55916 20884 55922 20936
rect 55950 20884 55956 20936
rect 56008 20884 56014 20936
rect 56045 20927 56103 20933
rect 56045 20893 56057 20927
rect 56091 20893 56103 20927
rect 56045 20887 56103 20893
rect 50706 20856 50712 20868
rect 50448 20828 50712 20856
rect 50249 20819 50307 20825
rect 50706 20816 50712 20828
rect 50764 20816 50770 20868
rect 49421 20791 49479 20797
rect 49421 20788 49433 20791
rect 49252 20760 49433 20788
rect 49421 20757 49433 20760
rect 49467 20757 49479 20791
rect 49421 20751 49479 20757
rect 55122 20748 55128 20800
rect 55180 20788 55186 20800
rect 55309 20791 55367 20797
rect 55309 20788 55321 20791
rect 55180 20760 55321 20788
rect 55180 20748 55186 20760
rect 55309 20757 55321 20760
rect 55355 20757 55367 20791
rect 56060 20788 56088 20887
rect 56410 20884 56416 20936
rect 56468 20884 56474 20936
rect 57974 20884 57980 20936
rect 58032 20884 58038 20936
rect 58161 20927 58219 20933
rect 58161 20893 58173 20927
rect 58207 20893 58219 20927
rect 58161 20887 58219 20893
rect 58253 20927 58311 20933
rect 58253 20893 58265 20927
rect 58299 20924 58311 20927
rect 58342 20924 58348 20936
rect 58299 20896 58348 20924
rect 58299 20893 58311 20896
rect 58253 20887 58311 20893
rect 56321 20859 56379 20865
rect 56321 20825 56333 20859
rect 56367 20856 56379 20859
rect 56658 20859 56716 20865
rect 56658 20856 56670 20859
rect 56367 20828 56670 20856
rect 56367 20825 56379 20828
rect 56321 20819 56379 20825
rect 56658 20825 56670 20828
rect 56704 20825 56716 20859
rect 58176 20856 58204 20887
rect 58342 20884 58348 20896
rect 58400 20884 58406 20936
rect 56658 20819 56716 20825
rect 57992 20828 58204 20856
rect 57992 20788 58020 20828
rect 56060 20760 58020 20788
rect 58176 20788 58204 20828
rect 58345 20791 58403 20797
rect 58345 20788 58357 20791
rect 58176 20760 58357 20788
rect 55309 20751 55367 20757
rect 58345 20757 58357 20760
rect 58391 20757 58403 20791
rect 58345 20751 58403 20757
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 3973 20587 4031 20593
rect 3973 20553 3985 20587
rect 4019 20584 4031 20587
rect 4338 20584 4344 20596
rect 4019 20556 4344 20584
rect 4019 20553 4031 20556
rect 3973 20547 4031 20553
rect 4338 20544 4344 20556
rect 4396 20544 4402 20596
rect 6454 20544 6460 20596
rect 6512 20584 6518 20596
rect 6549 20587 6607 20593
rect 6549 20584 6561 20587
rect 6512 20556 6561 20584
rect 6512 20544 6518 20556
rect 6549 20553 6561 20556
rect 6595 20553 6607 20587
rect 6549 20547 6607 20553
rect 6914 20544 6920 20596
rect 6972 20544 6978 20596
rect 8110 20544 8116 20596
rect 8168 20544 8174 20596
rect 8202 20544 8208 20596
rect 8260 20544 8266 20596
rect 10686 20544 10692 20596
rect 10744 20584 10750 20596
rect 10965 20587 11023 20593
rect 10965 20584 10977 20587
rect 10744 20556 10977 20584
rect 10744 20544 10750 20556
rect 10965 20553 10977 20556
rect 11011 20553 11023 20587
rect 10965 20547 11023 20553
rect 13170 20544 13176 20596
rect 13228 20544 13234 20596
rect 19705 20587 19763 20593
rect 19705 20553 19717 20587
rect 19751 20584 19763 20587
rect 19978 20584 19984 20596
rect 19751 20556 19984 20584
rect 19751 20553 19763 20556
rect 19705 20547 19763 20553
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 47305 20587 47363 20593
rect 47305 20553 47317 20587
rect 47351 20584 47363 20587
rect 48222 20584 48228 20596
rect 47351 20556 48228 20584
rect 47351 20553 47363 20556
rect 47305 20547 47363 20553
rect 48222 20544 48228 20556
rect 48280 20544 48286 20596
rect 48498 20544 48504 20596
rect 48556 20544 48562 20596
rect 48774 20544 48780 20596
rect 48832 20544 48838 20596
rect 49142 20544 49148 20596
rect 49200 20584 49206 20596
rect 49326 20584 49332 20596
rect 49200 20556 49332 20584
rect 49200 20544 49206 20556
rect 49326 20544 49332 20556
rect 49384 20584 49390 20596
rect 49421 20587 49479 20593
rect 49421 20584 49433 20587
rect 49384 20556 49433 20584
rect 49384 20544 49390 20556
rect 49421 20553 49433 20556
rect 49467 20553 49479 20587
rect 49421 20547 49479 20553
rect 49694 20544 49700 20596
rect 49752 20584 49758 20596
rect 50614 20584 50620 20596
rect 49752 20556 50620 20584
rect 49752 20544 49758 20556
rect 50614 20544 50620 20556
rect 50672 20544 50678 20596
rect 51442 20544 51448 20596
rect 51500 20584 51506 20596
rect 51905 20587 51963 20593
rect 51905 20584 51917 20587
rect 51500 20556 51917 20584
rect 51500 20544 51506 20556
rect 51905 20553 51917 20556
rect 51951 20553 51963 20587
rect 51905 20547 51963 20553
rect 55858 20544 55864 20596
rect 55916 20544 55922 20596
rect 55950 20544 55956 20596
rect 56008 20584 56014 20596
rect 56321 20587 56379 20593
rect 56321 20584 56333 20587
rect 56008 20556 56333 20584
rect 56008 20544 56014 20556
rect 56321 20553 56333 20556
rect 56367 20553 56379 20587
rect 56321 20547 56379 20553
rect 3329 20519 3387 20525
rect 3329 20485 3341 20519
rect 3375 20516 3387 20519
rect 6932 20516 6960 20544
rect 8220 20516 8248 20544
rect 8570 20516 8576 20528
rect 3375 20488 3832 20516
rect 3375 20485 3387 20488
rect 3329 20479 3387 20485
rect 2682 20408 2688 20460
rect 2740 20408 2746 20460
rect 3804 20457 3832 20488
rect 5920 20488 6776 20516
rect 5920 20460 5948 20488
rect 3513 20451 3571 20457
rect 3513 20417 3525 20451
rect 3559 20417 3571 20451
rect 3513 20411 3571 20417
rect 3697 20451 3755 20457
rect 3697 20417 3709 20451
rect 3743 20417 3755 20451
rect 3697 20411 3755 20417
rect 3789 20451 3847 20457
rect 3789 20417 3801 20451
rect 3835 20417 3847 20451
rect 3789 20411 3847 20417
rect 3528 20312 3556 20411
rect 3712 20380 3740 20411
rect 3970 20408 3976 20460
rect 4028 20408 4034 20460
rect 5074 20408 5080 20460
rect 5132 20448 5138 20460
rect 5362 20451 5420 20457
rect 5362 20448 5374 20451
rect 5132 20420 5374 20448
rect 5132 20408 5138 20420
rect 5362 20417 5374 20420
rect 5408 20417 5420 20451
rect 5362 20411 5420 20417
rect 5902 20408 5908 20460
rect 5960 20408 5966 20460
rect 6748 20457 6776 20488
rect 6932 20488 8576 20516
rect 6932 20457 6960 20488
rect 6365 20451 6423 20457
rect 6365 20448 6377 20451
rect 6288 20420 6377 20448
rect 4614 20380 4620 20392
rect 3712 20352 4620 20380
rect 4614 20340 4620 20352
rect 4672 20340 4678 20392
rect 5629 20383 5687 20389
rect 5629 20349 5641 20383
rect 5675 20380 5687 20383
rect 5675 20352 5856 20380
rect 5675 20349 5687 20352
rect 5629 20343 5687 20349
rect 3878 20312 3884 20324
rect 3528 20284 3884 20312
rect 3878 20272 3884 20284
rect 3936 20312 3942 20324
rect 4249 20315 4307 20321
rect 4249 20312 4261 20315
rect 3936 20284 4261 20312
rect 3936 20272 3942 20284
rect 4249 20281 4261 20284
rect 4295 20281 4307 20315
rect 4249 20275 4307 20281
rect 5828 20256 5856 20352
rect 6288 20312 6316 20420
rect 6365 20417 6377 20420
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 6641 20451 6699 20457
rect 6641 20417 6653 20451
rect 6687 20417 6699 20451
rect 6641 20411 6699 20417
rect 6733 20451 6791 20457
rect 6733 20417 6745 20451
rect 6779 20417 6791 20451
rect 6733 20411 6791 20417
rect 6917 20451 6975 20457
rect 6917 20417 6929 20451
rect 6963 20417 6975 20451
rect 6917 20411 6975 20417
rect 7929 20451 7987 20457
rect 7929 20417 7941 20451
rect 7975 20417 7987 20451
rect 7929 20411 7987 20417
rect 8205 20451 8263 20457
rect 8205 20417 8217 20451
rect 8251 20417 8263 20451
rect 8205 20411 8263 20417
rect 6656 20380 6684 20411
rect 6825 20383 6883 20389
rect 6825 20380 6837 20383
rect 6656 20352 6837 20380
rect 6825 20349 6837 20352
rect 6871 20349 6883 20383
rect 6825 20343 6883 20349
rect 7944 20312 7972 20411
rect 8220 20380 8248 20411
rect 8294 20408 8300 20460
rect 8352 20408 8358 20460
rect 8496 20457 8524 20488
rect 8570 20476 8576 20488
rect 8628 20476 8634 20528
rect 11238 20516 11244 20528
rect 11072 20488 11244 20516
rect 11072 20457 11100 20488
rect 11238 20476 11244 20488
rect 11296 20476 11302 20528
rect 12897 20519 12955 20525
rect 12897 20485 12909 20519
rect 12943 20516 12955 20519
rect 13188 20516 13216 20544
rect 47581 20519 47639 20525
rect 47581 20516 47593 20519
rect 12943 20488 13216 20516
rect 47228 20488 47593 20516
rect 12943 20485 12955 20488
rect 12897 20479 12955 20485
rect 8481 20451 8539 20457
rect 8481 20417 8493 20451
rect 8527 20417 8539 20451
rect 8481 20411 8539 20417
rect 10781 20451 10839 20457
rect 10781 20417 10793 20451
rect 10827 20448 10839 20451
rect 10873 20451 10931 20457
rect 10873 20448 10885 20451
rect 10827 20420 10885 20448
rect 10827 20417 10839 20420
rect 10781 20411 10839 20417
rect 10873 20417 10885 20420
rect 10919 20417 10931 20451
rect 10873 20411 10931 20417
rect 11057 20451 11115 20457
rect 11057 20417 11069 20451
rect 11103 20417 11115 20451
rect 11057 20411 11115 20417
rect 18230 20408 18236 20460
rect 18288 20448 18294 20460
rect 47228 20457 47256 20488
rect 47581 20485 47593 20488
rect 47627 20485 47639 20519
rect 47581 20479 47639 20485
rect 48317 20519 48375 20525
rect 48317 20485 48329 20519
rect 48363 20516 48375 20519
rect 48406 20516 48412 20528
rect 48363 20488 48412 20516
rect 48363 20485 48375 20488
rect 48317 20479 48375 20485
rect 48406 20476 48412 20488
rect 48464 20476 48470 20528
rect 48516 20516 48544 20544
rect 48516 20488 48728 20516
rect 47213 20451 47271 20457
rect 18288 20420 20392 20448
rect 18288 20408 18294 20420
rect 8389 20383 8447 20389
rect 8389 20380 8401 20383
rect 8220 20352 8401 20380
rect 8389 20349 8401 20352
rect 8435 20349 8447 20383
rect 8389 20343 8447 20349
rect 10134 20340 10140 20392
rect 10192 20340 10198 20392
rect 10318 20340 10324 20392
rect 10376 20380 10382 20392
rect 10962 20380 10968 20392
rect 10376 20352 10968 20380
rect 10376 20340 10382 20352
rect 10962 20340 10968 20352
rect 11020 20380 11026 20392
rect 12069 20383 12127 20389
rect 12069 20380 12081 20383
rect 11020 20352 12081 20380
rect 11020 20340 11026 20352
rect 12069 20349 12081 20352
rect 12115 20349 12127 20383
rect 12069 20343 12127 20349
rect 10594 20312 10600 20324
rect 6288 20284 10600 20312
rect 6288 20256 6316 20284
rect 10594 20272 10600 20284
rect 10652 20272 10658 20324
rect 3605 20247 3663 20253
rect 3605 20213 3617 20247
rect 3651 20244 3663 20247
rect 4614 20244 4620 20256
rect 3651 20216 4620 20244
rect 3651 20213 3663 20216
rect 3605 20207 3663 20213
rect 4614 20204 4620 20216
rect 4672 20204 4678 20256
rect 5810 20204 5816 20256
rect 5868 20204 5874 20256
rect 6270 20204 6276 20256
rect 6328 20204 6334 20256
rect 6365 20247 6423 20253
rect 6365 20213 6377 20247
rect 6411 20244 6423 20247
rect 6730 20244 6736 20256
rect 6411 20216 6736 20244
rect 6411 20213 6423 20216
rect 6365 20207 6423 20213
rect 6730 20204 6736 20216
rect 6788 20204 6794 20256
rect 7926 20204 7932 20256
rect 7984 20204 7990 20256
rect 8018 20204 8024 20256
rect 8076 20244 8082 20256
rect 9030 20244 9036 20256
rect 8076 20216 9036 20244
rect 8076 20204 8082 20216
rect 9030 20204 9036 20216
rect 9088 20204 9094 20256
rect 20364 20253 20392 20420
rect 47213 20417 47225 20451
rect 47259 20417 47271 20451
rect 47213 20411 47271 20417
rect 47397 20451 47455 20457
rect 47397 20417 47409 20451
rect 47443 20448 47455 20451
rect 47443 20420 48268 20448
rect 47443 20417 47455 20420
rect 47397 20411 47455 20417
rect 48133 20383 48191 20389
rect 48133 20380 48145 20383
rect 47044 20352 48145 20380
rect 20349 20247 20407 20253
rect 20349 20213 20361 20247
rect 20395 20244 20407 20247
rect 31110 20244 31116 20256
rect 20395 20216 31116 20244
rect 20395 20213 20407 20216
rect 20349 20207 20407 20213
rect 31110 20204 31116 20216
rect 31168 20204 31174 20256
rect 45738 20204 45744 20256
rect 45796 20244 45802 20256
rect 47044 20253 47072 20352
rect 48133 20349 48145 20352
rect 48179 20349 48191 20383
rect 48240 20380 48268 20420
rect 48498 20408 48504 20460
rect 48556 20408 48562 20460
rect 48590 20408 48596 20460
rect 48648 20408 48654 20460
rect 48700 20457 48728 20488
rect 53006 20476 53012 20528
rect 53064 20476 53070 20528
rect 55876 20516 55904 20544
rect 57146 20516 57152 20528
rect 55876 20488 57152 20516
rect 57146 20476 57152 20488
rect 57204 20516 57210 20528
rect 57333 20519 57391 20525
rect 57333 20516 57345 20519
rect 57204 20488 57345 20516
rect 57204 20476 57210 20488
rect 57333 20485 57345 20488
rect 57379 20485 57391 20519
rect 57333 20479 57391 20485
rect 48685 20451 48743 20457
rect 48685 20417 48697 20451
rect 48731 20417 48743 20451
rect 48685 20411 48743 20417
rect 48869 20451 48927 20457
rect 48869 20417 48881 20451
rect 48915 20448 48927 20451
rect 51819 20451 51877 20457
rect 48915 20420 48949 20448
rect 48915 20417 48927 20420
rect 48869 20411 48927 20417
rect 51819 20417 51831 20451
rect 51865 20417 51877 20451
rect 51819 20411 51877 20417
rect 51997 20451 52055 20457
rect 51997 20417 52009 20451
rect 52043 20417 52055 20451
rect 51997 20411 52055 20417
rect 52549 20451 52607 20457
rect 52549 20417 52561 20451
rect 52595 20448 52607 20451
rect 52733 20451 52791 20457
rect 52733 20448 52745 20451
rect 52595 20420 52745 20448
rect 52595 20417 52607 20420
rect 52549 20411 52607 20417
rect 52733 20417 52745 20420
rect 52779 20448 52791 20451
rect 52822 20448 52828 20460
rect 52779 20420 52828 20448
rect 52779 20417 52791 20420
rect 52733 20411 52791 20417
rect 48884 20380 48912 20411
rect 49050 20380 49056 20392
rect 48240 20352 49056 20380
rect 48133 20343 48191 20349
rect 49050 20340 49056 20352
rect 49108 20380 49114 20392
rect 49418 20380 49424 20392
rect 49108 20352 49424 20380
rect 49108 20340 49114 20352
rect 49418 20340 49424 20352
rect 49476 20340 49482 20392
rect 51828 20256 51856 20411
rect 52012 20312 52040 20411
rect 52822 20408 52828 20420
rect 52880 20408 52886 20460
rect 56229 20451 56287 20457
rect 56229 20448 56241 20451
rect 55508 20420 56241 20448
rect 52012 20284 52960 20312
rect 52932 20256 52960 20284
rect 47029 20247 47087 20253
rect 47029 20244 47041 20247
rect 45796 20216 47041 20244
rect 45796 20204 45802 20216
rect 47029 20213 47041 20216
rect 47075 20213 47087 20247
rect 47029 20207 47087 20213
rect 48314 20204 48320 20256
rect 48372 20204 48378 20256
rect 51810 20204 51816 20256
rect 51868 20204 51874 20256
rect 52914 20204 52920 20256
rect 52972 20204 52978 20256
rect 54294 20204 54300 20256
rect 54352 20244 54358 20256
rect 55508 20253 55536 20420
rect 56229 20417 56241 20420
rect 56275 20417 56287 20451
rect 56229 20411 56287 20417
rect 56318 20408 56324 20460
rect 56376 20448 56382 20460
rect 56413 20451 56471 20457
rect 56413 20448 56425 20451
rect 56376 20420 56425 20448
rect 56376 20408 56382 20420
rect 56413 20417 56425 20420
rect 56459 20417 56471 20451
rect 56413 20411 56471 20417
rect 57425 20451 57483 20457
rect 57425 20417 57437 20451
rect 57471 20448 57483 20451
rect 57701 20451 57759 20457
rect 57471 20420 57560 20448
rect 57471 20417 57483 20420
rect 57425 20411 57483 20417
rect 56137 20383 56195 20389
rect 56137 20349 56149 20383
rect 56183 20380 56195 20383
rect 56686 20380 56692 20392
rect 56183 20352 56692 20380
rect 56183 20349 56195 20352
rect 56137 20343 56195 20349
rect 56686 20340 56692 20352
rect 56744 20340 56750 20392
rect 57532 20321 57560 20420
rect 57701 20417 57713 20451
rect 57747 20417 57759 20451
rect 57701 20411 57759 20417
rect 57517 20315 57575 20321
rect 57517 20281 57529 20315
rect 57563 20281 57575 20315
rect 57716 20312 57744 20411
rect 58529 20383 58587 20389
rect 58529 20349 58541 20383
rect 58575 20380 58587 20383
rect 58575 20352 58940 20380
rect 58575 20349 58587 20352
rect 58529 20343 58587 20349
rect 57716 20284 58572 20312
rect 57517 20275 57575 20281
rect 58544 20256 58572 20284
rect 55493 20247 55551 20253
rect 55493 20244 55505 20247
rect 54352 20216 55505 20244
rect 54352 20204 54358 20216
rect 55493 20213 55505 20216
rect 55539 20213 55551 20247
rect 55493 20207 55551 20213
rect 57790 20204 57796 20256
rect 57848 20244 57854 20256
rect 57885 20247 57943 20253
rect 57885 20244 57897 20247
rect 57848 20216 57897 20244
rect 57848 20204 57854 20216
rect 57885 20213 57897 20216
rect 57931 20213 57943 20247
rect 57885 20207 57943 20213
rect 58526 20204 58532 20256
rect 58584 20204 58590 20256
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 3878 20000 3884 20052
rect 3936 20040 3942 20052
rect 4154 20040 4160 20052
rect 3936 20012 4160 20040
rect 3936 20000 3942 20012
rect 4154 20000 4160 20012
rect 4212 20000 4218 20052
rect 4709 20043 4767 20049
rect 4709 20009 4721 20043
rect 4755 20040 4767 20043
rect 5074 20040 5080 20052
rect 4755 20012 5080 20040
rect 4755 20009 4767 20012
rect 4709 20003 4767 20009
rect 5074 20000 5080 20012
rect 5132 20000 5138 20052
rect 5810 20000 5816 20052
rect 5868 20040 5874 20052
rect 7098 20040 7104 20052
rect 5868 20012 7104 20040
rect 5868 20000 5874 20012
rect 7098 20000 7104 20012
rect 7156 20040 7162 20052
rect 7156 20012 8800 20040
rect 7156 20000 7162 20012
rect 5902 19972 5908 19984
rect 3988 19944 5908 19972
rect 3988 19845 4016 19944
rect 5902 19932 5908 19944
rect 5960 19932 5966 19984
rect 4614 19904 4620 19916
rect 4448 19876 4620 19904
rect 2593 19839 2651 19845
rect 2593 19805 2605 19839
rect 2639 19836 2651 19839
rect 2869 19839 2927 19845
rect 2869 19836 2881 19839
rect 2639 19808 2881 19836
rect 2639 19805 2651 19808
rect 2593 19799 2651 19805
rect 2869 19805 2881 19808
rect 2915 19805 2927 19839
rect 2869 19799 2927 19805
rect 3789 19839 3847 19845
rect 3789 19805 3801 19839
rect 3835 19805 3847 19839
rect 3789 19799 3847 19805
rect 3973 19839 4031 19845
rect 3973 19805 3985 19839
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 934 19728 940 19780
rect 992 19768 998 19780
rect 1581 19771 1639 19777
rect 1581 19768 1593 19771
rect 992 19740 1593 19768
rect 992 19728 998 19740
rect 1581 19737 1593 19740
rect 1627 19737 1639 19771
rect 1581 19731 1639 19737
rect 1394 19660 1400 19712
rect 1452 19700 1458 19712
rect 2608 19700 2636 19799
rect 3804 19768 3832 19799
rect 4062 19796 4068 19848
rect 4120 19796 4126 19848
rect 4154 19796 4160 19848
rect 4212 19836 4218 19848
rect 4448 19845 4476 19876
rect 4614 19864 4620 19876
rect 4672 19864 4678 19916
rect 6270 19904 6276 19916
rect 4724 19876 6276 19904
rect 4249 19839 4307 19845
rect 4249 19836 4261 19839
rect 4212 19808 4261 19836
rect 4212 19796 4218 19808
rect 4249 19805 4261 19808
rect 4295 19805 4307 19839
rect 4249 19799 4307 19805
rect 4433 19839 4491 19845
rect 4433 19805 4445 19839
rect 4479 19805 4491 19839
rect 4433 19799 4491 19805
rect 4522 19796 4528 19848
rect 4580 19796 4586 19848
rect 4724 19845 4752 19876
rect 6270 19864 6276 19876
rect 6328 19864 6334 19916
rect 7300 19913 7328 20012
rect 8772 19913 8800 20012
rect 10042 20000 10048 20052
rect 10100 20040 10106 20052
rect 11701 20043 11759 20049
rect 11701 20040 11713 20043
rect 10100 20012 11713 20040
rect 10100 20000 10106 20012
rect 11701 20009 11713 20012
rect 11747 20009 11759 20043
rect 11701 20003 11759 20009
rect 48314 20000 48320 20052
rect 48372 20000 48378 20052
rect 48498 20000 48504 20052
rect 48556 20040 48562 20052
rect 49697 20043 49755 20049
rect 49697 20040 49709 20043
rect 48556 20012 49709 20040
rect 48556 20000 48562 20012
rect 49697 20009 49709 20012
rect 49743 20009 49755 20043
rect 49697 20003 49755 20009
rect 51074 20000 51080 20052
rect 51132 20040 51138 20052
rect 51169 20043 51227 20049
rect 51169 20040 51181 20043
rect 51132 20012 51181 20040
rect 51132 20000 51138 20012
rect 51169 20009 51181 20012
rect 51215 20009 51227 20043
rect 51169 20003 51227 20009
rect 51258 20000 51264 20052
rect 51316 20000 51322 20052
rect 51810 20000 51816 20052
rect 51868 20000 51874 20052
rect 52362 20000 52368 20052
rect 52420 20040 52426 20052
rect 53101 20043 53159 20049
rect 53101 20040 53113 20043
rect 52420 20012 53113 20040
rect 52420 20000 52426 20012
rect 53101 20009 53113 20012
rect 53147 20040 53159 20043
rect 53147 20012 53696 20040
rect 53147 20009 53159 20012
rect 53101 20003 53159 20009
rect 7285 19907 7343 19913
rect 7285 19873 7297 19907
rect 7331 19873 7343 19907
rect 7285 19867 7343 19873
rect 8757 19907 8815 19913
rect 8757 19873 8769 19907
rect 8803 19873 8815 19907
rect 8757 19867 8815 19873
rect 47026 19864 47032 19916
rect 47084 19864 47090 19916
rect 47949 19907 48007 19913
rect 47949 19873 47961 19907
rect 47995 19904 48007 19907
rect 48332 19904 48360 20000
rect 50801 19975 50859 19981
rect 50801 19972 50813 19975
rect 49252 19944 50476 19972
rect 49252 19904 49280 19944
rect 49418 19904 49424 19916
rect 47995 19876 48360 19904
rect 48516 19876 49280 19904
rect 47995 19873 48007 19876
rect 47949 19867 48007 19873
rect 4709 19839 4767 19845
rect 4709 19805 4721 19839
rect 4755 19805 4767 19839
rect 4709 19799 4767 19805
rect 4801 19839 4859 19845
rect 4801 19805 4813 19839
rect 4847 19805 4859 19839
rect 4801 19799 4859 19805
rect 4985 19839 5043 19845
rect 4985 19805 4997 19839
rect 5031 19805 5043 19839
rect 4985 19799 5043 19805
rect 4080 19768 4108 19796
rect 4816 19768 4844 19799
rect 3804 19740 4844 19768
rect 5000 19768 5028 19799
rect 6730 19796 6736 19848
rect 6788 19836 6794 19848
rect 7018 19839 7076 19845
rect 7018 19836 7030 19839
rect 6788 19808 7030 19836
rect 6788 19796 6794 19808
rect 7018 19805 7030 19808
rect 7064 19805 7076 19839
rect 7018 19799 7076 19805
rect 7926 19796 7932 19848
rect 7984 19836 7990 19848
rect 8490 19839 8548 19845
rect 8490 19836 8502 19839
rect 7984 19808 8502 19836
rect 7984 19796 7990 19808
rect 8490 19805 8502 19808
rect 8536 19805 8548 19839
rect 8490 19799 8548 19805
rect 9306 19796 9312 19848
rect 9364 19836 9370 19848
rect 10137 19839 10195 19845
rect 10137 19836 10149 19839
rect 9364 19808 10149 19836
rect 9364 19796 9370 19808
rect 10137 19805 10149 19808
rect 10183 19805 10195 19839
rect 10137 19799 10195 19805
rect 11422 19796 11428 19848
rect 11480 19796 11486 19848
rect 11793 19839 11851 19845
rect 11793 19805 11805 19839
rect 11839 19805 11851 19839
rect 11793 19799 11851 19805
rect 8294 19768 8300 19780
rect 5000 19740 8300 19768
rect 1452 19672 2636 19700
rect 1452 19660 1458 19672
rect 3510 19660 3516 19712
rect 3568 19660 3574 19712
rect 3786 19660 3792 19712
rect 3844 19660 3850 19712
rect 4157 19703 4215 19709
rect 4157 19669 4169 19703
rect 4203 19700 4215 19703
rect 4614 19700 4620 19712
rect 4203 19672 4620 19700
rect 4203 19669 4215 19672
rect 4157 19663 4215 19669
rect 4614 19660 4620 19672
rect 4672 19660 4678 19712
rect 4706 19660 4712 19712
rect 4764 19700 4770 19712
rect 7392 19709 7420 19740
rect 8294 19728 8300 19740
rect 8352 19728 8358 19780
rect 10781 19771 10839 19777
rect 10781 19737 10793 19771
rect 10827 19768 10839 19771
rect 10962 19768 10968 19780
rect 10827 19740 10968 19768
rect 10827 19737 10839 19740
rect 10781 19731 10839 19737
rect 10962 19728 10968 19740
rect 11020 19728 11026 19780
rect 11808 19712 11836 19799
rect 41782 19796 41788 19848
rect 41840 19836 41846 19848
rect 48516 19836 48544 19876
rect 41840 19808 48544 19836
rect 41840 19796 41846 19808
rect 48590 19796 48596 19848
rect 48648 19796 48654 19848
rect 49252 19845 49280 19876
rect 49350 19876 49424 19904
rect 49350 19845 49378 19876
rect 49418 19864 49424 19876
rect 49476 19864 49482 19916
rect 50249 19907 50307 19913
rect 50249 19904 50261 19907
rect 49528 19876 50261 19904
rect 49528 19845 49556 19876
rect 50249 19873 50261 19876
rect 50295 19873 50307 19907
rect 50448 19904 50476 19944
rect 50632 19944 50813 19972
rect 50448 19876 50568 19904
rect 50249 19867 50307 19873
rect 49237 19839 49295 19845
rect 49237 19805 49249 19839
rect 49283 19805 49295 19839
rect 49237 19799 49295 19805
rect 49329 19839 49387 19845
rect 49329 19805 49341 19839
rect 49375 19805 49387 19839
rect 49329 19799 49387 19805
rect 49513 19839 49571 19845
rect 49513 19805 49525 19839
rect 49559 19805 49571 19839
rect 49513 19799 49571 19805
rect 49602 19796 49608 19848
rect 49660 19796 49666 19848
rect 49786 19796 49792 19848
rect 49844 19796 49850 19848
rect 50157 19839 50215 19845
rect 50157 19805 50169 19839
rect 50203 19805 50215 19839
rect 50157 19799 50215 19805
rect 46784 19771 46842 19777
rect 46784 19737 46796 19771
rect 46830 19768 46842 19771
rect 47305 19771 47363 19777
rect 47305 19768 47317 19771
rect 46830 19740 47317 19768
rect 46830 19737 46842 19740
rect 46784 19731 46842 19737
rect 47305 19737 47317 19740
rect 47351 19737 47363 19771
rect 47305 19731 47363 19737
rect 48961 19771 49019 19777
rect 48961 19737 48973 19771
rect 49007 19768 49019 19771
rect 49007 19740 49556 19768
rect 49007 19737 49019 19740
rect 48961 19731 49019 19737
rect 49528 19712 49556 19740
rect 4801 19703 4859 19709
rect 4801 19700 4813 19703
rect 4764 19672 4813 19700
rect 4764 19660 4770 19672
rect 4801 19669 4813 19672
rect 4847 19669 4859 19703
rect 4801 19663 4859 19669
rect 7377 19703 7435 19709
rect 7377 19669 7389 19703
rect 7423 19669 7435 19703
rect 7377 19663 7435 19669
rect 10870 19660 10876 19712
rect 10928 19660 10934 19712
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 12069 19703 12127 19709
rect 12069 19700 12081 19703
rect 11848 19672 12081 19700
rect 11848 19660 11854 19672
rect 12069 19669 12081 19672
rect 12115 19669 12127 19703
rect 12069 19663 12127 19669
rect 45649 19703 45707 19709
rect 45649 19669 45661 19703
rect 45695 19700 45707 19703
rect 45738 19700 45744 19712
rect 45695 19672 45744 19700
rect 45695 19669 45707 19672
rect 45649 19663 45707 19669
rect 45738 19660 45744 19672
rect 45796 19660 45802 19712
rect 47210 19660 47216 19712
rect 47268 19700 47274 19712
rect 48041 19703 48099 19709
rect 48041 19700 48053 19703
rect 47268 19672 48053 19700
rect 47268 19660 47274 19672
rect 48041 19669 48053 19672
rect 48087 19669 48099 19703
rect 48041 19663 48099 19669
rect 48406 19660 48412 19712
rect 48464 19700 48470 19712
rect 49421 19703 49479 19709
rect 49421 19700 49433 19703
rect 48464 19672 49433 19700
rect 48464 19660 48470 19672
rect 49421 19669 49433 19672
rect 49467 19669 49479 19703
rect 49421 19663 49479 19669
rect 49510 19660 49516 19712
rect 49568 19660 49574 19712
rect 50172 19700 50200 19799
rect 50338 19796 50344 19848
rect 50396 19796 50402 19848
rect 50430 19796 50436 19848
rect 50488 19796 50494 19848
rect 50540 19768 50568 19876
rect 50632 19845 50660 19944
rect 50801 19941 50813 19944
rect 50847 19941 50859 19975
rect 50801 19935 50859 19941
rect 50890 19932 50896 19984
rect 50948 19972 50954 19984
rect 51092 19972 51120 20000
rect 50948 19944 51120 19972
rect 50948 19932 50954 19944
rect 51092 19904 51120 19944
rect 50724 19876 51120 19904
rect 51276 19904 51304 20000
rect 53561 19975 53619 19981
rect 53561 19941 53573 19975
rect 53607 19941 53619 19975
rect 53561 19935 53619 19941
rect 53377 19907 53435 19913
rect 53377 19904 53389 19907
rect 51276 19876 52040 19904
rect 50724 19845 50752 19876
rect 50617 19839 50675 19845
rect 50617 19805 50629 19839
rect 50663 19805 50675 19839
rect 50617 19799 50675 19805
rect 50709 19839 50767 19845
rect 50709 19805 50721 19839
rect 50755 19805 50767 19839
rect 50709 19799 50767 19805
rect 50893 19839 50951 19845
rect 50893 19805 50905 19839
rect 50939 19836 50951 19839
rect 51350 19836 51356 19848
rect 50939 19808 51356 19836
rect 50939 19805 50951 19808
rect 50893 19799 50951 19805
rect 51350 19796 51356 19808
rect 51408 19796 51414 19848
rect 51721 19839 51779 19845
rect 51721 19805 51733 19839
rect 51767 19836 51779 19839
rect 51810 19836 51816 19848
rect 51767 19808 51816 19836
rect 51767 19805 51779 19808
rect 51721 19799 51779 19805
rect 51810 19796 51816 19808
rect 51868 19796 51874 19848
rect 52012 19845 52040 19876
rect 52196 19876 53389 19904
rect 52196 19845 52224 19876
rect 53377 19873 53389 19876
rect 53423 19873 53435 19907
rect 53576 19904 53604 19935
rect 53377 19867 53435 19873
rect 53484 19876 53604 19904
rect 53484 19845 53512 19876
rect 51905 19839 51963 19845
rect 51905 19805 51917 19839
rect 51951 19805 51963 19839
rect 51905 19799 51963 19805
rect 51997 19839 52055 19845
rect 51997 19805 52009 19839
rect 52043 19805 52055 19839
rect 51997 19799 52055 19805
rect 52181 19839 52239 19845
rect 52181 19805 52193 19839
rect 52227 19805 52239 19839
rect 52181 19799 52239 19805
rect 53285 19839 53343 19845
rect 53285 19805 53297 19839
rect 53331 19805 53343 19839
rect 53285 19799 53343 19805
rect 53469 19839 53527 19845
rect 53469 19805 53481 19839
rect 53515 19805 53527 19839
rect 53469 19799 53527 19805
rect 53561 19839 53619 19845
rect 53561 19805 53573 19839
rect 53607 19805 53619 19839
rect 53561 19799 53619 19805
rect 51920 19768 51948 19799
rect 52089 19771 52147 19777
rect 52089 19768 52101 19771
rect 50540 19740 50660 19768
rect 51920 19740 52101 19768
rect 50525 19703 50583 19709
rect 50525 19700 50537 19703
rect 50172 19672 50537 19700
rect 50525 19669 50537 19672
rect 50571 19669 50583 19703
rect 50632 19700 50660 19740
rect 52089 19737 52101 19740
rect 52135 19737 52147 19771
rect 53300 19768 53328 19799
rect 53300 19740 53512 19768
rect 52089 19731 52147 19737
rect 53484 19712 53512 19740
rect 51166 19700 51172 19712
rect 50632 19672 51172 19700
rect 50525 19663 50583 19669
rect 51166 19660 51172 19672
rect 51224 19700 51230 19712
rect 51626 19700 51632 19712
rect 51224 19672 51632 19700
rect 51224 19660 51230 19672
rect 51626 19660 51632 19672
rect 51684 19660 51690 19712
rect 53466 19660 53472 19712
rect 53524 19660 53530 19712
rect 53576 19700 53604 19799
rect 53668 19780 53696 20012
rect 55214 20000 55220 20052
rect 55272 20040 55278 20052
rect 55272 20012 56272 20040
rect 55272 20000 55278 20012
rect 56244 19972 56272 20012
rect 56686 20000 56692 20052
rect 56744 20000 56750 20052
rect 58161 20043 58219 20049
rect 56796 20012 57744 20040
rect 56796 19972 56824 20012
rect 56244 19944 56824 19972
rect 57716 19972 57744 20012
rect 58161 20009 58173 20043
rect 58207 20040 58219 20043
rect 58912 20040 58940 20352
rect 58207 20012 58940 20040
rect 58207 20009 58219 20012
rect 58161 20003 58219 20009
rect 58345 19975 58403 19981
rect 58345 19972 58357 19975
rect 57716 19944 58357 19972
rect 58345 19941 58357 19944
rect 58391 19941 58403 19975
rect 58345 19935 58403 19941
rect 55033 19907 55091 19913
rect 55033 19904 55045 19907
rect 53944 19876 55045 19904
rect 53944 19836 53972 19876
rect 55033 19873 55045 19876
rect 55079 19873 55091 19907
rect 55033 19867 55091 19873
rect 53760 19808 53972 19836
rect 53650 19728 53656 19780
rect 53708 19728 53714 19780
rect 53760 19700 53788 19808
rect 54018 19796 54024 19848
rect 54076 19796 54082 19848
rect 54113 19839 54171 19845
rect 54113 19805 54125 19839
rect 54159 19836 54171 19839
rect 54202 19836 54208 19848
rect 54159 19808 54208 19836
rect 54159 19805 54171 19808
rect 54113 19799 54171 19805
rect 54202 19796 54208 19808
rect 54260 19796 54266 19848
rect 54294 19796 54300 19848
rect 54352 19796 54358 19848
rect 54941 19839 54999 19845
rect 54941 19805 54953 19839
rect 54987 19836 54999 19839
rect 55125 19839 55183 19845
rect 54987 19808 55076 19836
rect 54987 19805 54999 19808
rect 54941 19799 54999 19805
rect 55048 19780 55076 19808
rect 55125 19805 55137 19839
rect 55171 19805 55183 19839
rect 55125 19799 55183 19805
rect 53837 19771 53895 19777
rect 53837 19737 53849 19771
rect 53883 19768 53895 19771
rect 53883 19740 54064 19768
rect 53883 19737 53895 19740
rect 53837 19731 53895 19737
rect 54036 19709 54064 19740
rect 55030 19728 55036 19780
rect 55088 19728 55094 19780
rect 53576 19672 53788 19700
rect 54021 19703 54079 19709
rect 54021 19669 54033 19703
rect 54067 19669 54079 19703
rect 55140 19700 55168 19799
rect 55306 19796 55312 19848
rect 55364 19836 55370 19848
rect 56410 19836 56416 19848
rect 55364 19808 56416 19836
rect 55364 19796 55370 19808
rect 56410 19796 56416 19808
rect 56468 19836 56474 19848
rect 56781 19839 56839 19845
rect 56781 19836 56793 19839
rect 56468 19808 56793 19836
rect 56468 19796 56474 19808
rect 56781 19805 56793 19808
rect 56827 19805 56839 19839
rect 56781 19799 56839 19805
rect 58250 19796 58256 19848
rect 58308 19796 58314 19848
rect 55214 19728 55220 19780
rect 55272 19768 55278 19780
rect 57054 19777 57060 19780
rect 55554 19771 55612 19777
rect 55554 19768 55566 19771
rect 55272 19740 55566 19768
rect 55272 19728 55278 19740
rect 55554 19737 55566 19740
rect 55600 19737 55612 19771
rect 55554 19731 55612 19737
rect 57048 19731 57060 19777
rect 57054 19728 57060 19731
rect 57112 19728 57118 19780
rect 55674 19700 55680 19712
rect 55140 19672 55680 19700
rect 54021 19663 54079 19669
rect 55674 19660 55680 19672
rect 55732 19660 55738 19712
rect 56318 19660 56324 19712
rect 56376 19700 56382 19712
rect 57330 19700 57336 19712
rect 56376 19672 57336 19700
rect 56376 19660 56382 19672
rect 57330 19660 57336 19672
rect 57388 19660 57394 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 1394 19456 1400 19508
rect 1452 19456 1458 19508
rect 8846 19456 8852 19508
rect 8904 19456 8910 19508
rect 9125 19499 9183 19505
rect 9125 19465 9137 19499
rect 9171 19496 9183 19499
rect 10870 19496 10876 19508
rect 9171 19468 9352 19496
rect 9171 19465 9183 19468
rect 9125 19459 9183 19465
rect 2406 19388 2412 19440
rect 2464 19428 2470 19440
rect 5350 19428 5356 19440
rect 2464 19400 5356 19428
rect 2464 19388 2470 19400
rect 5350 19388 5356 19400
rect 5408 19388 5414 19440
rect 9324 19372 9352 19468
rect 10612 19468 10876 19496
rect 10318 19428 10324 19440
rect 10166 19400 10324 19428
rect 10318 19388 10324 19400
rect 10376 19388 10382 19440
rect 10612 19437 10640 19468
rect 10870 19456 10876 19468
rect 10928 19456 10934 19508
rect 11793 19499 11851 19505
rect 11793 19465 11805 19499
rect 11839 19496 11851 19499
rect 11974 19496 11980 19508
rect 11839 19468 11980 19496
rect 11839 19465 11851 19468
rect 11793 19459 11851 19465
rect 10597 19431 10655 19437
rect 10597 19397 10609 19431
rect 10643 19397 10655 19431
rect 11808 19428 11836 19459
rect 11974 19456 11980 19468
rect 12032 19456 12038 19508
rect 47210 19456 47216 19508
rect 47268 19456 47274 19508
rect 47946 19496 47952 19508
rect 47412 19468 47952 19496
rect 10597 19391 10655 19397
rect 10888 19400 11836 19428
rect 3142 19320 3148 19372
rect 3200 19320 3206 19372
rect 3510 19320 3516 19372
rect 3568 19360 3574 19372
rect 3973 19363 4031 19369
rect 3973 19360 3985 19363
rect 3568 19332 3985 19360
rect 3568 19320 3574 19332
rect 3973 19329 3985 19332
rect 4019 19329 4031 19363
rect 3973 19323 4031 19329
rect 4157 19363 4215 19369
rect 4157 19329 4169 19363
rect 4203 19329 4215 19363
rect 4157 19323 4215 19329
rect 8941 19363 8999 19369
rect 8941 19329 8953 19363
rect 8987 19329 8999 19363
rect 8941 19323 8999 19329
rect 2866 19252 2872 19304
rect 2924 19252 2930 19304
rect 3881 19295 3939 19301
rect 3881 19261 3893 19295
rect 3927 19292 3939 19295
rect 4065 19295 4123 19301
rect 4065 19292 4077 19295
rect 3927 19264 4077 19292
rect 3927 19261 3939 19264
rect 3881 19255 3939 19261
rect 4065 19261 4077 19264
rect 4111 19261 4123 19295
rect 4065 19255 4123 19261
rect 4172 19224 4200 19323
rect 6822 19252 6828 19304
rect 6880 19292 6886 19304
rect 7653 19295 7711 19301
rect 7653 19292 7665 19295
rect 6880 19264 7665 19292
rect 6880 19252 6886 19264
rect 7653 19261 7665 19264
rect 7699 19261 7711 19295
rect 7653 19255 7711 19261
rect 8665 19295 8723 19301
rect 8665 19261 8677 19295
rect 8711 19292 8723 19295
rect 8956 19292 8984 19323
rect 9306 19320 9312 19372
rect 9364 19320 9370 19372
rect 10888 19369 10916 19400
rect 10873 19363 10931 19369
rect 10873 19329 10885 19363
rect 10919 19329 10931 19363
rect 10873 19323 10931 19329
rect 10962 19320 10968 19372
rect 11020 19320 11026 19372
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19360 11207 19363
rect 11238 19360 11244 19372
rect 11195 19332 11244 19360
rect 11195 19329 11207 19332
rect 11149 19323 11207 19329
rect 11238 19320 11244 19332
rect 11296 19320 11302 19372
rect 47228 19369 47256 19456
rect 47412 19369 47440 19468
rect 47946 19456 47952 19468
rect 48004 19456 48010 19508
rect 49142 19456 49148 19508
rect 49200 19456 49206 19508
rect 49326 19456 49332 19508
rect 49384 19456 49390 19508
rect 50433 19499 50491 19505
rect 50433 19465 50445 19499
rect 50479 19496 50491 19499
rect 50614 19496 50620 19508
rect 50479 19468 50620 19496
rect 50479 19465 50491 19468
rect 50433 19459 50491 19465
rect 50614 19456 50620 19468
rect 50672 19456 50678 19508
rect 51350 19456 51356 19508
rect 51408 19496 51414 19508
rect 51721 19499 51779 19505
rect 51721 19496 51733 19499
rect 51408 19468 51733 19496
rect 51408 19456 51414 19468
rect 51721 19465 51733 19468
rect 51767 19465 51779 19499
rect 51721 19459 51779 19465
rect 53650 19456 53656 19508
rect 53708 19456 53714 19508
rect 55033 19499 55091 19505
rect 55033 19465 55045 19499
rect 55079 19496 55091 19499
rect 55214 19496 55220 19508
rect 55079 19468 55220 19496
rect 55079 19465 55091 19468
rect 55033 19459 55091 19465
rect 55214 19456 55220 19468
rect 55272 19456 55278 19508
rect 56965 19499 57023 19505
rect 56965 19465 56977 19499
rect 57011 19496 57023 19499
rect 57054 19496 57060 19508
rect 57011 19468 57060 19496
rect 57011 19465 57023 19468
rect 56965 19459 57023 19465
rect 57054 19456 57060 19468
rect 57112 19456 57118 19508
rect 57425 19499 57483 19505
rect 57425 19465 57437 19499
rect 57471 19496 57483 19499
rect 57471 19468 57560 19496
rect 57471 19465 57483 19468
rect 57425 19459 57483 19465
rect 49160 19369 49188 19456
rect 53668 19428 53696 19456
rect 56594 19428 56600 19440
rect 49252 19400 49464 19428
rect 47213 19363 47271 19369
rect 47213 19329 47225 19363
rect 47259 19329 47271 19363
rect 47213 19323 47271 19329
rect 47397 19363 47455 19369
rect 47397 19329 47409 19363
rect 47443 19329 47455 19363
rect 49145 19363 49203 19369
rect 47397 19323 47455 19329
rect 47504 19332 48912 19360
rect 42610 19292 42616 19304
rect 8711 19264 42616 19292
rect 8711 19261 8723 19264
rect 8665 19255 8723 19261
rect 42610 19252 42616 19264
rect 42668 19252 42674 19304
rect 47305 19295 47363 19301
rect 47305 19261 47317 19295
rect 47351 19292 47363 19295
rect 47504 19292 47532 19332
rect 48884 19301 48912 19332
rect 49145 19329 49157 19363
rect 49191 19329 49203 19363
rect 49145 19323 49203 19329
rect 47351 19264 47532 19292
rect 48133 19295 48191 19301
rect 47351 19261 47363 19264
rect 47305 19255 47363 19261
rect 48133 19261 48145 19295
rect 48179 19261 48191 19295
rect 48133 19255 48191 19261
rect 48869 19295 48927 19301
rect 48869 19261 48881 19295
rect 48915 19261 48927 19295
rect 48869 19255 48927 19261
rect 4080 19196 4200 19224
rect 4080 19168 4108 19196
rect 47210 19184 47216 19236
rect 47268 19224 47274 19236
rect 48148 19224 48176 19255
rect 49050 19252 49056 19304
rect 49108 19292 49114 19304
rect 49252 19292 49280 19400
rect 49436 19369 49464 19400
rect 49620 19400 50568 19428
rect 53668 19400 56600 19428
rect 49620 19369 49648 19400
rect 49329 19363 49387 19369
rect 49329 19329 49341 19363
rect 49375 19329 49387 19363
rect 49329 19323 49387 19329
rect 49421 19363 49479 19369
rect 49421 19329 49433 19363
rect 49467 19329 49479 19363
rect 49421 19323 49479 19329
rect 49605 19363 49663 19369
rect 49605 19329 49617 19363
rect 49651 19329 49663 19363
rect 49605 19323 49663 19329
rect 49108 19264 49280 19292
rect 49108 19252 49114 19264
rect 47268 19196 48176 19224
rect 49344 19224 49372 19323
rect 49694 19320 49700 19372
rect 49752 19320 49758 19372
rect 49878 19320 49884 19372
rect 49936 19320 49942 19372
rect 50154 19320 50160 19372
rect 50212 19360 50218 19372
rect 50540 19369 50568 19400
rect 56594 19388 56600 19400
rect 56652 19388 56658 19440
rect 57532 19428 57560 19468
rect 57606 19456 57612 19508
rect 57664 19496 57670 19508
rect 58342 19496 58348 19508
rect 57664 19468 58348 19496
rect 57664 19456 57670 19468
rect 58342 19456 58348 19468
rect 58400 19456 58406 19508
rect 57532 19400 58480 19428
rect 50341 19363 50399 19369
rect 50341 19360 50353 19363
rect 50212 19332 50353 19360
rect 50212 19320 50218 19332
rect 50341 19329 50353 19332
rect 50387 19329 50399 19363
rect 50341 19323 50399 19329
rect 50525 19363 50583 19369
rect 50525 19329 50537 19363
rect 50571 19360 50583 19363
rect 50982 19360 50988 19372
rect 50571 19332 50988 19360
rect 50571 19329 50583 19332
rect 50525 19323 50583 19329
rect 50982 19320 50988 19332
rect 51040 19320 51046 19372
rect 51353 19363 51411 19369
rect 51353 19360 51365 19363
rect 51184 19332 51365 19360
rect 51184 19304 51212 19332
rect 51353 19329 51365 19332
rect 51399 19360 51411 19363
rect 51399 19332 51580 19360
rect 51399 19329 51411 19332
rect 51353 19323 51411 19329
rect 49513 19295 49571 19301
rect 49513 19261 49525 19295
rect 49559 19292 49571 19295
rect 49786 19292 49792 19304
rect 49559 19264 49792 19292
rect 49559 19261 49571 19264
rect 49513 19255 49571 19261
rect 49786 19252 49792 19264
rect 49844 19252 49850 19304
rect 50249 19295 50307 19301
rect 50249 19261 50261 19295
rect 50295 19292 50307 19295
rect 50890 19292 50896 19304
rect 50295 19264 50896 19292
rect 50295 19261 50307 19264
rect 50249 19255 50307 19261
rect 50890 19252 50896 19264
rect 50948 19252 50954 19304
rect 51166 19252 51172 19304
rect 51224 19252 51230 19304
rect 51552 19292 51580 19332
rect 51626 19320 51632 19372
rect 51684 19320 51690 19372
rect 51718 19320 51724 19372
rect 51776 19320 51782 19372
rect 51902 19320 51908 19372
rect 51960 19320 51966 19372
rect 52012 19332 53604 19360
rect 52012 19292 52040 19332
rect 51552 19264 52040 19292
rect 53576 19292 53604 19332
rect 53650 19320 53656 19372
rect 53708 19360 53714 19372
rect 54202 19360 54208 19372
rect 53708 19332 54208 19360
rect 53708 19320 53714 19332
rect 54202 19320 54208 19332
rect 54260 19320 54266 19372
rect 54757 19363 54815 19369
rect 54757 19329 54769 19363
rect 54803 19360 54815 19363
rect 55401 19363 55459 19369
rect 55401 19360 55413 19363
rect 54803 19332 55413 19360
rect 54803 19329 54815 19332
rect 54757 19323 54815 19329
rect 55401 19329 55413 19332
rect 55447 19329 55459 19363
rect 55401 19323 55459 19329
rect 55493 19363 55551 19369
rect 55493 19329 55505 19363
rect 55539 19360 55551 19363
rect 55674 19360 55680 19372
rect 55539 19332 55680 19360
rect 55539 19329 55551 19332
rect 55493 19323 55551 19329
rect 55674 19320 55680 19332
rect 55732 19360 55738 19372
rect 56134 19360 56140 19372
rect 55732 19332 56140 19360
rect 55732 19320 55738 19332
rect 56134 19320 56140 19332
rect 56192 19320 56198 19372
rect 57241 19363 57299 19369
rect 57241 19329 57253 19363
rect 57287 19329 57299 19363
rect 57241 19323 57299 19329
rect 53834 19292 53840 19304
rect 53576 19264 53840 19292
rect 53834 19252 53840 19264
rect 53892 19252 53898 19304
rect 55033 19295 55091 19301
rect 55033 19261 55045 19295
rect 55079 19292 55091 19295
rect 55122 19292 55128 19304
rect 55079 19264 55128 19292
rect 55079 19261 55091 19264
rect 55033 19255 55091 19261
rect 55122 19252 55128 19264
rect 55180 19252 55186 19304
rect 56965 19295 57023 19301
rect 56965 19261 56977 19295
rect 57011 19292 57023 19295
rect 57054 19292 57060 19304
rect 57011 19264 57060 19292
rect 57011 19261 57023 19264
rect 56965 19255 57023 19261
rect 57054 19252 57060 19264
rect 57112 19252 57118 19304
rect 57149 19227 57207 19233
rect 57149 19224 57161 19227
rect 49344 19196 49832 19224
rect 47268 19184 47274 19196
rect 3234 19116 3240 19168
rect 3292 19116 3298 19168
rect 4062 19116 4068 19168
rect 4120 19116 4126 19168
rect 8297 19159 8355 19165
rect 8297 19125 8309 19159
rect 8343 19156 8355 19159
rect 8386 19156 8392 19168
rect 8343 19128 8392 19156
rect 8343 19125 8355 19128
rect 8297 19119 8355 19125
rect 8386 19116 8392 19128
rect 8444 19116 8450 19168
rect 11054 19116 11060 19168
rect 11112 19116 11118 19168
rect 47394 19116 47400 19168
rect 47452 19156 47458 19168
rect 47581 19159 47639 19165
rect 47581 19156 47593 19159
rect 47452 19128 47593 19156
rect 47452 19116 47458 19128
rect 47581 19125 47593 19128
rect 47627 19125 47639 19159
rect 47581 19119 47639 19125
rect 48314 19116 48320 19168
rect 48372 19116 48378 19168
rect 49804 19165 49832 19196
rect 54864 19196 57161 19224
rect 54864 19168 54892 19196
rect 57149 19193 57161 19196
rect 57195 19193 57207 19227
rect 57256 19224 57284 19323
rect 57330 19320 57336 19372
rect 57388 19320 57394 19372
rect 57517 19363 57575 19369
rect 57517 19329 57529 19363
rect 57563 19360 57575 19363
rect 57790 19360 57796 19372
rect 57563 19332 57796 19360
rect 57563 19329 57575 19332
rect 57517 19323 57575 19329
rect 57790 19320 57796 19332
rect 57848 19320 57854 19372
rect 57422 19252 57428 19304
rect 57480 19292 57486 19304
rect 58452 19301 58480 19400
rect 57885 19295 57943 19301
rect 57885 19292 57897 19295
rect 57480 19264 57897 19292
rect 57480 19252 57486 19264
rect 57885 19261 57897 19264
rect 57931 19261 57943 19295
rect 57885 19255 57943 19261
rect 58437 19295 58495 19301
rect 58437 19261 58449 19295
rect 58483 19261 58495 19295
rect 58437 19255 58495 19261
rect 57606 19224 57612 19236
rect 57256 19196 57612 19224
rect 57149 19187 57207 19193
rect 57606 19184 57612 19196
rect 57664 19184 57670 19236
rect 49789 19159 49847 19165
rect 49789 19125 49801 19159
rect 49835 19125 49847 19159
rect 49789 19119 49847 19125
rect 52270 19116 52276 19168
rect 52328 19156 52334 19168
rect 54846 19156 54852 19168
rect 52328 19128 54852 19156
rect 52328 19116 52334 19128
rect 54846 19116 54852 19128
rect 54904 19116 54910 19168
rect 55030 19116 55036 19168
rect 55088 19156 55094 19168
rect 57330 19156 57336 19168
rect 55088 19128 57336 19156
rect 55088 19116 55094 19128
rect 57330 19116 57336 19128
rect 57388 19116 57394 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 2148 18924 2774 18952
rect 2148 18757 2176 18924
rect 2746 18884 2774 18924
rect 2866 18912 2872 18964
rect 2924 18952 2930 18964
rect 3329 18955 3387 18961
rect 3329 18952 3341 18955
rect 2924 18924 3341 18952
rect 2924 18912 2930 18924
rect 3329 18921 3341 18924
rect 3375 18921 3387 18955
rect 3329 18915 3387 18921
rect 3786 18912 3792 18964
rect 3844 18912 3850 18964
rect 4617 18955 4675 18961
rect 4617 18921 4629 18955
rect 4663 18952 4675 18955
rect 4798 18952 4804 18964
rect 4663 18924 4804 18952
rect 4663 18921 4675 18924
rect 4617 18915 4675 18921
rect 4798 18912 4804 18924
rect 4856 18952 4862 18964
rect 6733 18955 6791 18961
rect 4856 18924 6684 18952
rect 4856 18912 4862 18924
rect 3804 18884 3832 18912
rect 2746 18856 3832 18884
rect 4706 18844 4712 18896
rect 4764 18844 4770 18896
rect 2409 18819 2467 18825
rect 2409 18785 2421 18819
rect 2455 18816 2467 18819
rect 3234 18816 3240 18828
rect 2455 18788 3240 18816
rect 2455 18785 2467 18788
rect 2409 18779 2467 18785
rect 3234 18776 3240 18788
rect 3292 18776 3298 18828
rect 3513 18819 3571 18825
rect 3513 18785 3525 18819
rect 3559 18816 3571 18819
rect 4341 18819 4399 18825
rect 4341 18816 4353 18819
rect 3559 18788 4353 18816
rect 3559 18785 3571 18788
rect 3513 18779 3571 18785
rect 4341 18785 4353 18788
rect 4387 18785 4399 18819
rect 4341 18779 4399 18785
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18717 2191 18751
rect 2133 18711 2191 18717
rect 2222 18708 2228 18760
rect 2280 18708 2286 18760
rect 2685 18751 2743 18757
rect 2685 18748 2697 18751
rect 2424 18720 2697 18748
rect 2424 18689 2452 18720
rect 2685 18717 2697 18720
rect 2731 18717 2743 18751
rect 2685 18711 2743 18717
rect 3421 18751 3479 18757
rect 3421 18717 3433 18751
rect 3467 18717 3479 18751
rect 3421 18711 3479 18717
rect 2409 18683 2467 18689
rect 2409 18649 2421 18683
rect 2455 18649 2467 18683
rect 3436 18680 3464 18711
rect 3602 18708 3608 18760
rect 3660 18708 3666 18760
rect 4062 18708 4068 18760
rect 4120 18708 4126 18760
rect 4525 18751 4583 18757
rect 4525 18717 4537 18751
rect 4571 18748 4583 18751
rect 4724 18748 4752 18844
rect 4801 18819 4859 18825
rect 4801 18785 4813 18819
rect 4847 18816 4859 18819
rect 4890 18816 4896 18828
rect 4847 18788 4896 18816
rect 4847 18785 4859 18788
rect 4801 18779 4859 18785
rect 4890 18776 4896 18788
rect 4948 18776 4954 18828
rect 6656 18760 6684 18924
rect 6733 18921 6745 18955
rect 6779 18952 6791 18955
rect 6822 18952 6828 18964
rect 6779 18924 6828 18952
rect 6779 18921 6791 18924
rect 6733 18915 6791 18921
rect 6822 18912 6828 18924
rect 6880 18912 6886 18964
rect 9769 18955 9827 18961
rect 9769 18921 9781 18955
rect 9815 18952 9827 18955
rect 11422 18952 11428 18964
rect 9815 18924 11428 18952
rect 9815 18921 9827 18924
rect 9769 18915 9827 18921
rect 11422 18912 11428 18924
rect 11480 18912 11486 18964
rect 49878 18912 49884 18964
rect 49936 18952 49942 18964
rect 50157 18955 50215 18961
rect 50157 18952 50169 18955
rect 49936 18924 50169 18952
rect 49936 18912 49942 18924
rect 50157 18921 50169 18924
rect 50203 18921 50215 18955
rect 50157 18915 50215 18921
rect 51718 18912 51724 18964
rect 51776 18912 51782 18964
rect 51902 18912 51908 18964
rect 51960 18952 51966 18964
rect 51960 18924 57192 18952
rect 51960 18912 51966 18924
rect 9677 18887 9735 18893
rect 9677 18853 9689 18887
rect 9723 18884 9735 18887
rect 9950 18884 9956 18896
rect 9723 18856 9956 18884
rect 9723 18853 9735 18856
rect 9677 18847 9735 18853
rect 9950 18844 9956 18856
rect 10008 18844 10014 18896
rect 48961 18887 49019 18893
rect 47044 18856 47624 18884
rect 47044 18828 47072 18856
rect 6822 18776 6828 18828
rect 6880 18776 6886 18828
rect 8386 18776 8392 18828
rect 8444 18816 8450 18828
rect 8481 18819 8539 18825
rect 8481 18816 8493 18819
rect 8444 18788 8493 18816
rect 8444 18776 8450 18788
rect 8481 18785 8493 18788
rect 8527 18785 8539 18819
rect 8481 18779 8539 18785
rect 8757 18819 8815 18825
rect 8757 18785 8769 18819
rect 8803 18816 8815 18819
rect 9766 18816 9772 18828
rect 8803 18788 9772 18816
rect 8803 18785 8815 18788
rect 8757 18779 8815 18785
rect 9766 18776 9772 18788
rect 9824 18776 9830 18828
rect 9861 18819 9919 18825
rect 9861 18785 9873 18819
rect 9907 18816 9919 18819
rect 10505 18819 10563 18825
rect 10505 18816 10517 18819
rect 9907 18788 10517 18816
rect 9907 18785 9919 18788
rect 9861 18779 9919 18785
rect 10505 18785 10517 18788
rect 10551 18785 10563 18819
rect 10505 18779 10563 18785
rect 11054 18776 11060 18828
rect 11112 18776 11118 18828
rect 47026 18776 47032 18828
rect 47084 18776 47090 18828
rect 47596 18825 47624 18856
rect 48961 18853 48973 18887
rect 49007 18884 49019 18887
rect 49007 18856 49372 18884
rect 49007 18853 49019 18856
rect 48961 18847 49019 18853
rect 47581 18819 47639 18825
rect 47320 18788 47532 18816
rect 5261 18751 5319 18757
rect 5261 18748 5273 18751
rect 4571 18720 4752 18748
rect 4816 18720 5273 18748
rect 4571 18717 4583 18720
rect 4525 18711 4583 18717
rect 4080 18680 4108 18708
rect 4816 18689 4844 18720
rect 5261 18717 5273 18720
rect 5307 18717 5319 18751
rect 5261 18711 5319 18717
rect 6362 18708 6368 18760
rect 6420 18748 6426 18760
rect 6549 18751 6607 18757
rect 6549 18748 6561 18751
rect 6420 18720 6561 18748
rect 6420 18708 6426 18720
rect 6549 18717 6561 18720
rect 6595 18717 6607 18751
rect 6549 18711 6607 18717
rect 6638 18708 6644 18760
rect 6696 18708 6702 18760
rect 47320 18757 47348 18788
rect 9585 18751 9643 18757
rect 9585 18717 9597 18751
rect 9631 18717 9643 18751
rect 9585 18711 9643 18717
rect 47121 18751 47179 18757
rect 47121 18717 47133 18751
rect 47167 18717 47179 18751
rect 47121 18711 47179 18717
rect 47305 18751 47363 18757
rect 47305 18717 47317 18751
rect 47351 18717 47363 18751
rect 47305 18711 47363 18717
rect 3436 18652 4108 18680
rect 4801 18683 4859 18689
rect 2409 18643 2467 18649
rect 4801 18649 4813 18683
rect 4847 18649 4859 18683
rect 9600 18680 9628 18711
rect 12066 18680 12072 18692
rect 4801 18643 4859 18649
rect 5828 18652 7052 18680
rect 8050 18652 8156 18680
rect 9600 18652 12072 18680
rect 3786 18572 3792 18624
rect 3844 18572 3850 18624
rect 4522 18572 4528 18624
rect 4580 18612 4586 18624
rect 5828 18612 5856 18652
rect 7024 18624 7052 18652
rect 4580 18584 5856 18612
rect 4580 18572 4586 18584
rect 5902 18572 5908 18624
rect 5960 18572 5966 18624
rect 7006 18572 7012 18624
rect 7064 18572 7070 18624
rect 8128 18612 8156 18652
rect 12066 18640 12072 18652
rect 12124 18640 12130 18692
rect 46784 18683 46842 18689
rect 46784 18649 46796 18683
rect 46830 18680 46842 18683
rect 46934 18680 46940 18692
rect 46830 18652 46940 18680
rect 46830 18649 46842 18652
rect 46784 18643 46842 18649
rect 46934 18640 46940 18652
rect 46992 18640 46998 18692
rect 47136 18680 47164 18711
rect 47394 18708 47400 18760
rect 47452 18708 47458 18760
rect 47412 18680 47440 18708
rect 47136 18652 47440 18680
rect 47504 18680 47532 18788
rect 47581 18785 47593 18819
rect 47627 18785 47639 18819
rect 47581 18779 47639 18785
rect 47848 18751 47906 18757
rect 47848 18717 47860 18751
rect 47894 18748 47906 18751
rect 48314 18748 48320 18760
rect 47894 18720 48320 18748
rect 47894 18717 47906 18720
rect 47848 18711 47906 18717
rect 48314 18708 48320 18720
rect 48372 18708 48378 18760
rect 48406 18708 48412 18760
rect 48464 18708 48470 18760
rect 49344 18748 49372 18856
rect 49436 18856 50936 18884
rect 49436 18828 49464 18856
rect 49418 18776 49424 18828
rect 49476 18776 49482 18828
rect 49510 18776 49516 18828
rect 49568 18816 49574 18828
rect 50908 18816 50936 18856
rect 50982 18844 50988 18896
rect 51040 18884 51046 18896
rect 51040 18856 52592 18884
rect 51040 18844 51046 18856
rect 52270 18816 52276 18828
rect 49568 18788 50200 18816
rect 50908 18788 52276 18816
rect 49568 18776 49574 18788
rect 49786 18748 49792 18760
rect 49344 18720 49792 18748
rect 49786 18708 49792 18720
rect 49844 18708 49850 18760
rect 50172 18757 50200 18788
rect 52270 18776 52276 18788
rect 52328 18776 52334 18828
rect 52564 18825 52592 18856
rect 53834 18844 53840 18896
rect 53892 18884 53898 18896
rect 53892 18856 54984 18884
rect 53892 18844 53898 18856
rect 52457 18819 52515 18825
rect 52457 18785 52469 18819
rect 52503 18785 52515 18819
rect 52457 18779 52515 18785
rect 52549 18819 52607 18825
rect 52549 18785 52561 18819
rect 52595 18785 52607 18819
rect 52549 18779 52607 18785
rect 54665 18819 54723 18825
rect 54665 18785 54677 18819
rect 54711 18816 54723 18819
rect 54849 18819 54907 18825
rect 54849 18816 54861 18819
rect 54711 18788 54861 18816
rect 54711 18785 54723 18788
rect 54665 18779 54723 18785
rect 54849 18785 54861 18788
rect 54895 18785 54907 18819
rect 54849 18779 54907 18785
rect 50157 18751 50215 18757
rect 50157 18717 50169 18751
rect 50203 18717 50215 18751
rect 50157 18711 50215 18717
rect 50341 18751 50399 18757
rect 50341 18717 50353 18751
rect 50387 18717 50399 18751
rect 50341 18711 50399 18717
rect 50433 18751 50491 18757
rect 50433 18717 50445 18751
rect 50479 18717 50491 18751
rect 50433 18711 50491 18717
rect 48424 18680 48452 18708
rect 47504 18652 48452 18680
rect 49326 18640 49332 18692
rect 49384 18680 49390 18692
rect 50356 18680 50384 18711
rect 49384 18652 50384 18680
rect 50448 18680 50476 18711
rect 50614 18708 50620 18760
rect 50672 18708 50678 18760
rect 51258 18708 51264 18760
rect 51316 18708 51322 18760
rect 51537 18751 51595 18757
rect 51537 18717 51549 18751
rect 51583 18748 51595 18751
rect 51626 18748 51632 18760
rect 51583 18720 51632 18748
rect 51583 18717 51595 18720
rect 51537 18711 51595 18717
rect 51626 18708 51632 18720
rect 51684 18708 51690 18760
rect 51718 18708 51724 18760
rect 51776 18708 51782 18760
rect 52181 18751 52239 18757
rect 52181 18717 52193 18751
rect 52227 18717 52239 18751
rect 52472 18748 52500 18779
rect 52181 18711 52239 18717
rect 52380 18720 52500 18748
rect 51276 18680 51304 18708
rect 50448 18652 51304 18680
rect 49384 18640 49390 18652
rect 8294 18612 8300 18624
rect 8128 18584 8300 18612
rect 8294 18572 8300 18584
rect 8352 18612 8358 18624
rect 10318 18612 10324 18624
rect 8352 18584 10324 18612
rect 8352 18572 8358 18584
rect 10318 18572 10324 18584
rect 10376 18572 10382 18624
rect 45646 18572 45652 18624
rect 45704 18572 45710 18624
rect 47302 18572 47308 18624
rect 47360 18572 47366 18624
rect 49142 18572 49148 18624
rect 49200 18572 49206 18624
rect 49878 18572 49884 18624
rect 49936 18612 49942 18624
rect 50525 18615 50583 18621
rect 50525 18612 50537 18615
rect 49936 18584 50537 18612
rect 49936 18572 49942 18584
rect 50525 18581 50537 18584
rect 50571 18581 50583 18615
rect 51276 18612 51304 18652
rect 51534 18612 51540 18624
rect 51276 18584 51540 18612
rect 50525 18575 50583 18581
rect 51534 18572 51540 18584
rect 51592 18572 51598 18624
rect 52196 18612 52224 18711
rect 52270 18612 52276 18624
rect 52196 18584 52276 18612
rect 52270 18572 52276 18584
rect 52328 18572 52334 18624
rect 52380 18612 52408 18720
rect 54754 18708 54760 18760
rect 54812 18708 54818 18760
rect 54956 18757 54984 18856
rect 56778 18844 56784 18896
rect 56836 18884 56842 18896
rect 57057 18887 57115 18893
rect 57057 18884 57069 18887
rect 56836 18856 57069 18884
rect 56836 18844 56842 18856
rect 57057 18853 57069 18856
rect 57103 18853 57115 18887
rect 57164 18884 57192 18924
rect 57606 18912 57612 18964
rect 57664 18912 57670 18964
rect 58342 18912 58348 18964
rect 58400 18912 58406 18964
rect 58158 18884 58164 18896
rect 57164 18856 58164 18884
rect 57057 18847 57115 18853
rect 54941 18751 54999 18757
rect 54941 18717 54953 18751
rect 54987 18748 54999 18751
rect 55398 18748 55404 18760
rect 54987 18720 55404 18748
rect 54987 18717 54999 18720
rect 54941 18711 54999 18717
rect 55398 18708 55404 18720
rect 55456 18748 55462 18760
rect 56318 18748 56324 18760
rect 55456 18720 56324 18748
rect 55456 18708 55462 18720
rect 56318 18708 56324 18720
rect 56376 18708 56382 18760
rect 52457 18683 52515 18689
rect 52457 18649 52469 18683
rect 52503 18680 52515 18683
rect 52794 18683 52852 18689
rect 52794 18680 52806 18683
rect 52503 18652 52806 18680
rect 52503 18649 52515 18652
rect 52457 18643 52515 18649
rect 52794 18649 52806 18652
rect 52840 18649 52852 18683
rect 54021 18683 54079 18689
rect 54021 18680 54033 18683
rect 52794 18643 52852 18649
rect 52932 18652 54033 18680
rect 52932 18612 52960 18652
rect 54021 18649 54033 18652
rect 54067 18649 54079 18683
rect 54021 18643 54079 18649
rect 52380 18584 52960 18612
rect 53926 18572 53932 18624
rect 53984 18572 53990 18624
rect 57072 18612 57100 18847
rect 58158 18844 58164 18856
rect 58216 18844 58222 18896
rect 57330 18816 57336 18828
rect 57256 18788 57336 18816
rect 57256 18757 57284 18788
rect 57330 18776 57336 18788
rect 57388 18776 57394 18828
rect 57716 18788 58388 18816
rect 57716 18757 57744 18788
rect 58360 18760 58388 18788
rect 57241 18751 57299 18757
rect 57241 18717 57253 18751
rect 57287 18717 57299 18751
rect 57241 18711 57299 18717
rect 57425 18751 57483 18757
rect 57425 18717 57437 18751
rect 57471 18748 57483 18751
rect 57701 18751 57759 18757
rect 57701 18748 57713 18751
rect 57471 18720 57713 18748
rect 57471 18717 57483 18720
rect 57425 18711 57483 18717
rect 57701 18717 57713 18720
rect 57747 18717 57759 18751
rect 57701 18711 57759 18717
rect 57790 18708 57796 18760
rect 57848 18748 57854 18760
rect 57885 18751 57943 18757
rect 57885 18748 57897 18751
rect 57848 18720 57897 18748
rect 57848 18708 57854 18720
rect 57885 18717 57897 18720
rect 57931 18717 57943 18751
rect 57885 18711 57943 18717
rect 58066 18708 58072 18760
rect 58124 18708 58130 18760
rect 58342 18708 58348 18760
rect 58400 18708 58406 18760
rect 58529 18751 58587 18757
rect 58529 18717 58541 18751
rect 58575 18748 58587 18751
rect 58894 18748 58900 18760
rect 58575 18720 58900 18748
rect 58575 18717 58587 18720
rect 58529 18711 58587 18717
rect 58894 18708 58900 18720
rect 58952 18708 58958 18760
rect 57333 18683 57391 18689
rect 57333 18649 57345 18683
rect 57379 18680 57391 18683
rect 57379 18652 58112 18680
rect 57379 18649 57391 18652
rect 57333 18643 57391 18649
rect 58084 18624 58112 18652
rect 57882 18612 57888 18624
rect 57072 18584 57888 18612
rect 57882 18572 57888 18584
rect 57940 18572 57946 18624
rect 57974 18572 57980 18624
rect 58032 18572 58038 18624
rect 58066 18572 58072 18624
rect 58124 18572 58130 18624
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 3602 18368 3608 18420
rect 3660 18408 3666 18420
rect 3697 18411 3755 18417
rect 3697 18408 3709 18411
rect 3660 18380 3709 18408
rect 3660 18368 3666 18380
rect 3697 18377 3709 18380
rect 3743 18377 3755 18411
rect 3697 18371 3755 18377
rect 6822 18368 6828 18420
rect 6880 18408 6886 18420
rect 7929 18411 7987 18417
rect 7929 18408 7941 18411
rect 6880 18380 7941 18408
rect 6880 18368 6886 18380
rect 7929 18377 7941 18380
rect 7975 18377 7987 18411
rect 7929 18371 7987 18377
rect 46934 18368 46940 18420
rect 46992 18368 46998 18420
rect 47210 18368 47216 18420
rect 47268 18368 47274 18420
rect 47670 18368 47676 18420
rect 47728 18368 47734 18420
rect 48409 18411 48467 18417
rect 48409 18377 48421 18411
rect 48455 18408 48467 18411
rect 48590 18408 48596 18420
rect 48455 18380 48596 18408
rect 48455 18377 48467 18380
rect 48409 18371 48467 18377
rect 48590 18368 48596 18380
rect 48648 18368 48654 18420
rect 49142 18368 49148 18420
rect 49200 18368 49206 18420
rect 49326 18368 49332 18420
rect 49384 18368 49390 18420
rect 49878 18368 49884 18420
rect 49936 18368 49942 18420
rect 51718 18368 51724 18420
rect 51776 18408 51782 18420
rect 51905 18411 51963 18417
rect 51905 18408 51917 18411
rect 51776 18380 51917 18408
rect 51776 18368 51782 18380
rect 51905 18377 51917 18380
rect 51951 18377 51963 18411
rect 51905 18371 51963 18377
rect 52270 18368 52276 18420
rect 52328 18408 52334 18420
rect 53009 18411 53067 18417
rect 53009 18408 53021 18411
rect 52328 18380 53021 18408
rect 52328 18368 52334 18380
rect 53009 18377 53021 18380
rect 53055 18377 53067 18411
rect 53009 18371 53067 18377
rect 53650 18368 53656 18420
rect 53708 18408 53714 18420
rect 53708 18380 53788 18408
rect 53708 18368 53714 18380
rect 2498 18300 2504 18352
rect 2556 18340 2562 18352
rect 4522 18340 4528 18352
rect 2556 18312 4528 18340
rect 2556 18300 2562 18312
rect 4522 18300 4528 18312
rect 4580 18300 4586 18352
rect 5442 18300 5448 18352
rect 5500 18340 5506 18352
rect 5500 18312 6868 18340
rect 5500 18300 5506 18312
rect 2682 18232 2688 18284
rect 2740 18272 2746 18284
rect 4249 18275 4307 18281
rect 4249 18272 4261 18275
rect 2740 18244 4261 18272
rect 2740 18232 2746 18244
rect 4249 18241 4261 18244
rect 4295 18241 4307 18275
rect 4249 18235 4307 18241
rect 1578 18164 1584 18216
rect 1636 18164 1642 18216
rect 3510 18164 3516 18216
rect 3568 18164 3574 18216
rect 5902 18164 5908 18216
rect 5960 18164 5966 18216
rect 6181 18207 6239 18213
rect 6181 18173 6193 18207
rect 6227 18204 6239 18207
rect 6270 18204 6276 18216
rect 6227 18176 6276 18204
rect 6227 18173 6239 18176
rect 6181 18167 6239 18173
rect 6270 18164 6276 18176
rect 6328 18164 6334 18216
rect 6840 18204 6868 18312
rect 7006 18300 7012 18352
rect 7064 18340 7070 18352
rect 7064 18312 7788 18340
rect 7064 18300 7070 18312
rect 6914 18232 6920 18284
rect 6972 18232 6978 18284
rect 7760 18281 7788 18312
rect 8294 18300 8300 18352
rect 8352 18300 8358 18352
rect 9861 18343 9919 18349
rect 9861 18309 9873 18343
rect 9907 18309 9919 18343
rect 46952 18340 46980 18368
rect 47688 18340 47716 18368
rect 49160 18340 49188 18368
rect 46952 18312 47164 18340
rect 9861 18303 9919 18309
rect 7101 18275 7159 18281
rect 7101 18241 7113 18275
rect 7147 18272 7159 18275
rect 7193 18275 7251 18281
rect 7193 18272 7205 18275
rect 7147 18244 7205 18272
rect 7147 18241 7159 18244
rect 7101 18235 7159 18241
rect 7193 18241 7205 18244
rect 7239 18241 7251 18275
rect 7193 18235 7251 18241
rect 7745 18275 7803 18281
rect 7745 18241 7757 18275
rect 7791 18241 7803 18275
rect 7745 18235 7803 18241
rect 8312 18204 8340 18300
rect 9585 18275 9643 18281
rect 9585 18241 9597 18275
rect 9631 18272 9643 18275
rect 9674 18272 9680 18284
rect 9631 18244 9680 18272
rect 9631 18241 9643 18244
rect 9585 18235 9643 18241
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 9876 18272 9904 18303
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 9876 18244 11529 18272
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 11517 18235 11575 18241
rect 46937 18275 46995 18281
rect 46937 18241 46949 18275
rect 46983 18272 46995 18275
rect 47029 18275 47087 18281
rect 47029 18272 47041 18275
rect 46983 18244 47041 18272
rect 46983 18241 46995 18244
rect 46937 18235 46995 18241
rect 47029 18241 47041 18244
rect 47075 18241 47087 18275
rect 47029 18235 47087 18241
rect 6840 18176 8340 18204
rect 8481 18207 8539 18213
rect 8481 18173 8493 18207
rect 8527 18173 8539 18207
rect 8481 18167 8539 18173
rect 9861 18207 9919 18213
rect 9861 18173 9873 18207
rect 9907 18204 9919 18207
rect 10137 18207 10195 18213
rect 10137 18204 10149 18207
rect 9907 18176 10149 18204
rect 9907 18173 9919 18176
rect 9861 18167 9919 18173
rect 10137 18173 10149 18176
rect 10183 18173 10195 18207
rect 10137 18167 10195 18173
rect 10781 18207 10839 18213
rect 10781 18173 10793 18207
rect 10827 18204 10839 18207
rect 11054 18204 11060 18216
rect 10827 18176 11060 18204
rect 10827 18173 10839 18176
rect 10781 18167 10839 18173
rect 7009 18139 7067 18145
rect 7009 18105 7021 18139
rect 7055 18136 7067 18139
rect 8496 18136 8524 18167
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 46293 18207 46351 18213
rect 46293 18204 46305 18207
rect 46124 18176 46305 18204
rect 7055 18108 8524 18136
rect 9677 18139 9735 18145
rect 7055 18105 7067 18108
rect 7009 18099 7067 18105
rect 9677 18105 9689 18139
rect 9723 18136 9735 18139
rect 9950 18136 9956 18148
rect 9723 18108 9956 18136
rect 9723 18105 9735 18108
rect 9677 18099 9735 18105
rect 9950 18096 9956 18108
rect 10008 18096 10014 18148
rect 2866 18028 2872 18080
rect 2924 18068 2930 18080
rect 2961 18071 3019 18077
rect 2961 18068 2973 18071
rect 2924 18040 2973 18068
rect 2924 18028 2930 18040
rect 2961 18037 2973 18040
rect 3007 18037 3019 18071
rect 2961 18031 3019 18037
rect 4433 18071 4491 18077
rect 4433 18037 4445 18071
rect 4479 18068 4491 18071
rect 4706 18068 4712 18080
rect 4479 18040 4712 18068
rect 4479 18037 4491 18040
rect 4433 18031 4491 18037
rect 4706 18028 4712 18040
rect 4764 18028 4770 18080
rect 9214 18028 9220 18080
rect 9272 18028 9278 18080
rect 12158 18028 12164 18080
rect 12216 18028 12222 18080
rect 38654 18028 38660 18080
rect 38712 18068 38718 18080
rect 45646 18068 45652 18080
rect 38712 18040 45652 18068
rect 38712 18028 38718 18040
rect 45646 18028 45652 18040
rect 45704 18068 45710 18080
rect 46124 18077 46152 18176
rect 46293 18173 46305 18176
rect 46339 18173 46351 18207
rect 47136 18204 47164 18312
rect 47228 18312 48360 18340
rect 47228 18281 47256 18312
rect 47213 18275 47271 18281
rect 47213 18241 47225 18275
rect 47259 18241 47271 18275
rect 47213 18235 47271 18241
rect 47302 18232 47308 18284
rect 47360 18272 47366 18284
rect 48332 18281 48360 18312
rect 48516 18312 49188 18340
rect 49421 18343 49479 18349
rect 48516 18281 48544 18312
rect 49421 18309 49433 18343
rect 49467 18340 49479 18343
rect 49602 18340 49608 18352
rect 49467 18312 49608 18340
rect 49467 18309 49479 18312
rect 49421 18303 49479 18309
rect 49602 18300 49608 18312
rect 49660 18300 49666 18352
rect 48133 18275 48191 18281
rect 48133 18272 48145 18275
rect 47360 18244 48145 18272
rect 47360 18232 47366 18244
rect 48133 18241 48145 18244
rect 48179 18241 48191 18275
rect 48133 18235 48191 18241
rect 48317 18275 48375 18281
rect 48317 18241 48329 18275
rect 48363 18241 48375 18275
rect 48317 18235 48375 18241
rect 48501 18275 48559 18281
rect 48501 18241 48513 18275
rect 48547 18241 48559 18275
rect 48501 18235 48559 18241
rect 48866 18232 48872 18284
rect 48924 18272 48930 18284
rect 49145 18275 49203 18281
rect 49145 18272 49157 18275
rect 48924 18244 49157 18272
rect 48924 18232 48930 18244
rect 49145 18241 49157 18244
rect 49191 18241 49203 18275
rect 49145 18235 49203 18241
rect 49329 18275 49387 18281
rect 49329 18241 49341 18275
rect 49375 18272 49387 18275
rect 49896 18272 49924 18368
rect 53760 18349 53788 18380
rect 53926 18368 53932 18420
rect 53984 18368 53990 18420
rect 54665 18411 54723 18417
rect 54665 18377 54677 18411
rect 54711 18408 54723 18411
rect 54754 18408 54760 18420
rect 54711 18380 54760 18408
rect 54711 18377 54723 18380
rect 54665 18371 54723 18377
rect 51629 18343 51687 18349
rect 51629 18340 51641 18343
rect 51460 18312 51641 18340
rect 51460 18281 51488 18312
rect 51629 18309 51641 18312
rect 51675 18309 51687 18343
rect 52181 18343 52239 18349
rect 52181 18340 52193 18343
rect 51629 18303 51687 18309
rect 52012 18312 52193 18340
rect 49375 18244 49924 18272
rect 51261 18275 51319 18281
rect 49375 18241 49387 18244
rect 49329 18235 49387 18241
rect 51261 18241 51273 18275
rect 51307 18241 51319 18275
rect 51261 18235 51319 18241
rect 51445 18275 51503 18281
rect 51445 18241 51457 18275
rect 51491 18241 51503 18275
rect 51445 18235 51503 18241
rect 47581 18207 47639 18213
rect 47581 18204 47593 18207
rect 47136 18176 47593 18204
rect 46293 18167 46351 18173
rect 47581 18173 47593 18176
rect 47627 18173 47639 18207
rect 49160 18204 49188 18235
rect 51276 18204 51304 18235
rect 51534 18232 51540 18284
rect 51592 18232 51598 18284
rect 51718 18232 51724 18284
rect 51776 18232 51782 18284
rect 51810 18232 51816 18284
rect 51868 18232 51874 18284
rect 52012 18281 52040 18312
rect 52181 18309 52193 18312
rect 52227 18309 52239 18343
rect 52181 18303 52239 18309
rect 53745 18343 53803 18349
rect 53745 18309 53757 18343
rect 53791 18340 53803 18343
rect 53834 18340 53840 18352
rect 53791 18312 53840 18340
rect 53791 18309 53803 18312
rect 53745 18303 53803 18309
rect 53834 18300 53840 18312
rect 53892 18300 53898 18352
rect 53944 18340 53972 18368
rect 53944 18312 54064 18340
rect 51997 18275 52055 18281
rect 51997 18241 52009 18275
rect 52043 18241 52055 18275
rect 51997 18235 52055 18241
rect 52089 18275 52147 18281
rect 52089 18241 52101 18275
rect 52135 18241 52147 18275
rect 52089 18235 52147 18241
rect 52273 18275 52331 18281
rect 52273 18241 52285 18275
rect 52319 18241 52331 18275
rect 52273 18235 52331 18241
rect 53101 18275 53159 18281
rect 53101 18241 53113 18275
rect 53147 18272 53159 18275
rect 53558 18272 53564 18284
rect 53147 18244 53564 18272
rect 53147 18241 53159 18244
rect 53101 18235 53159 18241
rect 51828 18204 51856 18232
rect 49160 18176 51856 18204
rect 47581 18167 47639 18173
rect 51534 18096 51540 18148
rect 51592 18136 51598 18148
rect 52104 18136 52132 18235
rect 52288 18204 52316 18235
rect 53558 18232 53564 18244
rect 53616 18232 53622 18284
rect 53650 18232 53656 18284
rect 53708 18232 53714 18284
rect 54036 18281 54064 18312
rect 53929 18275 53987 18281
rect 53929 18241 53941 18275
rect 53975 18241 53987 18275
rect 53929 18235 53987 18241
rect 54021 18275 54079 18281
rect 54021 18241 54033 18275
rect 54067 18241 54079 18275
rect 54021 18235 54079 18241
rect 53834 18204 53840 18216
rect 52288 18176 53840 18204
rect 53834 18164 53840 18176
rect 53892 18164 53898 18216
rect 53944 18204 53972 18235
rect 54680 18204 54708 18371
rect 54754 18368 54760 18380
rect 54812 18368 54818 18420
rect 56594 18368 56600 18420
rect 56652 18408 56658 18420
rect 57333 18411 57391 18417
rect 57333 18408 57345 18411
rect 56652 18380 57345 18408
rect 56652 18368 56658 18380
rect 57333 18377 57345 18380
rect 57379 18377 57391 18411
rect 57333 18371 57391 18377
rect 55953 18275 56011 18281
rect 55953 18241 55965 18275
rect 55999 18272 56011 18275
rect 56962 18272 56968 18284
rect 55999 18244 56968 18272
rect 55999 18241 56011 18244
rect 55953 18235 56011 18241
rect 56962 18232 56968 18244
rect 57020 18232 57026 18284
rect 53944 18176 54708 18204
rect 57348 18204 57376 18371
rect 57974 18368 57980 18420
rect 58032 18368 58038 18420
rect 58066 18368 58072 18420
rect 58124 18368 58130 18420
rect 58342 18368 58348 18420
rect 58400 18368 58406 18420
rect 58894 18368 58900 18420
rect 58952 18368 58958 18420
rect 57992 18340 58020 18368
rect 57900 18312 58020 18340
rect 57900 18281 57928 18312
rect 57701 18275 57759 18281
rect 57701 18241 57713 18275
rect 57747 18241 57759 18275
rect 57701 18235 57759 18241
rect 57885 18275 57943 18281
rect 57885 18241 57897 18275
rect 57931 18241 57943 18275
rect 57885 18235 57943 18241
rect 57977 18275 58035 18281
rect 57977 18241 57989 18275
rect 58023 18272 58035 18275
rect 58084 18272 58112 18368
rect 58023 18244 58112 18272
rect 58161 18275 58219 18281
rect 58023 18241 58035 18244
rect 57977 18235 58035 18241
rect 58161 18241 58173 18275
rect 58207 18241 58219 18275
rect 58161 18235 58219 18241
rect 58529 18275 58587 18281
rect 58529 18241 58541 18275
rect 58575 18272 58587 18275
rect 58912 18272 58940 18368
rect 58575 18244 58940 18272
rect 58575 18241 58587 18244
rect 58529 18235 58587 18241
rect 57716 18204 57744 18235
rect 57790 18204 57796 18216
rect 57348 18176 57652 18204
rect 57716 18176 57796 18204
rect 57624 18148 57652 18176
rect 57790 18164 57796 18176
rect 57848 18164 57854 18216
rect 51592 18108 52132 18136
rect 51592 18096 51598 18108
rect 53558 18096 53564 18148
rect 53616 18136 53622 18148
rect 57517 18139 57575 18145
rect 57517 18136 57529 18139
rect 53616 18108 57529 18136
rect 53616 18096 53622 18108
rect 57517 18105 57529 18108
rect 57563 18105 57575 18139
rect 57517 18099 57575 18105
rect 57606 18096 57612 18148
rect 57664 18136 57670 18148
rect 58176 18136 58204 18235
rect 57664 18108 58204 18136
rect 57664 18096 57670 18108
rect 46109 18071 46167 18077
rect 46109 18068 46121 18071
rect 45704 18040 46121 18068
rect 45704 18028 45710 18040
rect 46109 18037 46121 18040
rect 46155 18037 46167 18071
rect 46109 18031 46167 18037
rect 49053 18071 49111 18077
rect 49053 18037 49065 18071
rect 49099 18068 49111 18071
rect 49786 18068 49792 18080
rect 49099 18040 49792 18068
rect 49099 18037 49111 18040
rect 49053 18031 49111 18037
rect 49786 18028 49792 18040
rect 49844 18028 49850 18080
rect 50893 18071 50951 18077
rect 50893 18037 50905 18071
rect 50939 18068 50951 18071
rect 50982 18068 50988 18080
rect 50939 18040 50988 18068
rect 50939 18037 50951 18040
rect 50893 18031 50951 18037
rect 50982 18028 50988 18040
rect 51040 18028 51046 18080
rect 51350 18028 51356 18080
rect 51408 18028 51414 18080
rect 53653 18071 53711 18077
rect 53653 18037 53665 18071
rect 53699 18068 53711 18071
rect 53742 18068 53748 18080
rect 53699 18040 53748 18068
rect 53699 18037 53711 18040
rect 53653 18031 53711 18037
rect 53742 18028 53748 18040
rect 53800 18028 53806 18080
rect 55214 18028 55220 18080
rect 55272 18068 55278 18080
rect 55861 18071 55919 18077
rect 55861 18068 55873 18071
rect 55272 18040 55873 18068
rect 55272 18028 55278 18040
rect 55861 18037 55873 18040
rect 55907 18037 55919 18071
rect 55861 18031 55919 18037
rect 58069 18071 58127 18077
rect 58069 18037 58081 18071
rect 58115 18068 58127 18071
rect 58342 18068 58348 18080
rect 58115 18040 58348 18068
rect 58115 18037 58127 18040
rect 58069 18031 58127 18037
rect 58342 18028 58348 18040
rect 58400 18028 58406 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 1397 17867 1455 17873
rect 1397 17833 1409 17867
rect 1443 17864 1455 17867
rect 2682 17864 2688 17876
rect 1443 17836 2688 17864
rect 1443 17833 1455 17836
rect 1397 17827 1455 17833
rect 2682 17824 2688 17836
rect 2740 17824 2746 17876
rect 3329 17867 3387 17873
rect 3329 17833 3341 17867
rect 3375 17864 3387 17867
rect 3510 17864 3516 17876
rect 3375 17836 3516 17864
rect 3375 17833 3387 17836
rect 3329 17827 3387 17833
rect 3510 17824 3516 17836
rect 3568 17824 3574 17876
rect 3786 17824 3792 17876
rect 3844 17824 3850 17876
rect 4614 17824 4620 17876
rect 4672 17824 4678 17876
rect 4801 17867 4859 17873
rect 4801 17833 4813 17867
rect 4847 17864 4859 17867
rect 4890 17864 4896 17876
rect 4847 17836 4896 17864
rect 4847 17833 4859 17836
rect 4801 17827 4859 17833
rect 4890 17824 4896 17836
rect 4948 17824 4954 17876
rect 9858 17864 9864 17876
rect 8404 17836 9864 17864
rect 2866 17688 2872 17740
rect 2924 17688 2930 17740
rect 3237 17731 3295 17737
rect 3237 17697 3249 17731
rect 3283 17728 3295 17731
rect 3804 17728 3832 17824
rect 4632 17796 4660 17824
rect 3283 17700 3832 17728
rect 3896 17768 4660 17796
rect 3283 17697 3295 17700
rect 3237 17691 3295 17697
rect 3142 17620 3148 17672
rect 3200 17620 3206 17672
rect 3421 17663 3479 17669
rect 3421 17629 3433 17663
rect 3467 17629 3479 17663
rect 3421 17623 3479 17629
rect 3513 17663 3571 17669
rect 3513 17629 3525 17663
rect 3559 17660 3571 17663
rect 3896 17660 3924 17768
rect 4706 17756 4712 17808
rect 4764 17796 4770 17808
rect 4764 17768 6132 17796
rect 4764 17756 4770 17768
rect 6104 17737 6132 17768
rect 4617 17731 4675 17737
rect 4617 17697 4629 17731
rect 4663 17728 4675 17731
rect 5353 17731 5411 17737
rect 5353 17728 5365 17731
rect 4663 17700 5365 17728
rect 4663 17697 4675 17700
rect 4617 17691 4675 17697
rect 5353 17697 5365 17700
rect 5399 17697 5411 17731
rect 5353 17691 5411 17697
rect 6089 17731 6147 17737
rect 6089 17697 6101 17731
rect 6135 17697 6147 17731
rect 6089 17691 6147 17697
rect 3559 17632 3924 17660
rect 3559 17629 3571 17632
rect 3513 17623 3571 17629
rect 2406 17552 2412 17604
rect 2464 17552 2470 17604
rect 2222 17484 2228 17536
rect 2280 17524 2286 17536
rect 3436 17524 3464 17623
rect 4062 17620 4068 17672
rect 4120 17660 4126 17672
rect 4525 17663 4583 17669
rect 4525 17660 4537 17663
rect 4120 17632 4537 17660
rect 4120 17620 4126 17632
rect 4525 17629 4537 17632
rect 4571 17629 4583 17663
rect 4525 17623 4583 17629
rect 4709 17663 4767 17669
rect 4709 17629 4721 17663
rect 4755 17660 4767 17663
rect 5537 17663 5595 17669
rect 5537 17660 5549 17663
rect 4755 17632 5549 17660
rect 4755 17629 4767 17632
rect 4709 17623 4767 17629
rect 5537 17629 5549 17632
rect 5583 17629 5595 17663
rect 6914 17660 6920 17672
rect 5537 17623 5595 17629
rect 5644 17632 6920 17660
rect 4540 17592 4568 17623
rect 5644 17592 5672 17632
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 8404 17669 8432 17836
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 11974 17824 11980 17876
rect 12032 17864 12038 17876
rect 12253 17867 12311 17873
rect 12253 17864 12265 17867
rect 12032 17836 12265 17864
rect 12032 17824 12038 17836
rect 12253 17833 12265 17836
rect 12299 17833 12311 17867
rect 12253 17827 12311 17833
rect 48314 17824 48320 17876
rect 48372 17864 48378 17876
rect 49602 17864 49608 17876
rect 48372 17836 49608 17864
rect 48372 17824 48378 17836
rect 49602 17824 49608 17836
rect 49660 17864 49666 17876
rect 49697 17867 49755 17873
rect 49697 17864 49709 17867
rect 49660 17836 49709 17864
rect 49660 17824 49666 17836
rect 49697 17833 49709 17836
rect 49743 17833 49755 17867
rect 49697 17827 49755 17833
rect 50062 17824 50068 17876
rect 50120 17864 50126 17876
rect 50157 17867 50215 17873
rect 50157 17864 50169 17867
rect 50120 17836 50169 17864
rect 50120 17824 50126 17836
rect 50157 17833 50169 17836
rect 50203 17833 50215 17867
rect 50157 17827 50215 17833
rect 53558 17824 53564 17876
rect 53616 17824 53622 17876
rect 53834 17824 53840 17876
rect 53892 17864 53898 17876
rect 54021 17867 54079 17873
rect 54021 17864 54033 17867
rect 53892 17836 54033 17864
rect 53892 17824 53898 17836
rect 54021 17833 54033 17836
rect 54067 17833 54079 17867
rect 54021 17827 54079 17833
rect 54846 17824 54852 17876
rect 54904 17864 54910 17876
rect 54941 17867 54999 17873
rect 54941 17864 54953 17867
rect 54904 17836 54953 17864
rect 54904 17824 54910 17836
rect 54941 17833 54953 17836
rect 54987 17833 54999 17867
rect 54941 17827 54999 17833
rect 55214 17824 55220 17876
rect 55272 17824 55278 17876
rect 57882 17824 57888 17876
rect 57940 17864 57946 17876
rect 57974 17864 57980 17876
rect 57940 17836 57980 17864
rect 57940 17824 57946 17836
rect 57974 17824 57980 17836
rect 58032 17824 58038 17876
rect 58250 17824 58256 17876
rect 58308 17824 58314 17876
rect 8573 17799 8631 17805
rect 8573 17765 8585 17799
rect 8619 17796 8631 17799
rect 8619 17768 9444 17796
rect 8619 17765 8631 17768
rect 8573 17759 8631 17765
rect 8662 17688 8668 17740
rect 8720 17688 8726 17740
rect 9416 17737 9444 17768
rect 11992 17737 12020 17824
rect 49421 17799 49479 17805
rect 49421 17765 49433 17799
rect 49467 17765 49479 17799
rect 53576 17796 53604 17824
rect 55232 17796 55260 17824
rect 49421 17759 49479 17765
rect 53300 17768 53604 17796
rect 54864 17768 55260 17796
rect 56689 17799 56747 17805
rect 9401 17731 9459 17737
rect 8772 17700 9352 17728
rect 8389 17663 8447 17669
rect 8389 17629 8401 17663
rect 8435 17629 8447 17663
rect 8389 17623 8447 17629
rect 8481 17663 8539 17669
rect 8481 17629 8493 17663
rect 8527 17660 8539 17663
rect 8772 17660 8800 17700
rect 8527 17632 8800 17660
rect 9125 17663 9183 17669
rect 8527 17629 8539 17632
rect 8481 17623 8539 17629
rect 9125 17629 9137 17663
rect 9171 17660 9183 17663
rect 9324 17660 9352 17700
rect 9401 17697 9413 17731
rect 9447 17697 9459 17731
rect 9401 17691 9459 17697
rect 11977 17731 12035 17737
rect 11977 17697 11989 17731
rect 12023 17697 12035 17731
rect 11977 17691 12035 17697
rect 9950 17660 9956 17672
rect 9171 17632 9260 17660
rect 9324 17632 9956 17660
rect 9171 17629 9183 17632
rect 9125 17623 9183 17629
rect 4540 17564 5672 17592
rect 6638 17552 6644 17604
rect 6696 17592 6702 17604
rect 8496 17592 8524 17623
rect 6696 17564 8524 17592
rect 6696 17552 6702 17564
rect 9030 17552 9036 17604
rect 9088 17552 9094 17604
rect 9232 17536 9260 17632
rect 9950 17620 9956 17632
rect 10008 17620 10014 17672
rect 10318 17620 10324 17672
rect 10376 17660 10382 17672
rect 10376 17632 10626 17660
rect 10376 17620 10382 17632
rect 47854 17620 47860 17672
rect 47912 17620 47918 17672
rect 49145 17663 49203 17669
rect 49145 17629 49157 17663
rect 49191 17629 49203 17663
rect 49145 17623 49203 17629
rect 11701 17595 11759 17601
rect 11701 17561 11713 17595
rect 11747 17592 11759 17595
rect 12158 17592 12164 17604
rect 11747 17564 12164 17592
rect 11747 17561 11759 17564
rect 11701 17555 11759 17561
rect 12158 17552 12164 17564
rect 12216 17552 12222 17604
rect 49160 17536 49188 17623
rect 49234 17620 49240 17672
rect 49292 17620 49298 17672
rect 49436 17660 49464 17759
rect 50157 17663 50215 17669
rect 50157 17660 50169 17663
rect 49436 17632 50169 17660
rect 50157 17629 50169 17632
rect 50203 17629 50215 17663
rect 50157 17623 50215 17629
rect 50341 17663 50399 17669
rect 50341 17629 50353 17663
rect 50387 17660 50399 17663
rect 51350 17660 51356 17672
rect 50387 17632 51356 17660
rect 50387 17629 50399 17632
rect 50341 17623 50399 17629
rect 51350 17620 51356 17632
rect 51408 17620 51414 17672
rect 53300 17669 53328 17768
rect 53377 17731 53435 17737
rect 53377 17697 53389 17731
rect 53423 17728 53435 17731
rect 53423 17700 53604 17728
rect 53423 17697 53435 17700
rect 53377 17691 53435 17697
rect 53576 17669 53604 17700
rect 53285 17663 53343 17669
rect 53285 17629 53297 17663
rect 53331 17629 53343 17663
rect 53285 17623 53343 17629
rect 53469 17663 53527 17669
rect 53469 17629 53481 17663
rect 53515 17629 53527 17663
rect 53469 17623 53527 17629
rect 53561 17663 53619 17669
rect 53561 17629 53573 17663
rect 53607 17629 53619 17663
rect 53561 17623 53619 17629
rect 49252 17592 49280 17620
rect 49421 17595 49479 17601
rect 49421 17592 49433 17595
rect 49252 17564 49433 17592
rect 49421 17561 49433 17564
rect 49467 17592 49479 17595
rect 49602 17592 49608 17604
rect 49467 17564 49608 17592
rect 49467 17561 49479 17564
rect 49421 17555 49479 17561
rect 49602 17552 49608 17564
rect 49660 17552 49666 17604
rect 53374 17552 53380 17604
rect 53432 17592 53438 17604
rect 53484 17592 53512 17623
rect 53742 17620 53748 17672
rect 53800 17660 53806 17672
rect 53837 17663 53895 17669
rect 53837 17660 53849 17663
rect 53800 17632 53849 17660
rect 53800 17620 53806 17632
rect 53837 17629 53849 17632
rect 53883 17629 53895 17663
rect 53837 17623 53895 17629
rect 53926 17620 53932 17672
rect 53984 17620 53990 17672
rect 54864 17669 54892 17768
rect 56689 17765 56701 17799
rect 56735 17765 56747 17799
rect 56689 17759 56747 17765
rect 57793 17799 57851 17805
rect 57793 17765 57805 17799
rect 57839 17796 57851 17799
rect 57839 17768 58388 17796
rect 57839 17765 57851 17768
rect 57793 17759 57851 17765
rect 55122 17688 55128 17740
rect 55180 17688 55186 17740
rect 56704 17728 56732 17759
rect 56781 17731 56839 17737
rect 56781 17728 56793 17731
rect 56704 17700 56793 17728
rect 56781 17697 56793 17700
rect 56827 17697 56839 17731
rect 56781 17691 56839 17697
rect 57440 17700 57928 17728
rect 54113 17663 54171 17669
rect 54113 17629 54125 17663
rect 54159 17629 54171 17663
rect 54113 17623 54171 17629
rect 54849 17663 54907 17669
rect 54849 17629 54861 17663
rect 54895 17629 54907 17663
rect 54849 17623 54907 17629
rect 53432 17564 53512 17592
rect 53653 17595 53711 17601
rect 53432 17552 53438 17564
rect 53653 17561 53665 17595
rect 53699 17561 53711 17595
rect 54128 17592 54156 17623
rect 55306 17620 55312 17672
rect 55364 17620 55370 17672
rect 53653 17555 53711 17561
rect 53760 17564 54156 17592
rect 55125 17595 55183 17601
rect 2280 17496 3464 17524
rect 2280 17484 2286 17496
rect 9214 17484 9220 17536
rect 9272 17484 9278 17536
rect 10042 17484 10048 17536
rect 10100 17484 10106 17536
rect 10226 17484 10232 17536
rect 10284 17484 10290 17536
rect 47302 17484 47308 17536
rect 47360 17484 47366 17536
rect 49142 17484 49148 17536
rect 49200 17484 49206 17536
rect 49234 17484 49240 17536
rect 49292 17484 49298 17536
rect 52730 17484 52736 17536
rect 52788 17524 52794 17536
rect 53101 17527 53159 17533
rect 53101 17524 53113 17527
rect 52788 17496 53113 17524
rect 52788 17484 52794 17496
rect 53101 17493 53113 17496
rect 53147 17524 53159 17527
rect 53668 17524 53696 17555
rect 53760 17533 53788 17564
rect 55125 17561 55137 17595
rect 55171 17592 55183 17595
rect 55554 17595 55612 17601
rect 55554 17592 55566 17595
rect 55171 17564 55566 17592
rect 55171 17561 55183 17564
rect 55125 17555 55183 17561
rect 55554 17561 55566 17564
rect 55600 17561 55612 17595
rect 55554 17555 55612 17561
rect 53147 17496 53696 17524
rect 53745 17527 53803 17533
rect 53147 17493 53159 17496
rect 53101 17487 53159 17493
rect 53745 17493 53757 17527
rect 53791 17493 53803 17527
rect 53745 17487 53803 17493
rect 56502 17484 56508 17536
rect 56560 17524 56566 17536
rect 57440 17533 57468 17700
rect 57517 17663 57575 17669
rect 57517 17629 57529 17663
rect 57563 17660 57575 17663
rect 57606 17660 57612 17672
rect 57563 17632 57612 17660
rect 57563 17629 57575 17632
rect 57517 17623 57575 17629
rect 57606 17620 57612 17632
rect 57664 17620 57670 17672
rect 57900 17669 57928 17700
rect 58066 17671 58072 17672
rect 57793 17663 57851 17669
rect 57793 17629 57805 17663
rect 57839 17629 57851 17663
rect 57793 17623 57851 17629
rect 57885 17663 57943 17669
rect 57885 17629 57897 17663
rect 57931 17629 57943 17663
rect 57885 17623 57943 17629
rect 58044 17665 58072 17671
rect 58044 17631 58056 17665
rect 58044 17625 58072 17631
rect 57698 17552 57704 17604
rect 57756 17552 57762 17604
rect 57425 17527 57483 17533
rect 57425 17524 57437 17527
rect 56560 17496 57437 17524
rect 56560 17484 56566 17496
rect 57425 17493 57437 17496
rect 57471 17493 57483 17527
rect 57808 17524 57836 17623
rect 58066 17620 58072 17625
rect 58124 17620 58130 17672
rect 58161 17663 58219 17669
rect 58161 17629 58173 17663
rect 58207 17662 58219 17663
rect 58250 17662 58256 17672
rect 58207 17634 58256 17662
rect 58207 17629 58219 17634
rect 58161 17623 58219 17629
rect 58250 17620 58256 17634
rect 58308 17620 58314 17672
rect 58360 17669 58388 17768
rect 58345 17663 58403 17669
rect 58345 17629 58357 17663
rect 58391 17629 58403 17663
rect 58345 17623 58403 17629
rect 58069 17527 58127 17533
rect 58069 17524 58081 17527
rect 57808 17496 58081 17524
rect 57425 17487 57483 17493
rect 58069 17493 58081 17496
rect 58115 17493 58127 17527
rect 58069 17487 58127 17493
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 5534 17320 5540 17332
rect 2424 17292 4384 17320
rect 2222 17144 2228 17196
rect 2280 17144 2286 17196
rect 2424 17193 2452 17292
rect 2685 17255 2743 17261
rect 2685 17221 2697 17255
rect 2731 17252 2743 17255
rect 2731 17224 2820 17252
rect 2731 17221 2743 17224
rect 2685 17215 2743 17221
rect 2792 17193 2820 17224
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17153 2467 17187
rect 2409 17147 2467 17153
rect 2777 17187 2835 17193
rect 2777 17153 2789 17187
rect 2823 17153 2835 17187
rect 2777 17147 2835 17153
rect 2240 17116 2268 17144
rect 2501 17119 2559 17125
rect 2501 17116 2513 17119
rect 2240 17088 2513 17116
rect 2501 17085 2513 17088
rect 2547 17085 2559 17119
rect 2501 17079 2559 17085
rect 2685 17119 2743 17125
rect 2685 17085 2697 17119
rect 2731 17116 2743 17119
rect 3513 17119 3571 17125
rect 3513 17116 3525 17119
rect 2731 17088 3525 17116
rect 2731 17085 2743 17088
rect 2685 17079 2743 17085
rect 3513 17085 3525 17088
rect 3559 17085 3571 17119
rect 3513 17079 3571 17085
rect 2516 17048 2544 17079
rect 4154 17076 4160 17128
rect 4212 17076 4218 17128
rect 4356 17048 4384 17292
rect 4448 17292 5540 17320
rect 4448 17193 4476 17292
rect 5534 17280 5540 17292
rect 5592 17280 5598 17332
rect 6178 17280 6184 17332
rect 6236 17280 6242 17332
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8720 17292 9045 17320
rect 8720 17280 8726 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9033 17283 9091 17289
rect 11054 17280 11060 17332
rect 11112 17280 11118 17332
rect 11238 17280 11244 17332
rect 11296 17280 11302 17332
rect 47302 17280 47308 17332
rect 47360 17280 47366 17332
rect 47673 17323 47731 17329
rect 47673 17289 47685 17323
rect 47719 17320 47731 17323
rect 47854 17320 47860 17332
rect 47719 17292 47860 17320
rect 47719 17289 47731 17292
rect 47673 17283 47731 17289
rect 47854 17280 47860 17292
rect 47912 17280 47918 17332
rect 48682 17280 48688 17332
rect 48740 17320 48746 17332
rect 49145 17323 49203 17329
rect 48740 17292 49096 17320
rect 48740 17280 48746 17292
rect 4709 17255 4767 17261
rect 4709 17221 4721 17255
rect 4755 17221 4767 17255
rect 4709 17215 4767 17221
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17153 4491 17187
rect 4724 17184 4752 17215
rect 4801 17187 4859 17193
rect 4801 17184 4813 17187
rect 4724 17156 4813 17184
rect 4433 17147 4491 17153
rect 4801 17153 4813 17156
rect 4847 17153 4859 17187
rect 6196 17184 6224 17280
rect 6733 17255 6791 17261
rect 6733 17221 6745 17255
rect 6779 17252 6791 17255
rect 6779 17224 6868 17252
rect 6779 17221 6791 17224
rect 6733 17215 6791 17221
rect 4801 17147 4859 17153
rect 5644 17156 6224 17184
rect 4709 17119 4767 17125
rect 4709 17085 4721 17119
rect 4755 17116 4767 17119
rect 5537 17119 5595 17125
rect 5537 17116 5549 17119
rect 4755 17088 5549 17116
rect 4755 17085 4767 17088
rect 4709 17079 4767 17085
rect 5537 17085 5549 17088
rect 5583 17085 5595 17119
rect 5537 17079 5595 17085
rect 5644 17048 5672 17156
rect 6454 17144 6460 17196
rect 6512 17144 6518 17196
rect 6549 17187 6607 17193
rect 6549 17153 6561 17187
rect 6595 17184 6607 17187
rect 6638 17184 6644 17196
rect 6595 17156 6644 17184
rect 6595 17153 6607 17156
rect 6549 17147 6607 17153
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 6840 17193 6868 17224
rect 6914 17212 6920 17264
rect 6972 17252 6978 17264
rect 11256 17252 11284 17280
rect 47320 17252 47348 17280
rect 6972 17224 11284 17252
rect 6972 17212 6978 17224
rect 9968 17193 9996 17224
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 8941 17187 8999 17193
rect 8941 17153 8953 17187
rect 8987 17184 8999 17187
rect 9769 17187 9827 17193
rect 9769 17184 9781 17187
rect 8987 17156 9781 17184
rect 8987 17153 8999 17156
rect 8941 17147 8999 17153
rect 9769 17153 9781 17156
rect 9815 17153 9827 17187
rect 9769 17147 9827 17153
rect 9953 17187 10011 17193
rect 9953 17153 9965 17187
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 10873 17187 10931 17193
rect 10873 17153 10885 17187
rect 10919 17184 10931 17187
rect 10965 17187 11023 17193
rect 10965 17184 10977 17187
rect 10919 17156 10977 17184
rect 10919 17153 10931 17156
rect 10873 17147 10931 17153
rect 10965 17153 10977 17156
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 11149 17187 11207 17193
rect 11149 17153 11161 17187
rect 11195 17184 11207 17187
rect 11256 17184 11284 17224
rect 11195 17156 11284 17184
rect 46952 17224 47348 17252
rect 11195 17153 11207 17156
rect 11149 17147 11207 17153
rect 6178 17076 6184 17128
rect 6236 17076 6242 17128
rect 6733 17119 6791 17125
rect 6733 17085 6745 17119
rect 6779 17116 6791 17119
rect 7561 17119 7619 17125
rect 7561 17116 7573 17119
rect 6779 17088 7573 17116
rect 6779 17085 6791 17088
rect 6733 17079 6791 17085
rect 7561 17085 7573 17088
rect 7607 17085 7619 17119
rect 7561 17079 7619 17085
rect 8110 17076 8116 17128
rect 8168 17076 8174 17128
rect 8389 17119 8447 17125
rect 8389 17085 8401 17119
rect 8435 17116 8447 17119
rect 9030 17116 9036 17128
rect 8435 17088 9036 17116
rect 8435 17085 8447 17088
rect 8389 17079 8447 17085
rect 9030 17076 9036 17088
rect 9088 17076 9094 17128
rect 9677 17119 9735 17125
rect 9677 17085 9689 17119
rect 9723 17116 9735 17119
rect 9861 17119 9919 17125
rect 9861 17116 9873 17119
rect 9723 17088 9873 17116
rect 9723 17085 9735 17088
rect 9677 17079 9735 17085
rect 9861 17085 9873 17088
rect 9907 17085 9919 17119
rect 9861 17079 9919 17085
rect 10226 17076 10232 17128
rect 10284 17076 10290 17128
rect 46952 17125 46980 17224
rect 48038 17212 48044 17264
rect 48096 17252 48102 17264
rect 48961 17255 49019 17261
rect 48096 17224 48820 17252
rect 48096 17212 48102 17224
rect 48792 17196 48820 17224
rect 48961 17221 48973 17255
rect 49007 17221 49019 17255
rect 49068 17252 49096 17292
rect 49145 17289 49157 17323
rect 49191 17320 49203 17323
rect 49234 17320 49240 17332
rect 49191 17292 49240 17320
rect 49191 17289 49203 17292
rect 49145 17283 49203 17289
rect 49234 17280 49240 17292
rect 49292 17280 49298 17332
rect 55122 17280 55128 17332
rect 55180 17320 55186 17332
rect 55585 17323 55643 17329
rect 55585 17320 55597 17323
rect 55180 17292 55597 17320
rect 55180 17280 55186 17292
rect 55585 17289 55597 17292
rect 55631 17289 55643 17323
rect 55585 17283 55643 17289
rect 56962 17280 56968 17332
rect 57020 17280 57026 17332
rect 57241 17323 57299 17329
rect 57241 17289 57253 17323
rect 57287 17320 57299 17323
rect 57698 17320 57704 17332
rect 57287 17292 57704 17320
rect 57287 17289 57299 17292
rect 57241 17283 57299 17289
rect 57698 17280 57704 17292
rect 57756 17280 57762 17332
rect 57974 17280 57980 17332
rect 58032 17320 58038 17332
rect 58250 17320 58256 17332
rect 58032 17292 58256 17320
rect 58032 17280 58038 17292
rect 58250 17280 58256 17292
rect 58308 17280 58314 17332
rect 58345 17323 58403 17329
rect 58345 17289 58357 17323
rect 58391 17289 58403 17323
rect 58345 17283 58403 17289
rect 49068 17224 49280 17252
rect 48961 17215 49019 17221
rect 47213 17187 47271 17193
rect 47213 17153 47225 17187
rect 47259 17184 47271 17187
rect 47581 17187 47639 17193
rect 47259 17156 47532 17184
rect 47259 17153 47271 17156
rect 47213 17147 47271 17153
rect 46937 17119 46995 17125
rect 46937 17085 46949 17119
rect 46983 17085 46995 17119
rect 46937 17079 46995 17085
rect 2516 17020 4292 17048
rect 4356 17020 5672 17048
rect 47504 17048 47532 17156
rect 47581 17153 47593 17187
rect 47627 17184 47639 17187
rect 47765 17187 47823 17193
rect 47627 17156 47716 17184
rect 47627 17153 47639 17156
rect 47581 17147 47639 17153
rect 47688 17128 47716 17156
rect 47765 17153 47777 17187
rect 47811 17184 47823 17187
rect 48593 17187 48651 17193
rect 48593 17184 48605 17187
rect 47811 17156 48605 17184
rect 47811 17153 47823 17156
rect 47765 17147 47823 17153
rect 48593 17153 48605 17156
rect 48639 17184 48651 17187
rect 48685 17187 48743 17193
rect 48685 17184 48697 17187
rect 48639 17156 48697 17184
rect 48639 17153 48651 17156
rect 48593 17147 48651 17153
rect 48685 17153 48697 17156
rect 48731 17153 48743 17187
rect 48685 17147 48743 17153
rect 48774 17144 48780 17196
rect 48832 17144 48838 17196
rect 48976 17184 49004 17215
rect 49252 17193 49280 17224
rect 55398 17212 55404 17264
rect 55456 17252 55462 17264
rect 56980 17252 57008 17280
rect 58360 17252 58388 17283
rect 55456 17224 56364 17252
rect 55456 17212 55462 17224
rect 49053 17187 49111 17193
rect 49053 17184 49065 17187
rect 48976 17156 49065 17184
rect 49053 17153 49065 17156
rect 49099 17153 49111 17187
rect 49053 17147 49111 17153
rect 49237 17187 49295 17193
rect 49237 17153 49249 17187
rect 49283 17153 49295 17187
rect 49237 17147 49295 17153
rect 49326 17144 49332 17196
rect 49384 17144 49390 17196
rect 56336 17193 56364 17224
rect 56980 17224 58388 17252
rect 49513 17187 49571 17193
rect 49513 17153 49525 17187
rect 49559 17153 49571 17187
rect 49513 17147 49571 17153
rect 56321 17187 56379 17193
rect 56321 17153 56333 17187
rect 56367 17153 56379 17187
rect 56321 17147 56379 17153
rect 47670 17076 47676 17128
rect 47728 17076 47734 17128
rect 48038 17076 48044 17128
rect 48096 17076 48102 17128
rect 48961 17119 49019 17125
rect 48148 17088 48912 17116
rect 48148 17048 48176 17088
rect 47504 17020 48176 17048
rect 3418 16940 3424 16992
rect 3476 16940 3482 16992
rect 4264 16980 4292 17020
rect 48774 17008 48780 17060
rect 48832 17008 48838 17060
rect 48884 17048 48912 17088
rect 48961 17085 48973 17119
rect 49007 17116 49019 17119
rect 49421 17119 49479 17125
rect 49421 17116 49433 17119
rect 49007 17088 49433 17116
rect 49007 17085 49019 17088
rect 48961 17079 49019 17085
rect 49421 17085 49433 17088
rect 49467 17085 49479 17119
rect 49421 17079 49479 17085
rect 49528 17048 49556 17147
rect 56502 17144 56508 17196
rect 56560 17144 56566 17196
rect 56980 17184 57008 17224
rect 57057 17187 57115 17193
rect 57057 17184 57069 17187
rect 56980 17156 57069 17184
rect 57057 17153 57069 17156
rect 57103 17153 57115 17187
rect 57057 17147 57115 17153
rect 57241 17187 57299 17193
rect 57241 17153 57253 17187
rect 57287 17184 57299 17187
rect 57330 17184 57336 17196
rect 57287 17156 57336 17184
rect 57287 17153 57299 17156
rect 57241 17147 57299 17153
rect 57330 17144 57336 17156
rect 57388 17144 57394 17196
rect 57606 17144 57612 17196
rect 57664 17144 57670 17196
rect 57977 17187 58035 17193
rect 57977 17153 57989 17187
rect 58023 17153 58035 17187
rect 57977 17147 58035 17153
rect 58161 17187 58219 17193
rect 58161 17153 58173 17187
rect 58207 17184 58219 17187
rect 58342 17184 58348 17196
rect 58207 17156 58348 17184
rect 58207 17153 58219 17156
rect 58161 17147 58219 17153
rect 56229 17119 56287 17125
rect 56229 17085 56241 17119
rect 56275 17116 56287 17119
rect 56413 17119 56471 17125
rect 56413 17116 56425 17119
rect 56275 17088 56425 17116
rect 56275 17085 56287 17088
rect 56229 17079 56287 17085
rect 56413 17085 56425 17088
rect 56459 17085 56471 17119
rect 56413 17079 56471 17085
rect 48884 17020 49556 17048
rect 4525 16983 4583 16989
rect 4525 16980 4537 16983
rect 4264 16952 4537 16980
rect 4525 16949 4537 16952
rect 4571 16980 4583 16983
rect 4798 16980 4804 16992
rect 4571 16952 4804 16980
rect 4571 16949 4583 16952
rect 4525 16943 4583 16949
rect 4798 16940 4804 16952
rect 4856 16940 4862 16992
rect 5442 16940 5448 16992
rect 5500 16940 5506 16992
rect 7466 16940 7472 16992
rect 7524 16940 7530 16992
rect 46934 16940 46940 16992
rect 46992 16980 46998 16992
rect 47029 16983 47087 16989
rect 47029 16980 47041 16983
rect 46992 16952 47041 16980
rect 46992 16940 46998 16952
rect 47029 16949 47041 16952
rect 47075 16949 47087 16983
rect 47029 16943 47087 16949
rect 47118 16940 47124 16992
rect 47176 16940 47182 16992
rect 48792 16980 48820 17008
rect 49344 16992 49372 17020
rect 57992 16992 58020 17147
rect 58342 17144 58348 17156
rect 58400 17144 58406 17196
rect 58529 17187 58587 17193
rect 58529 17153 58541 17187
rect 58575 17184 58587 17187
rect 58575 17156 58940 17184
rect 58575 17153 58587 17156
rect 58529 17147 58587 17153
rect 58912 17060 58940 17156
rect 58069 17051 58127 17057
rect 58069 17017 58081 17051
rect 58115 17048 58127 17051
rect 58158 17048 58164 17060
rect 58115 17020 58164 17048
rect 58115 17017 58127 17020
rect 58069 17011 58127 17017
rect 58158 17008 58164 17020
rect 58216 17008 58222 17060
rect 58894 17008 58900 17060
rect 58952 17008 58958 17060
rect 49234 16980 49240 16992
rect 48792 16952 49240 16980
rect 49234 16940 49240 16952
rect 49292 16940 49298 16992
rect 49326 16940 49332 16992
rect 49384 16940 49390 16992
rect 52730 16940 52736 16992
rect 52788 16980 52794 16992
rect 53101 16983 53159 16989
rect 53101 16980 53113 16983
rect 52788 16952 53113 16980
rect 52788 16940 52794 16952
rect 53101 16949 53113 16952
rect 53147 16949 53159 16983
rect 53101 16943 53159 16949
rect 57974 16940 57980 16992
rect 58032 16940 58038 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 3163 16779 3221 16785
rect 3163 16745 3175 16779
rect 3209 16776 3221 16779
rect 3418 16776 3424 16788
rect 3209 16748 3424 16776
rect 3209 16745 3221 16748
rect 3163 16739 3221 16745
rect 3418 16736 3424 16748
rect 3476 16736 3482 16788
rect 5442 16736 5448 16788
rect 5500 16776 5506 16788
rect 5825 16779 5883 16785
rect 5825 16776 5837 16779
rect 5500 16748 5837 16776
rect 5500 16736 5506 16748
rect 5825 16745 5837 16748
rect 5871 16745 5883 16779
rect 5825 16739 5883 16745
rect 6178 16736 6184 16788
rect 6236 16776 6242 16788
rect 6273 16779 6331 16785
rect 6273 16776 6285 16779
rect 6236 16748 6285 16776
rect 6236 16736 6242 16748
rect 6273 16745 6285 16748
rect 6319 16745 6331 16779
rect 6273 16739 6331 16745
rect 7466 16736 7472 16788
rect 7524 16776 7530 16788
rect 8217 16779 8275 16785
rect 8217 16776 8229 16779
rect 7524 16748 8229 16776
rect 7524 16736 7530 16748
rect 8217 16745 8229 16748
rect 8263 16745 8275 16779
rect 8217 16739 8275 16745
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 10517 16779 10575 16785
rect 10517 16776 10529 16779
rect 10100 16748 10529 16776
rect 10100 16736 10106 16748
rect 10517 16745 10529 16748
rect 10563 16745 10575 16779
rect 47026 16776 47032 16788
rect 10517 16739 10575 16745
rect 46676 16748 47032 16776
rect 3142 16600 3148 16652
rect 3200 16640 3206 16652
rect 3421 16643 3479 16649
rect 3421 16640 3433 16643
rect 3200 16612 3433 16640
rect 3200 16600 3206 16612
rect 3421 16609 3433 16612
rect 3467 16640 3479 16643
rect 6089 16643 6147 16649
rect 6089 16640 6101 16643
rect 3467 16612 6101 16640
rect 3467 16609 3479 16612
rect 3421 16603 3479 16609
rect 6089 16609 6101 16612
rect 6135 16640 6147 16643
rect 6270 16640 6276 16652
rect 6135 16612 6276 16640
rect 6135 16609 6147 16612
rect 6089 16603 6147 16609
rect 6270 16600 6276 16612
rect 6328 16640 6334 16652
rect 8481 16643 8539 16649
rect 8481 16640 8493 16643
rect 6328 16612 8493 16640
rect 6328 16600 6334 16612
rect 8481 16609 8493 16612
rect 8527 16640 8539 16643
rect 9766 16640 9772 16652
rect 8527 16612 9772 16640
rect 8527 16609 8539 16612
rect 8481 16603 8539 16609
rect 9766 16600 9772 16612
rect 9824 16640 9830 16652
rect 10781 16643 10839 16649
rect 10781 16640 10793 16643
rect 9824 16612 10793 16640
rect 9824 16600 9830 16612
rect 10781 16609 10793 16612
rect 10827 16609 10839 16643
rect 10781 16603 10839 16609
rect 45922 16600 45928 16652
rect 45980 16640 45986 16652
rect 46676 16649 46704 16748
rect 47026 16736 47032 16748
rect 47084 16736 47090 16788
rect 48038 16736 48044 16788
rect 48096 16736 48102 16788
rect 48682 16736 48688 16788
rect 48740 16776 48746 16788
rect 48869 16779 48927 16785
rect 48869 16776 48881 16779
rect 48740 16748 48881 16776
rect 48740 16736 48746 16748
rect 48869 16745 48881 16748
rect 48915 16776 48927 16779
rect 49234 16776 49240 16788
rect 48915 16748 49240 16776
rect 48915 16745 48927 16748
rect 48869 16739 48927 16745
rect 49234 16736 49240 16748
rect 49292 16736 49298 16788
rect 49418 16736 49424 16788
rect 49476 16776 49482 16788
rect 49789 16779 49847 16785
rect 49789 16776 49801 16779
rect 49476 16748 49801 16776
rect 49476 16736 49482 16748
rect 49789 16745 49801 16748
rect 49835 16745 49847 16779
rect 50890 16776 50896 16788
rect 49789 16739 49847 16745
rect 50172 16748 50896 16776
rect 46661 16643 46719 16649
rect 46661 16640 46673 16643
rect 45980 16612 46673 16640
rect 45980 16600 45986 16612
rect 46661 16609 46673 16612
rect 46707 16609 46719 16643
rect 46661 16603 46719 16609
rect 49620 16612 49832 16640
rect 3786 16532 3792 16584
rect 3844 16532 3850 16584
rect 3970 16532 3976 16584
rect 4028 16532 4034 16584
rect 4062 16532 4068 16584
rect 4120 16532 4126 16584
rect 6181 16575 6239 16581
rect 4264 16558 4738 16572
rect 4264 16544 4752 16558
rect 3881 16507 3939 16513
rect 2714 16476 2774 16504
rect 1670 16396 1676 16448
rect 1728 16396 1734 16448
rect 2406 16396 2412 16448
rect 2464 16436 2470 16448
rect 2746 16436 2774 16476
rect 3881 16473 3893 16507
rect 3927 16504 3939 16507
rect 4080 16504 4108 16532
rect 3927 16476 4108 16504
rect 3927 16473 3939 16476
rect 3881 16467 3939 16473
rect 4264 16436 4292 16544
rect 2464 16408 4292 16436
rect 4341 16439 4399 16445
rect 2464 16396 2470 16408
rect 4341 16405 4353 16439
rect 4387 16436 4399 16439
rect 4522 16436 4528 16448
rect 4387 16408 4528 16436
rect 4387 16405 4399 16408
rect 4341 16399 4399 16405
rect 4522 16396 4528 16408
rect 4580 16396 4586 16448
rect 4724 16436 4752 16544
rect 6181 16541 6193 16575
rect 6227 16541 6239 16575
rect 6181 16535 6239 16541
rect 5350 16464 5356 16516
rect 5408 16504 5414 16516
rect 6196 16504 6224 16535
rect 6362 16532 6368 16584
rect 6420 16532 6426 16584
rect 6914 16532 6920 16584
rect 6972 16532 6978 16584
rect 46934 16581 46940 16584
rect 46928 16572 46940 16581
rect 46895 16544 46940 16572
rect 46928 16535 46940 16544
rect 46934 16532 46940 16535
rect 46992 16532 46998 16584
rect 47670 16532 47676 16584
rect 47728 16572 47734 16584
rect 49620 16572 49648 16612
rect 47728 16544 49648 16572
rect 49697 16575 49755 16581
rect 47728 16532 47734 16544
rect 49697 16541 49709 16575
rect 49743 16541 49755 16575
rect 49804 16572 49832 16612
rect 49970 16600 49976 16652
rect 50028 16600 50034 16652
rect 50172 16649 50200 16748
rect 50890 16736 50896 16748
rect 50948 16736 50954 16788
rect 52822 16736 52828 16788
rect 52880 16736 52886 16788
rect 52914 16736 52920 16788
rect 52972 16736 52978 16788
rect 53466 16736 53472 16788
rect 53524 16776 53530 16788
rect 53653 16779 53711 16785
rect 53653 16776 53665 16779
rect 53524 16748 53665 16776
rect 53524 16736 53530 16748
rect 53653 16745 53665 16748
rect 53699 16745 53711 16779
rect 53653 16739 53711 16745
rect 57790 16736 57796 16788
rect 57848 16736 57854 16788
rect 57974 16736 57980 16788
rect 58032 16736 58038 16788
rect 51537 16711 51595 16717
rect 51537 16677 51549 16711
rect 51583 16677 51595 16711
rect 52840 16708 52868 16736
rect 53558 16708 53564 16720
rect 52840 16680 53564 16708
rect 51537 16671 51595 16677
rect 50157 16643 50215 16649
rect 50157 16609 50169 16643
rect 50203 16609 50215 16643
rect 51552 16640 51580 16671
rect 53558 16668 53564 16680
rect 53616 16708 53622 16720
rect 54205 16711 54263 16717
rect 54205 16708 54217 16711
rect 53616 16680 54217 16708
rect 53616 16668 53622 16680
rect 51629 16643 51687 16649
rect 51629 16640 51641 16643
rect 51552 16612 51641 16640
rect 50157 16603 50215 16609
rect 51629 16609 51641 16612
rect 51675 16609 51687 16643
rect 51629 16603 51687 16609
rect 52730 16600 52736 16652
rect 52788 16640 52794 16652
rect 52788 16612 53512 16640
rect 52788 16600 52794 16612
rect 51166 16572 51172 16584
rect 49804 16544 51172 16572
rect 49697 16535 49755 16541
rect 6932 16504 6960 16532
rect 5408 16476 5488 16504
rect 6196 16476 6960 16504
rect 7774 16476 9168 16504
rect 10074 16476 10364 16504
rect 5408 16464 5414 16476
rect 5460 16436 5488 16476
rect 4724 16408 5488 16436
rect 6730 16396 6736 16448
rect 6788 16396 6794 16448
rect 9030 16396 9036 16448
rect 9088 16396 9094 16448
rect 9140 16436 9168 16476
rect 10336 16448 10364 16476
rect 10318 16436 10324 16448
rect 9140 16408 10324 16436
rect 10318 16396 10324 16408
rect 10376 16396 10382 16448
rect 49712 16436 49740 16535
rect 51166 16532 51172 16544
rect 51224 16532 51230 16584
rect 52457 16575 52515 16581
rect 52457 16572 52469 16575
rect 52288 16544 52469 16572
rect 49973 16507 50031 16513
rect 49973 16473 49985 16507
rect 50019 16504 50031 16507
rect 50402 16507 50460 16513
rect 50402 16504 50414 16507
rect 50019 16476 50414 16504
rect 50019 16473 50031 16476
rect 49973 16467 50031 16473
rect 50402 16473 50414 16476
rect 50448 16473 50460 16507
rect 51810 16504 51816 16516
rect 50402 16467 50460 16473
rect 51046 16476 51816 16504
rect 51046 16436 51074 16476
rect 51810 16464 51816 16476
rect 51868 16464 51874 16516
rect 49712 16408 51074 16436
rect 51258 16396 51264 16448
rect 51316 16436 51322 16448
rect 52288 16445 52316 16544
rect 52457 16541 52469 16544
rect 52503 16541 52515 16575
rect 52457 16535 52515 16541
rect 52549 16575 52607 16581
rect 52549 16541 52561 16575
rect 52595 16541 52607 16575
rect 52549 16535 52607 16541
rect 52641 16575 52699 16581
rect 52641 16541 52653 16575
rect 52687 16572 52699 16575
rect 52687 16544 53162 16572
rect 52687 16541 52699 16544
rect 52641 16535 52699 16541
rect 52564 16448 52592 16535
rect 52914 16464 52920 16516
rect 52972 16464 52978 16516
rect 53134 16504 53162 16544
rect 53190 16532 53196 16584
rect 53248 16532 53254 16584
rect 53282 16532 53288 16584
rect 53340 16532 53346 16584
rect 53484 16581 53512 16612
rect 53469 16575 53527 16581
rect 53469 16541 53481 16575
rect 53515 16541 53527 16575
rect 53469 16535 53527 16541
rect 53558 16532 53564 16584
rect 53616 16572 53622 16584
rect 53760 16581 53788 16680
rect 54205 16677 54217 16680
rect 54251 16708 54263 16711
rect 56413 16711 56471 16717
rect 56413 16708 56425 16711
rect 54251 16680 56425 16708
rect 54251 16677 54263 16680
rect 54205 16671 54263 16677
rect 56413 16677 56425 16680
rect 56459 16708 56471 16711
rect 56870 16708 56876 16720
rect 56459 16680 56876 16708
rect 56459 16677 56471 16680
rect 56413 16671 56471 16677
rect 56870 16668 56876 16680
rect 56928 16668 56934 16720
rect 58345 16711 58403 16717
rect 58345 16677 58357 16711
rect 58391 16677 58403 16711
rect 58345 16671 58403 16677
rect 58360 16640 58388 16671
rect 55600 16612 57974 16640
rect 55600 16584 55628 16612
rect 53653 16575 53711 16581
rect 53653 16572 53665 16575
rect 53616 16544 53665 16572
rect 53616 16532 53622 16544
rect 53653 16541 53665 16544
rect 53699 16541 53711 16575
rect 53653 16535 53711 16541
rect 53745 16575 53803 16581
rect 53745 16541 53757 16575
rect 53791 16541 53803 16575
rect 53745 16535 53803 16541
rect 55582 16532 55588 16584
rect 55640 16532 55646 16584
rect 56594 16532 56600 16584
rect 56652 16532 56658 16584
rect 57946 16572 57974 16612
rect 58084 16612 58388 16640
rect 58084 16572 58112 16612
rect 57946 16544 58112 16572
rect 58158 16532 58164 16584
rect 58216 16532 58222 16584
rect 58529 16575 58587 16581
rect 58529 16541 58541 16575
rect 58575 16572 58587 16575
rect 58575 16544 58940 16572
rect 58575 16541 58587 16544
rect 58529 16535 58587 16541
rect 53929 16507 53987 16513
rect 53134 16476 53696 16504
rect 53668 16448 53696 16476
rect 53929 16473 53941 16507
rect 53975 16473 53987 16507
rect 53929 16467 53987 16473
rect 52273 16439 52331 16445
rect 52273 16436 52285 16439
rect 51316 16408 52285 16436
rect 51316 16396 51322 16408
rect 52273 16405 52285 16408
rect 52319 16405 52331 16439
rect 52273 16399 52331 16405
rect 52546 16396 52552 16448
rect 52604 16396 52610 16448
rect 52822 16396 52828 16448
rect 52880 16396 52886 16448
rect 53101 16439 53159 16445
rect 53101 16405 53113 16439
rect 53147 16436 53159 16439
rect 53285 16439 53343 16445
rect 53285 16436 53297 16439
rect 53147 16408 53297 16436
rect 53147 16405 53159 16408
rect 53101 16399 53159 16405
rect 53285 16405 53297 16408
rect 53331 16405 53343 16439
rect 53285 16399 53343 16405
rect 53650 16396 53656 16448
rect 53708 16396 53714 16448
rect 53944 16436 53972 16467
rect 56870 16464 56876 16516
rect 56928 16504 56934 16516
rect 57885 16507 57943 16513
rect 57885 16504 57897 16507
rect 56928 16476 57897 16504
rect 56928 16464 56934 16476
rect 57885 16473 57897 16476
rect 57931 16473 57943 16507
rect 57885 16467 57943 16473
rect 58069 16507 58127 16513
rect 58069 16473 58081 16507
rect 58115 16473 58127 16507
rect 58069 16467 58127 16473
rect 54110 16436 54116 16448
rect 53944 16408 54116 16436
rect 54110 16396 54116 16408
rect 54168 16396 54174 16448
rect 55490 16396 55496 16448
rect 55548 16396 55554 16448
rect 56778 16396 56784 16448
rect 56836 16436 56842 16448
rect 57241 16439 57299 16445
rect 57241 16436 57253 16439
rect 56836 16408 57253 16436
rect 56836 16396 56842 16408
rect 57241 16405 57253 16408
rect 57287 16405 57299 16439
rect 57241 16399 57299 16405
rect 57974 16396 57980 16448
rect 58032 16436 58038 16448
rect 58084 16436 58112 16467
rect 58912 16448 58940 16544
rect 58032 16408 58112 16436
rect 58032 16396 58038 16408
rect 58894 16396 58900 16448
rect 58952 16396 58958 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 3513 16235 3571 16241
rect 3513 16201 3525 16235
rect 3559 16232 3571 16235
rect 3786 16232 3792 16244
rect 3559 16204 3792 16232
rect 3559 16201 3571 16204
rect 3513 16195 3571 16201
rect 3786 16192 3792 16204
rect 3844 16192 3850 16244
rect 6362 16192 6368 16244
rect 6420 16192 6426 16244
rect 6914 16192 6920 16244
rect 6972 16192 6978 16244
rect 7285 16235 7343 16241
rect 7285 16201 7297 16235
rect 7331 16232 7343 16235
rect 8110 16232 8116 16244
rect 7331 16204 8116 16232
rect 7331 16201 7343 16204
rect 7285 16195 7343 16201
rect 8110 16192 8116 16204
rect 8168 16192 8174 16244
rect 48501 16235 48559 16241
rect 48501 16201 48513 16235
rect 48547 16232 48559 16235
rect 48869 16235 48927 16241
rect 48869 16232 48881 16235
rect 48547 16204 48881 16232
rect 48547 16201 48559 16204
rect 48501 16195 48559 16201
rect 48869 16201 48881 16204
rect 48915 16201 48927 16235
rect 49145 16235 49203 16241
rect 49145 16232 49157 16235
rect 48869 16195 48927 16201
rect 48976 16204 49157 16232
rect 6932 16164 6960 16192
rect 44085 16167 44143 16173
rect 6932 16136 7236 16164
rect 934 16056 940 16108
rect 992 16096 998 16108
rect 1581 16099 1639 16105
rect 1581 16096 1593 16099
rect 992 16068 1593 16096
rect 992 16056 998 16068
rect 1581 16065 1593 16068
rect 1627 16065 1639 16099
rect 1581 16059 1639 16065
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16096 2743 16099
rect 4706 16096 4712 16108
rect 2731 16068 4712 16096
rect 2731 16065 2743 16068
rect 2685 16059 2743 16065
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 6730 16056 6736 16108
rect 6788 16096 6794 16108
rect 7208 16105 7236 16136
rect 44085 16133 44097 16167
rect 44131 16164 44143 16167
rect 44177 16167 44235 16173
rect 44177 16164 44189 16167
rect 44131 16136 44189 16164
rect 44131 16133 44143 16136
rect 44085 16127 44143 16133
rect 44177 16133 44189 16136
rect 44223 16164 44235 16167
rect 48314 16164 48320 16176
rect 44223 16136 48320 16164
rect 44223 16133 44235 16136
rect 44177 16127 44235 16133
rect 48314 16124 48320 16136
rect 48372 16124 48378 16176
rect 7193 16099 7251 16105
rect 6788 16068 7052 16096
rect 6788 16056 6794 16068
rect 1670 15988 1676 16040
rect 1728 16028 1734 16040
rect 2869 16031 2927 16037
rect 2869 16028 2881 16031
rect 1728 16000 2881 16028
rect 1728 15988 1734 16000
rect 2700 15904 2728 16000
rect 2869 15997 2881 16000
rect 2915 15997 2927 16031
rect 2869 15991 2927 15997
rect 4614 15988 4620 16040
rect 4672 16028 4678 16040
rect 6917 16031 6975 16037
rect 6917 16028 6929 16031
rect 4672 16000 6929 16028
rect 4672 15988 4678 16000
rect 6917 15997 6929 16000
rect 6963 15997 6975 16031
rect 7024 16028 7052 16068
rect 7193 16065 7205 16099
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 7377 16099 7435 16105
rect 7377 16065 7389 16099
rect 7423 16096 7435 16099
rect 7929 16099 7987 16105
rect 7929 16096 7941 16099
rect 7423 16068 7941 16096
rect 7423 16065 7435 16068
rect 7377 16059 7435 16065
rect 7929 16065 7941 16068
rect 7975 16065 7987 16099
rect 7929 16059 7987 16065
rect 45922 16056 45928 16108
rect 45980 16056 45986 16108
rect 47670 16056 47676 16108
rect 47728 16096 47734 16108
rect 47857 16099 47915 16105
rect 47857 16096 47869 16099
rect 47728 16068 47869 16096
rect 47728 16056 47734 16068
rect 47857 16065 47869 16068
rect 47903 16065 47915 16099
rect 47857 16059 47915 16065
rect 48038 16056 48044 16108
rect 48096 16056 48102 16108
rect 48406 16056 48412 16108
rect 48464 16056 48470 16108
rect 48593 16099 48651 16105
rect 48593 16065 48605 16099
rect 48639 16096 48651 16099
rect 48682 16096 48688 16108
rect 48639 16068 48688 16096
rect 48639 16065 48651 16068
rect 48593 16059 48651 16065
rect 48682 16056 48688 16068
rect 48740 16056 48746 16108
rect 48777 16099 48835 16105
rect 48777 16065 48789 16099
rect 48823 16065 48835 16099
rect 48777 16059 48835 16065
rect 8481 16031 8539 16037
rect 8481 16028 8493 16031
rect 7024 16000 8493 16028
rect 6917 15991 6975 15997
rect 8481 15997 8493 16000
rect 8527 15997 8539 16031
rect 8481 15991 8539 15997
rect 44818 15988 44824 16040
rect 44876 16028 44882 16040
rect 48498 16028 48504 16040
rect 44876 16000 48504 16028
rect 44876 15988 44882 16000
rect 48498 15988 48504 16000
rect 48556 15988 48562 16040
rect 48792 16028 48820 16059
rect 48976 16028 49004 16204
rect 49145 16201 49157 16204
rect 49191 16201 49203 16235
rect 49145 16195 49203 16201
rect 49234 16192 49240 16244
rect 49292 16232 49298 16244
rect 49697 16235 49755 16241
rect 49697 16232 49709 16235
rect 49292 16204 49709 16232
rect 49292 16192 49298 16204
rect 49697 16201 49709 16204
rect 49743 16201 49755 16235
rect 49697 16195 49755 16201
rect 49970 16192 49976 16244
rect 50028 16232 50034 16244
rect 50341 16235 50399 16241
rect 50341 16232 50353 16235
rect 50028 16204 50353 16232
rect 50028 16192 50034 16204
rect 50341 16201 50353 16204
rect 50387 16201 50399 16235
rect 50341 16195 50399 16201
rect 52822 16192 52828 16244
rect 52880 16192 52886 16244
rect 53009 16235 53067 16241
rect 53009 16201 53021 16235
rect 53055 16232 53067 16235
rect 53282 16232 53288 16244
rect 53055 16204 53288 16232
rect 53055 16201 53067 16204
rect 53009 16195 53067 16201
rect 53282 16192 53288 16204
rect 53340 16192 53346 16244
rect 53558 16192 53564 16244
rect 53616 16192 53622 16244
rect 54110 16192 54116 16244
rect 54168 16192 54174 16244
rect 55582 16232 55588 16244
rect 54220 16204 55588 16232
rect 49602 16164 49608 16176
rect 49068 16136 49608 16164
rect 49068 16105 49096 16136
rect 49602 16124 49608 16136
rect 49660 16124 49666 16176
rect 52181 16167 52239 16173
rect 52181 16133 52193 16167
rect 52227 16164 52239 16167
rect 52840 16164 52868 16192
rect 52227 16136 52592 16164
rect 52840 16136 53052 16164
rect 52227 16133 52239 16136
rect 52181 16127 52239 16133
rect 49053 16099 49111 16105
rect 49053 16065 49065 16099
rect 49099 16065 49111 16099
rect 49053 16059 49111 16065
rect 49145 16099 49203 16105
rect 49145 16065 49157 16099
rect 49191 16065 49203 16099
rect 49145 16059 49203 16065
rect 49329 16099 49387 16105
rect 49329 16065 49341 16099
rect 49375 16096 49387 16099
rect 49375 16068 49464 16096
rect 49375 16065 49387 16068
rect 49329 16059 49387 16065
rect 48792 16000 49004 16028
rect 48314 15920 48320 15972
rect 48372 15960 48378 15972
rect 49160 15960 49188 16059
rect 49436 15972 49464 16068
rect 51074 16056 51080 16108
rect 51132 16056 51138 16108
rect 51258 16056 51264 16108
rect 51316 16056 51322 16108
rect 52089 16099 52147 16105
rect 52089 16065 52101 16099
rect 52135 16065 52147 16099
rect 52089 16059 52147 16065
rect 52273 16099 52331 16105
rect 52273 16065 52285 16099
rect 52319 16065 52331 16099
rect 52564 16096 52592 16136
rect 53024 16105 53052 16136
rect 53374 16124 53380 16176
rect 53432 16124 53438 16176
rect 53650 16124 53656 16176
rect 53708 16124 53714 16176
rect 54220 16164 54248 16204
rect 55582 16192 55588 16204
rect 55640 16192 55646 16244
rect 56505 16235 56563 16241
rect 56505 16201 56517 16235
rect 56551 16232 56563 16235
rect 56594 16232 56600 16244
rect 56551 16204 56600 16232
rect 56551 16201 56563 16204
rect 56505 16195 56563 16201
rect 56594 16192 56600 16204
rect 56652 16192 56658 16244
rect 57330 16192 57336 16244
rect 57388 16192 57394 16244
rect 58161 16235 58219 16241
rect 58161 16232 58173 16235
rect 57532 16204 58173 16232
rect 53760 16136 54248 16164
rect 54389 16167 54447 16173
rect 52825 16099 52883 16105
rect 52825 16096 52837 16099
rect 52564 16068 52837 16096
rect 52273 16059 52331 16065
rect 52825 16065 52837 16068
rect 52871 16065 52883 16099
rect 52825 16059 52883 16065
rect 53009 16099 53067 16105
rect 53009 16065 53021 16099
rect 53055 16065 53067 16099
rect 53392 16096 53420 16124
rect 53561 16099 53619 16105
rect 53561 16096 53573 16099
rect 53392 16068 53573 16096
rect 53009 16059 53067 16065
rect 53561 16065 53573 16068
rect 53607 16065 53619 16099
rect 53561 16059 53619 16065
rect 50985 16031 51043 16037
rect 50985 15997 50997 16031
rect 51031 16028 51043 16031
rect 51169 16031 51227 16037
rect 51169 16028 51181 16031
rect 51031 16000 51181 16028
rect 51031 15997 51043 16000
rect 50985 15991 51043 15997
rect 51169 15997 51181 16000
rect 51215 15997 51227 16031
rect 51169 15991 51227 15997
rect 48372 15932 49188 15960
rect 48372 15920 48378 15932
rect 49418 15920 49424 15972
rect 49476 15920 49482 15972
rect 2682 15852 2688 15904
rect 2740 15852 2746 15904
rect 47946 15852 47952 15904
rect 48004 15852 48010 15904
rect 49053 15895 49111 15901
rect 49053 15861 49065 15895
rect 49099 15892 49111 15895
rect 49510 15892 49516 15904
rect 49099 15864 49516 15892
rect 49099 15861 49111 15864
rect 49053 15855 49111 15861
rect 49510 15852 49516 15864
rect 49568 15852 49574 15904
rect 51810 15852 51816 15904
rect 51868 15892 51874 15904
rect 52104 15892 52132 16059
rect 52288 15960 52316 16059
rect 52546 15988 52552 16040
rect 52604 16028 52610 16040
rect 53668 16028 53696 16124
rect 53760 16105 53788 16136
rect 54389 16133 54401 16167
rect 54435 16164 54447 16167
rect 56778 16164 56784 16176
rect 54435 16136 56784 16164
rect 54435 16133 54447 16136
rect 54389 16127 54447 16133
rect 56778 16124 56784 16136
rect 56836 16124 56842 16176
rect 56870 16124 56876 16176
rect 56928 16124 56934 16176
rect 57348 16164 57376 16192
rect 57532 16173 57560 16204
rect 58161 16201 58173 16204
rect 58207 16201 58219 16235
rect 58161 16195 58219 16201
rect 57517 16167 57575 16173
rect 57348 16136 57468 16164
rect 55398 16105 55404 16108
rect 53745 16099 53803 16105
rect 53745 16065 53757 16099
rect 53791 16065 53803 16099
rect 53745 16059 53803 16065
rect 54113 16099 54171 16105
rect 54113 16065 54125 16099
rect 54159 16065 54171 16099
rect 54113 16059 54171 16065
rect 54205 16099 54263 16105
rect 54205 16065 54217 16099
rect 54251 16065 54263 16099
rect 54205 16059 54263 16065
rect 55392 16059 55404 16105
rect 54128 16028 54156 16059
rect 52604 16000 53512 16028
rect 53668 16000 54156 16028
rect 52604 15988 52610 16000
rect 53374 15960 53380 15972
rect 52288 15932 53380 15960
rect 53374 15920 53380 15932
rect 53432 15920 53438 15972
rect 53484 15960 53512 16000
rect 54018 15960 54024 15972
rect 53484 15932 54024 15960
rect 54018 15920 54024 15932
rect 54076 15960 54082 15972
rect 54220 15960 54248 16059
rect 55398 16056 55404 16059
rect 55456 16056 55462 16108
rect 56888 16096 56916 16124
rect 57333 16099 57391 16105
rect 57333 16096 57345 16099
rect 56888 16068 57345 16096
rect 57333 16065 57345 16068
rect 57379 16065 57391 16099
rect 57333 16059 57391 16065
rect 55125 16031 55183 16037
rect 55125 15997 55137 16031
rect 55171 15997 55183 16031
rect 55125 15991 55183 15997
rect 54076 15932 54248 15960
rect 54076 15920 54082 15932
rect 53098 15892 53104 15904
rect 51868 15864 53104 15892
rect 51868 15852 51874 15864
rect 53098 15852 53104 15864
rect 53156 15852 53162 15904
rect 55140 15892 55168 15991
rect 57146 15988 57152 16040
rect 57204 15988 57210 16040
rect 57440 16028 57468 16136
rect 57517 16133 57529 16167
rect 57563 16133 57575 16167
rect 57977 16167 58035 16173
rect 57977 16164 57989 16167
rect 57517 16127 57575 16133
rect 57624 16136 57989 16164
rect 57624 16105 57652 16136
rect 57977 16133 57989 16136
rect 58023 16133 58035 16167
rect 58526 16164 58532 16176
rect 57977 16127 58035 16133
rect 58084 16136 58532 16164
rect 57609 16099 57667 16105
rect 57609 16065 57621 16099
rect 57655 16065 57667 16099
rect 57609 16059 57667 16065
rect 57790 16056 57796 16108
rect 57848 16096 57854 16108
rect 58084 16105 58112 16136
rect 58526 16124 58532 16136
rect 58584 16124 58590 16176
rect 57885 16099 57943 16105
rect 57885 16096 57897 16099
rect 57848 16068 57897 16096
rect 57848 16056 57854 16068
rect 57885 16065 57897 16068
rect 57931 16065 57943 16099
rect 57885 16059 57943 16065
rect 58069 16099 58127 16105
rect 58069 16065 58081 16099
rect 58115 16065 58127 16099
rect 58069 16059 58127 16065
rect 58161 16099 58219 16105
rect 58161 16065 58173 16099
rect 58207 16065 58219 16099
rect 58161 16059 58219 16065
rect 57698 16028 57704 16040
rect 57440 16000 57704 16028
rect 57698 15988 57704 16000
rect 57756 16028 57762 16040
rect 58176 16028 58204 16059
rect 58342 16056 58348 16108
rect 58400 16056 58406 16108
rect 57756 16000 58204 16028
rect 57756 15988 57762 16000
rect 57609 15963 57667 15969
rect 57609 15929 57621 15963
rect 57655 15960 57667 15963
rect 57882 15960 57888 15972
rect 57655 15932 57888 15960
rect 57655 15929 57667 15932
rect 57609 15923 57667 15929
rect 57882 15920 57888 15932
rect 57940 15920 57946 15972
rect 55306 15892 55312 15904
rect 55140 15864 55312 15892
rect 55306 15852 55312 15864
rect 55364 15852 55370 15904
rect 56594 15852 56600 15904
rect 56652 15852 56658 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 47946 15648 47952 15700
rect 48004 15648 48010 15700
rect 49697 15691 49755 15697
rect 49697 15657 49709 15691
rect 49743 15688 49755 15691
rect 49878 15688 49884 15700
rect 49743 15660 49884 15688
rect 49743 15657 49755 15660
rect 49697 15651 49755 15657
rect 49878 15648 49884 15660
rect 49936 15648 49942 15700
rect 50249 15691 50307 15697
rect 50249 15657 50261 15691
rect 50295 15688 50307 15691
rect 50706 15688 50712 15700
rect 50295 15660 50712 15688
rect 50295 15657 50307 15660
rect 50249 15651 50307 15657
rect 50706 15648 50712 15660
rect 50764 15648 50770 15700
rect 51626 15648 51632 15700
rect 51684 15688 51690 15700
rect 51905 15691 51963 15697
rect 51905 15688 51917 15691
rect 51684 15660 51917 15688
rect 51684 15648 51690 15660
rect 51905 15657 51917 15660
rect 51951 15657 51963 15691
rect 51905 15651 51963 15657
rect 52914 15648 52920 15700
rect 52972 15648 52978 15700
rect 53466 15648 53472 15700
rect 53524 15648 53530 15700
rect 53745 15691 53803 15697
rect 53745 15657 53757 15691
rect 53791 15688 53803 15691
rect 53926 15688 53932 15700
rect 53791 15660 53932 15688
rect 53791 15657 53803 15660
rect 53745 15651 53803 15657
rect 53926 15648 53932 15660
rect 53984 15648 53990 15700
rect 55398 15648 55404 15700
rect 55456 15688 55462 15700
rect 55493 15691 55551 15697
rect 55493 15688 55505 15691
rect 55456 15660 55505 15688
rect 55456 15648 55462 15660
rect 55493 15657 55505 15660
rect 55539 15657 55551 15691
rect 55493 15651 55551 15657
rect 56594 15648 56600 15700
rect 56652 15648 56658 15700
rect 56689 15691 56747 15697
rect 56689 15657 56701 15691
rect 56735 15688 56747 15691
rect 57146 15688 57152 15700
rect 56735 15660 57152 15688
rect 56735 15657 56747 15660
rect 56689 15651 56747 15657
rect 57146 15648 57152 15660
rect 57204 15648 57210 15700
rect 57698 15648 57704 15700
rect 57756 15648 57762 15700
rect 57974 15648 57980 15700
rect 58032 15648 58038 15700
rect 58158 15648 58164 15700
rect 58216 15688 58222 15700
rect 58253 15691 58311 15697
rect 58253 15688 58265 15691
rect 58216 15660 58265 15688
rect 58216 15648 58222 15660
rect 58253 15657 58265 15660
rect 58299 15657 58311 15691
rect 58253 15651 58311 15657
rect 47397 15623 47455 15629
rect 47397 15589 47409 15623
rect 47443 15589 47455 15623
rect 47397 15583 47455 15589
rect 45922 15512 45928 15564
rect 45980 15552 45986 15564
rect 46017 15555 46075 15561
rect 46017 15552 46029 15555
rect 45980 15524 46029 15552
rect 45980 15512 45986 15524
rect 46017 15521 46029 15524
rect 46063 15521 46075 15555
rect 46017 15515 46075 15521
rect 47412 15484 47440 15583
rect 47964 15552 47992 15648
rect 49234 15580 49240 15632
rect 49292 15620 49298 15632
rect 52549 15623 52607 15629
rect 52549 15620 52561 15623
rect 49292 15592 52561 15620
rect 49292 15580 49298 15592
rect 48041 15555 48099 15561
rect 48041 15552 48053 15555
rect 47964 15524 48053 15552
rect 48041 15521 48053 15524
rect 48087 15521 48099 15555
rect 51810 15552 51816 15564
rect 48041 15515 48099 15521
rect 50632 15524 51816 15552
rect 48777 15487 48835 15493
rect 48777 15484 48789 15487
rect 47412 15456 48789 15484
rect 48777 15453 48789 15456
rect 48823 15453 48835 15487
rect 48777 15447 48835 15453
rect 49053 15487 49111 15493
rect 49053 15453 49065 15487
rect 49099 15453 49111 15487
rect 49053 15447 49111 15453
rect 46284 15419 46342 15425
rect 46284 15385 46296 15419
rect 46330 15416 46342 15419
rect 46566 15416 46572 15428
rect 46330 15388 46572 15416
rect 46330 15385 46342 15388
rect 46284 15379 46342 15385
rect 46566 15376 46572 15388
rect 46624 15376 46630 15428
rect 48498 15376 48504 15428
rect 48556 15416 48562 15428
rect 49068 15416 49096 15447
rect 49234 15444 49240 15496
rect 49292 15444 49298 15496
rect 49326 15444 49332 15496
rect 49384 15444 49390 15496
rect 49418 15444 49424 15496
rect 49476 15493 49482 15496
rect 49476 15487 49525 15493
rect 49476 15453 49479 15487
rect 49513 15484 49525 15487
rect 50062 15484 50068 15496
rect 49513 15456 50068 15484
rect 49513 15453 49525 15456
rect 49476 15447 49525 15453
rect 49476 15444 49482 15447
rect 50062 15444 50068 15456
rect 50120 15484 50126 15496
rect 50632 15493 50660 15524
rect 51810 15512 51816 15524
rect 51868 15512 51874 15564
rect 50525 15487 50583 15493
rect 50525 15484 50537 15487
rect 50120 15456 50537 15484
rect 50120 15444 50126 15456
rect 50525 15453 50537 15456
rect 50571 15453 50583 15487
rect 50525 15447 50583 15453
rect 50617 15487 50675 15493
rect 50617 15453 50629 15487
rect 50663 15453 50675 15487
rect 50617 15447 50675 15453
rect 50709 15487 50767 15493
rect 50709 15453 50721 15487
rect 50755 15453 50767 15487
rect 50709 15447 50767 15453
rect 48556 15388 49096 15416
rect 49344 15416 49372 15444
rect 49970 15416 49976 15428
rect 49344 15388 49976 15416
rect 48556 15376 48562 15388
rect 49970 15376 49976 15388
rect 50028 15376 50034 15428
rect 50724 15416 50752 15447
rect 50798 15444 50804 15496
rect 50856 15484 50862 15496
rect 50893 15487 50951 15493
rect 50893 15484 50905 15487
rect 50856 15456 50905 15484
rect 50856 15444 50862 15456
rect 50893 15453 50905 15456
rect 50939 15453 50951 15487
rect 50893 15447 50951 15453
rect 51626 15444 51632 15496
rect 51684 15444 51690 15496
rect 52104 15493 52132 15592
rect 52549 15589 52561 15592
rect 52595 15620 52607 15623
rect 52730 15620 52736 15632
rect 52595 15592 52736 15620
rect 52595 15589 52607 15592
rect 52549 15583 52607 15589
rect 52730 15580 52736 15592
rect 52788 15580 52794 15632
rect 51905 15487 51963 15493
rect 51905 15453 51917 15487
rect 51951 15453 51963 15487
rect 51905 15447 51963 15453
rect 52089 15487 52147 15493
rect 52089 15453 52101 15487
rect 52135 15453 52147 15487
rect 52089 15447 52147 15453
rect 52273 15487 52331 15493
rect 52273 15453 52285 15487
rect 52319 15484 52331 15487
rect 52822 15484 52828 15496
rect 52319 15456 52828 15484
rect 52319 15453 52331 15456
rect 52273 15447 52331 15453
rect 51074 15416 51080 15428
rect 50724 15388 51080 15416
rect 51074 15376 51080 15388
rect 51132 15376 51138 15428
rect 51920 15416 51948 15447
rect 52822 15444 52828 15456
rect 52880 15444 52886 15496
rect 52932 15416 52960 15648
rect 53098 15580 53104 15632
rect 53156 15620 53162 15632
rect 56502 15620 56508 15632
rect 53156 15592 56508 15620
rect 53156 15580 53162 15592
rect 56502 15580 56508 15592
rect 56560 15580 56566 15632
rect 54846 15512 54852 15564
rect 54904 15512 54910 15564
rect 55490 15552 55496 15564
rect 55324 15524 55496 15552
rect 53466 15444 53472 15496
rect 53524 15444 53530 15496
rect 53558 15444 53564 15496
rect 53616 15444 53622 15496
rect 51644 15388 52960 15416
rect 53484 15416 53512 15444
rect 53653 15419 53711 15425
rect 53653 15416 53665 15419
rect 53484 15388 53665 15416
rect 47486 15308 47492 15360
rect 47544 15308 47550 15360
rect 47578 15308 47584 15360
rect 47636 15348 47642 15360
rect 48038 15348 48044 15360
rect 47636 15320 48044 15348
rect 47636 15308 47642 15320
rect 48038 15308 48044 15320
rect 48096 15348 48102 15360
rect 48225 15351 48283 15357
rect 48225 15348 48237 15351
rect 48096 15320 48237 15348
rect 48096 15308 48102 15320
rect 48225 15317 48237 15320
rect 48271 15317 48283 15351
rect 48225 15311 48283 15317
rect 49510 15308 49516 15360
rect 49568 15348 49574 15360
rect 51644 15348 51672 15388
rect 53653 15385 53665 15388
rect 53699 15385 53711 15419
rect 53653 15379 53711 15385
rect 53837 15419 53895 15425
rect 53837 15385 53849 15419
rect 53883 15416 53895 15419
rect 54018 15416 54024 15428
rect 53883 15388 54024 15416
rect 53883 15385 53895 15388
rect 53837 15379 53895 15385
rect 54018 15376 54024 15388
rect 54076 15376 54082 15428
rect 54864 15416 54892 15512
rect 55324 15493 55352 15524
rect 55490 15512 55496 15524
rect 55548 15512 55554 15564
rect 55585 15555 55643 15561
rect 55585 15521 55597 15555
rect 55631 15552 55643 15555
rect 56612 15552 56640 15648
rect 56778 15580 56784 15632
rect 56836 15580 56842 15632
rect 56870 15580 56876 15632
rect 56928 15620 56934 15632
rect 57241 15623 57299 15629
rect 57241 15620 57253 15623
rect 56928 15592 57253 15620
rect 56928 15580 56934 15592
rect 57241 15589 57253 15592
rect 57287 15589 57299 15623
rect 57241 15583 57299 15589
rect 55631 15524 56640 15552
rect 55631 15521 55643 15524
rect 55585 15515 55643 15521
rect 56796 15493 56824 15580
rect 57716 15552 57744 15648
rect 57790 15580 57796 15632
rect 57848 15620 57854 15632
rect 57848 15592 58204 15620
rect 57848 15580 57854 15592
rect 57716 15524 57928 15552
rect 55309 15487 55367 15493
rect 55309 15453 55321 15487
rect 55355 15453 55367 15487
rect 55309 15447 55367 15453
rect 55401 15487 55459 15493
rect 55401 15453 55413 15487
rect 55447 15453 55459 15487
rect 56597 15487 56655 15493
rect 56597 15484 56609 15487
rect 55401 15447 55459 15453
rect 56336 15456 56609 15484
rect 55416 15416 55444 15447
rect 54864 15388 55444 15416
rect 56336 15360 56364 15456
rect 56597 15453 56609 15456
rect 56643 15453 56655 15487
rect 56597 15447 56655 15453
rect 56781 15487 56839 15493
rect 56781 15453 56793 15487
rect 56827 15453 56839 15487
rect 56781 15447 56839 15453
rect 57517 15487 57575 15493
rect 57517 15453 57529 15487
rect 57563 15453 57575 15487
rect 57517 15447 57575 15453
rect 56612 15416 56640 15447
rect 57532 15416 57560 15447
rect 57698 15444 57704 15496
rect 57756 15444 57762 15496
rect 57900 15493 57928 15524
rect 57885 15487 57943 15493
rect 57885 15453 57897 15487
rect 57931 15453 57943 15487
rect 57885 15447 57943 15453
rect 58066 15444 58072 15496
rect 58124 15444 58130 15496
rect 58176 15493 58204 15592
rect 58161 15487 58219 15493
rect 58161 15453 58173 15487
rect 58207 15453 58219 15487
rect 58161 15447 58219 15453
rect 58345 15487 58403 15493
rect 58345 15453 58357 15487
rect 58391 15484 58403 15487
rect 58391 15456 58572 15484
rect 58391 15453 58403 15456
rect 58345 15447 58403 15453
rect 56612 15388 57560 15416
rect 57609 15419 57667 15425
rect 57609 15385 57621 15419
rect 57655 15416 57667 15419
rect 58434 15416 58440 15428
rect 57655 15388 58440 15416
rect 57655 15385 57667 15388
rect 57609 15379 57667 15385
rect 58434 15376 58440 15388
rect 58492 15376 58498 15428
rect 49568 15320 51672 15348
rect 51721 15351 51779 15357
rect 49568 15308 49574 15320
rect 51721 15317 51733 15351
rect 51767 15348 51779 15351
rect 52181 15351 52239 15357
rect 52181 15348 52193 15351
rect 51767 15320 52193 15348
rect 51767 15317 51779 15320
rect 51721 15311 51779 15317
rect 52181 15317 52193 15320
rect 52227 15317 52239 15351
rect 52181 15311 52239 15317
rect 56318 15308 56324 15360
rect 56376 15308 56382 15360
rect 56505 15351 56563 15357
rect 56505 15317 56517 15351
rect 56551 15348 56563 15351
rect 56962 15348 56968 15360
rect 56551 15320 56968 15348
rect 56551 15317 56563 15320
rect 56505 15311 56563 15317
rect 56962 15308 56968 15320
rect 57020 15348 57026 15360
rect 57514 15348 57520 15360
rect 57020 15320 57520 15348
rect 57020 15308 57026 15320
rect 57514 15308 57520 15320
rect 57572 15308 57578 15360
rect 57698 15308 57704 15360
rect 57756 15348 57762 15360
rect 58544 15348 58572 15456
rect 57756 15320 58572 15348
rect 57756 15308 57762 15320
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 46566 15104 46572 15156
rect 46624 15104 46630 15156
rect 47857 15147 47915 15153
rect 47857 15113 47869 15147
rect 47903 15144 47915 15147
rect 48406 15144 48412 15156
rect 47903 15116 48412 15144
rect 47903 15113 47915 15116
rect 47857 15107 47915 15113
rect 48406 15104 48412 15116
rect 48464 15104 48470 15156
rect 49050 15104 49056 15156
rect 49108 15144 49114 15156
rect 49145 15147 49203 15153
rect 49145 15144 49157 15147
rect 49108 15116 49157 15144
rect 49108 15104 49114 15116
rect 49145 15113 49157 15116
rect 49191 15113 49203 15147
rect 49145 15107 49203 15113
rect 49234 15104 49240 15156
rect 49292 15104 49298 15156
rect 50062 15104 50068 15156
rect 50120 15104 50126 15156
rect 50154 15104 50160 15156
rect 50212 15144 50218 15156
rect 50341 15147 50399 15153
rect 50341 15144 50353 15147
rect 50212 15116 50353 15144
rect 50212 15104 50218 15116
rect 50341 15113 50353 15116
rect 50387 15113 50399 15147
rect 50341 15107 50399 15113
rect 50614 15104 50620 15156
rect 50672 15144 50678 15156
rect 50672 15116 51028 15144
rect 50672 15104 50678 15116
rect 50080 15076 50108 15104
rect 50430 15076 50436 15088
rect 46860 15048 48820 15076
rect 2685 15011 2743 15017
rect 2685 14977 2697 15011
rect 2731 15008 2743 15011
rect 10134 15008 10140 15020
rect 2731 14980 10140 15008
rect 2731 14977 2743 14980
rect 2685 14971 2743 14977
rect 10134 14968 10140 14980
rect 10192 14968 10198 15020
rect 46860 15017 46888 15048
rect 46845 15011 46903 15017
rect 46845 14977 46857 15011
rect 46891 14977 46903 15011
rect 46845 14971 46903 14977
rect 47578 14968 47584 15020
rect 47636 14968 47642 15020
rect 47673 15011 47731 15017
rect 47673 14977 47685 15011
rect 47719 15008 47731 15011
rect 47946 15008 47952 15020
rect 47719 14980 47952 15008
rect 47719 14977 47731 14980
rect 47673 14971 47731 14977
rect 47946 14968 47952 14980
rect 48004 15008 48010 15020
rect 48130 15008 48136 15020
rect 48004 14980 48136 15008
rect 48004 14968 48010 14980
rect 48130 14968 48136 14980
rect 48188 14968 48194 15020
rect 48332 15017 48360 15048
rect 48792 15020 48820 15048
rect 49252 15048 50436 15076
rect 48317 15011 48375 15017
rect 48317 14977 48329 15011
rect 48363 14977 48375 15011
rect 48317 14971 48375 14977
rect 48498 14968 48504 15020
rect 48556 14968 48562 15020
rect 48682 14968 48688 15020
rect 48740 14968 48746 15020
rect 48774 14968 48780 15020
rect 48832 14968 48838 15020
rect 49252 15017 49280 15048
rect 50430 15036 50436 15048
rect 50488 15076 50494 15088
rect 50488 15048 50936 15076
rect 50488 15036 50494 15048
rect 48869 15011 48927 15017
rect 48869 14977 48881 15011
rect 48915 15008 48927 15011
rect 49237 15011 49295 15017
rect 49237 15008 49249 15011
rect 48915 14980 49249 15008
rect 48915 14977 48927 14980
rect 48869 14971 48927 14977
rect 49237 14977 49249 14980
rect 49283 14977 49295 15011
rect 49237 14971 49295 14977
rect 49421 15011 49479 15017
rect 49421 14977 49433 15011
rect 49467 15008 49479 15011
rect 50062 15008 50068 15020
rect 49467 14980 50068 15008
rect 49467 14977 49479 14980
rect 49421 14971 49479 14977
rect 50062 14968 50068 14980
rect 50120 14968 50126 15020
rect 50522 15008 50528 15020
rect 50172 14980 50528 15008
rect 934 14900 940 14952
rect 992 14940 998 14952
rect 1581 14943 1639 14949
rect 1581 14940 1593 14943
rect 992 14912 1593 14940
rect 992 14900 998 14912
rect 1581 14909 1593 14912
rect 1627 14909 1639 14943
rect 1581 14903 1639 14909
rect 46569 14943 46627 14949
rect 46569 14909 46581 14943
rect 46615 14940 46627 14943
rect 47486 14940 47492 14952
rect 46615 14912 47492 14940
rect 46615 14909 46627 14912
rect 46569 14903 46627 14909
rect 47486 14900 47492 14912
rect 47544 14900 47550 14952
rect 47857 14943 47915 14949
rect 47857 14909 47869 14943
rect 47903 14940 47915 14943
rect 48225 14943 48283 14949
rect 48225 14940 48237 14943
rect 47903 14912 48237 14940
rect 47903 14909 47915 14912
rect 47857 14903 47915 14909
rect 48225 14909 48237 14912
rect 48271 14909 48283 14943
rect 48516 14940 48544 14968
rect 50172 14949 50200 14980
rect 50522 14968 50528 14980
rect 50580 14968 50586 15020
rect 50632 15017 50660 15048
rect 50617 15011 50675 15017
rect 50617 14977 50629 15011
rect 50663 14977 50675 15011
rect 50617 14971 50675 14977
rect 50706 14968 50712 15020
rect 50764 14968 50770 15020
rect 50801 15011 50859 15017
rect 50801 14977 50813 15011
rect 50847 14977 50859 15011
rect 50801 14971 50859 14977
rect 49697 14943 49755 14949
rect 49697 14940 49709 14943
rect 48516 14912 49709 14940
rect 48225 14903 48283 14909
rect 49697 14909 49709 14912
rect 49743 14940 49755 14943
rect 50157 14943 50215 14949
rect 50157 14940 50169 14943
rect 49743 14912 50169 14940
rect 49743 14909 49755 14912
rect 49697 14903 49755 14909
rect 50157 14909 50169 14912
rect 50203 14909 50215 14943
rect 50816 14940 50844 14971
rect 50157 14903 50215 14909
rect 50540 14912 50844 14940
rect 50908 14940 50936 15048
rect 51000 15017 51028 15116
rect 51074 15104 51080 15156
rect 51132 15104 51138 15156
rect 51537 15147 51595 15153
rect 51537 15113 51549 15147
rect 51583 15144 51595 15147
rect 51626 15144 51632 15156
rect 51583 15116 51632 15144
rect 51583 15113 51595 15116
rect 51537 15107 51595 15113
rect 51626 15104 51632 15116
rect 51684 15104 51690 15156
rect 52822 15104 52828 15156
rect 52880 15104 52886 15156
rect 53006 15104 53012 15156
rect 53064 15104 53070 15156
rect 53190 15104 53196 15156
rect 53248 15104 53254 15156
rect 53558 15104 53564 15156
rect 53616 15104 53622 15156
rect 53650 15104 53656 15156
rect 53708 15104 53714 15156
rect 54018 15104 54024 15156
rect 54076 15104 54082 15156
rect 56873 15147 56931 15153
rect 56873 15113 56885 15147
rect 56919 15144 56931 15147
rect 56962 15144 56968 15156
rect 56919 15116 56968 15144
rect 56919 15113 56931 15116
rect 56873 15107 56931 15113
rect 56962 15104 56968 15116
rect 57020 15104 57026 15156
rect 57698 15104 57704 15156
rect 57756 15104 57762 15156
rect 53024 15076 53052 15104
rect 51092 15048 53052 15076
rect 51092 15017 51120 15048
rect 50985 15011 51043 15017
rect 50985 14977 50997 15011
rect 51031 14977 51043 15011
rect 50985 14971 51043 14977
rect 51077 15011 51135 15017
rect 51077 14977 51089 15011
rect 51123 14977 51135 15011
rect 51077 14971 51135 14977
rect 51261 15011 51319 15017
rect 51261 14977 51273 15011
rect 51307 14977 51319 15011
rect 51261 14971 51319 14977
rect 51092 14940 51120 14971
rect 50908 14912 51120 14940
rect 46753 14875 46811 14881
rect 46753 14841 46765 14875
rect 46799 14872 46811 14875
rect 47118 14872 47124 14884
rect 46799 14844 47124 14872
rect 46799 14841 46811 14844
rect 46753 14835 46811 14841
rect 47118 14832 47124 14844
rect 47176 14832 47182 14884
rect 50540 14816 50568 14912
rect 51276 14872 51304 14971
rect 51442 14968 51448 15020
rect 51500 14968 51506 15020
rect 51644 15017 51672 15048
rect 51629 15011 51687 15017
rect 51629 14977 51641 15011
rect 51675 14977 51687 15011
rect 51629 14971 51687 14977
rect 52730 14968 52736 15020
rect 52788 14968 52794 15020
rect 52914 14968 52920 15020
rect 52972 14968 52978 15020
rect 53024 15017 53052 15048
rect 53374 15036 53380 15088
rect 53432 15036 53438 15088
rect 53668 15076 53696 15104
rect 53668 15048 54064 15076
rect 53009 15011 53067 15017
rect 53009 14977 53021 15011
rect 53055 14977 53067 15011
rect 53009 14971 53067 14977
rect 53193 15011 53251 15017
rect 53193 14977 53205 15011
rect 53239 14977 53251 15011
rect 53392 15008 53420 15036
rect 53561 15011 53619 15017
rect 53561 15008 53573 15011
rect 53392 14980 53573 15008
rect 53193 14971 53251 14977
rect 53561 14977 53573 14980
rect 53607 14977 53619 15011
rect 53561 14971 53619 14977
rect 53745 15011 53803 15017
rect 53745 14977 53757 15011
rect 53791 15008 53803 15011
rect 53926 15008 53932 15020
rect 53791 14980 53932 15008
rect 53791 14977 53803 14980
rect 53745 14971 53803 14977
rect 53208 14940 53236 14971
rect 53926 14968 53932 14980
rect 53984 14968 53990 15020
rect 54036 15017 54064 15048
rect 54110 15036 54116 15088
rect 54168 15036 54174 15088
rect 54021 15011 54079 15017
rect 54021 14977 54033 15011
rect 54067 14977 54079 15011
rect 54021 14971 54079 14977
rect 54297 15011 54355 15017
rect 54297 14977 54309 15011
rect 54343 15008 54355 15011
rect 55582 15008 55588 15020
rect 54343 14980 55588 15008
rect 54343 14977 54355 14980
rect 54297 14971 54355 14977
rect 55582 14968 55588 14980
rect 55640 14968 55646 15020
rect 58434 14968 58440 15020
rect 58492 14968 58498 15020
rect 53834 14940 53840 14952
rect 53208 14912 53840 14940
rect 53834 14900 53840 14912
rect 53892 14900 53898 14952
rect 56134 14900 56140 14952
rect 56192 14900 56198 14952
rect 57146 14900 57152 14952
rect 57204 14900 57210 14952
rect 54018 14872 54024 14884
rect 51276 14844 54024 14872
rect 54018 14832 54024 14844
rect 54076 14832 54082 14884
rect 50522 14764 50528 14816
rect 50580 14764 50586 14816
rect 55490 14764 55496 14816
rect 55548 14764 55554 14816
rect 57882 14764 57888 14816
rect 57940 14764 57946 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 48409 14603 48467 14609
rect 48409 14569 48421 14603
rect 48455 14600 48467 14603
rect 48498 14600 48504 14612
rect 48455 14572 48504 14600
rect 48455 14569 48467 14572
rect 48409 14563 48467 14569
rect 48498 14560 48504 14572
rect 48556 14560 48562 14612
rect 48593 14603 48651 14609
rect 48593 14569 48605 14603
rect 48639 14600 48651 14603
rect 48682 14600 48688 14612
rect 48639 14572 48688 14600
rect 48639 14569 48651 14572
rect 48593 14563 48651 14569
rect 48682 14560 48688 14572
rect 48740 14560 48746 14612
rect 49142 14560 49148 14612
rect 49200 14600 49206 14612
rect 49237 14603 49295 14609
rect 49237 14600 49249 14603
rect 49200 14572 49249 14600
rect 49200 14560 49206 14572
rect 49237 14569 49249 14572
rect 49283 14569 49295 14603
rect 49237 14563 49295 14569
rect 50522 14560 50528 14612
rect 50580 14560 50586 14612
rect 50614 14560 50620 14612
rect 50672 14560 50678 14612
rect 50706 14560 50712 14612
rect 50764 14600 50770 14612
rect 52365 14603 52423 14609
rect 50764 14572 51074 14600
rect 50764 14560 50770 14572
rect 50632 14532 50660 14560
rect 50893 14535 50951 14541
rect 50893 14532 50905 14535
rect 50632 14504 50905 14532
rect 50893 14501 50905 14504
rect 50939 14501 50951 14535
rect 50893 14495 50951 14501
rect 51046 14464 51074 14572
rect 52365 14569 52377 14603
rect 52411 14600 52423 14603
rect 52730 14600 52736 14612
rect 52411 14572 52736 14600
rect 52411 14569 52423 14572
rect 52365 14563 52423 14569
rect 52730 14560 52736 14572
rect 52788 14560 52794 14612
rect 57146 14560 57152 14612
rect 57204 14600 57210 14612
rect 58253 14603 58311 14609
rect 58253 14600 58265 14603
rect 57204 14572 58265 14600
rect 57204 14560 57210 14572
rect 58253 14569 58265 14572
rect 58299 14569 58311 14603
rect 58253 14563 58311 14569
rect 58894 14560 58900 14612
rect 58952 14560 58958 14612
rect 56686 14492 56692 14544
rect 56744 14492 56750 14544
rect 58066 14492 58072 14544
rect 58124 14532 58130 14544
rect 58345 14535 58403 14541
rect 58345 14532 58357 14535
rect 58124 14504 58357 14532
rect 58124 14492 58130 14504
rect 58345 14501 58357 14504
rect 58391 14501 58403 14535
rect 58345 14495 58403 14501
rect 51046 14436 52316 14464
rect 52288 14408 52316 14436
rect 48501 14399 48559 14405
rect 48501 14365 48513 14399
rect 48547 14365 48559 14399
rect 48501 14359 48559 14365
rect 48685 14399 48743 14405
rect 48685 14365 48697 14399
rect 48731 14396 48743 14399
rect 49145 14399 49203 14405
rect 49145 14396 49157 14399
rect 48731 14368 49157 14396
rect 48731 14365 48743 14368
rect 48685 14359 48743 14365
rect 49145 14365 49157 14368
rect 49191 14365 49203 14399
rect 49145 14359 49203 14365
rect 48516 14272 48544 14359
rect 49160 14328 49188 14359
rect 49326 14356 49332 14408
rect 49384 14356 49390 14408
rect 50430 14356 50436 14408
rect 50488 14356 50494 14408
rect 50617 14399 50675 14405
rect 50617 14365 50629 14399
rect 50663 14396 50675 14399
rect 50663 14368 52132 14396
rect 50663 14365 50675 14368
rect 50617 14359 50675 14365
rect 50448 14328 50476 14356
rect 49160 14300 50476 14328
rect 52104 14272 52132 14368
rect 52270 14356 52276 14408
rect 52328 14356 52334 14408
rect 52457 14399 52515 14405
rect 52457 14365 52469 14399
rect 52503 14396 52515 14399
rect 53374 14396 53380 14408
rect 52503 14368 53380 14396
rect 52503 14365 52515 14368
rect 52457 14359 52515 14365
rect 53374 14356 53380 14368
rect 53432 14356 53438 14408
rect 53926 14356 53932 14408
rect 53984 14396 53990 14408
rect 55125 14399 55183 14405
rect 55125 14396 55137 14399
rect 53984 14368 55137 14396
rect 53984 14356 53990 14368
rect 55125 14365 55137 14368
rect 55171 14365 55183 14399
rect 55125 14359 55183 14365
rect 48498 14220 48504 14272
rect 48556 14220 48562 14272
rect 52086 14220 52092 14272
rect 52144 14220 52150 14272
rect 54018 14220 54024 14272
rect 54076 14260 54082 14272
rect 54754 14260 54760 14272
rect 54076 14232 54760 14260
rect 54076 14220 54082 14232
rect 54754 14220 54760 14232
rect 54812 14220 54818 14272
rect 55030 14220 55036 14272
rect 55088 14220 55094 14272
rect 55140 14260 55168 14359
rect 55306 14356 55312 14408
rect 55364 14396 55370 14408
rect 56873 14399 56931 14405
rect 56873 14396 56885 14399
rect 55364 14368 56885 14396
rect 55364 14356 55370 14368
rect 56873 14365 56885 14368
rect 56919 14365 56931 14399
rect 56873 14359 56931 14365
rect 58529 14399 58587 14405
rect 58529 14365 58541 14399
rect 58575 14396 58587 14399
rect 58912 14396 58940 14560
rect 58575 14368 58940 14396
rect 58575 14365 58587 14368
rect 58529 14359 58587 14365
rect 55214 14288 55220 14340
rect 55272 14328 55278 14340
rect 55554 14331 55612 14337
rect 55554 14328 55566 14331
rect 55272 14300 55566 14328
rect 55272 14288 55278 14300
rect 55554 14297 55566 14300
rect 55600 14297 55612 14331
rect 55554 14291 55612 14297
rect 55692 14300 56732 14328
rect 55692 14260 55720 14300
rect 55140 14232 55720 14260
rect 56704 14260 56732 14300
rect 56778 14288 56784 14340
rect 56836 14328 56842 14340
rect 57118 14331 57176 14337
rect 57118 14328 57130 14331
rect 56836 14300 57130 14328
rect 56836 14288 56842 14300
rect 57118 14297 57130 14300
rect 57164 14297 57176 14331
rect 57118 14291 57176 14297
rect 58158 14260 58164 14272
rect 56704 14232 58164 14260
rect 58158 14220 58164 14232
rect 58216 14220 58222 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 47857 14059 47915 14065
rect 47857 14025 47869 14059
rect 47903 14056 47915 14059
rect 48314 14056 48320 14068
rect 47903 14028 48320 14056
rect 47903 14025 47915 14028
rect 47857 14019 47915 14025
rect 48314 14016 48320 14028
rect 48372 14016 48378 14068
rect 49326 14016 49332 14068
rect 49384 14016 49390 14068
rect 51261 14059 51319 14065
rect 51261 14025 51273 14059
rect 51307 14025 51319 14059
rect 51261 14019 51319 14025
rect 51276 13988 51304 14019
rect 51442 14016 51448 14068
rect 51500 14016 51506 14068
rect 52733 14059 52791 14065
rect 52733 14025 52745 14059
rect 52779 14056 52791 14059
rect 52914 14056 52920 14068
rect 52779 14028 52920 14056
rect 52779 14025 52791 14028
rect 52733 14019 52791 14025
rect 52914 14016 52920 14028
rect 52972 14016 52978 14068
rect 53006 14016 53012 14068
rect 53064 14056 53070 14068
rect 53650 14056 53656 14068
rect 53064 14028 53656 14056
rect 53064 14016 53070 14028
rect 53650 14016 53656 14028
rect 53708 14016 53714 14068
rect 53834 14016 53840 14068
rect 53892 14056 53898 14068
rect 54205 14059 54263 14065
rect 54205 14056 54217 14059
rect 53892 14028 54217 14056
rect 53892 14016 53898 14028
rect 54205 14025 54217 14028
rect 54251 14025 54263 14059
rect 54205 14019 54263 14025
rect 55030 14016 55036 14068
rect 55088 14016 55094 14068
rect 55125 14059 55183 14065
rect 55125 14025 55137 14059
rect 55171 14056 55183 14059
rect 55214 14056 55220 14068
rect 55171 14028 55220 14056
rect 55171 14025 55183 14028
rect 55125 14019 55183 14025
rect 55214 14016 55220 14028
rect 55272 14016 55278 14068
rect 55490 14016 55496 14068
rect 55548 14016 55554 14068
rect 55582 14016 55588 14068
rect 55640 14016 55646 14068
rect 56134 14016 56140 14068
rect 56192 14056 56198 14068
rect 56321 14059 56379 14065
rect 56321 14056 56333 14059
rect 56192 14028 56333 14056
rect 56192 14016 56198 14028
rect 56321 14025 56333 14028
rect 56367 14025 56379 14059
rect 56321 14019 56379 14025
rect 56686 14016 56692 14068
rect 56744 14016 56750 14068
rect 56778 14016 56784 14068
rect 56836 14016 56842 14068
rect 58066 14016 58072 14068
rect 58124 14016 58130 14068
rect 58158 14016 58164 14068
rect 58216 14056 58222 14068
rect 58345 14059 58403 14065
rect 58345 14056 58357 14059
rect 58216 14028 58357 14056
rect 58216 14016 58222 14028
rect 58345 14025 58357 14028
rect 58391 14025 58403 14059
rect 58345 14019 58403 14025
rect 58894 14016 58900 14068
rect 58952 14016 58958 14068
rect 53668 13988 53696 14016
rect 47136 13960 48176 13988
rect 51276 13960 51402 13988
rect 47136 13932 47164 13960
rect 47118 13880 47124 13932
rect 47176 13880 47182 13932
rect 47578 13880 47584 13932
rect 47636 13880 47642 13932
rect 47673 13923 47731 13929
rect 47673 13889 47685 13923
rect 47719 13920 47731 13923
rect 47946 13920 47952 13932
rect 47719 13892 47952 13920
rect 47719 13889 47731 13892
rect 47673 13883 47731 13889
rect 47780 13784 47808 13892
rect 47946 13880 47952 13892
rect 48004 13880 48010 13932
rect 48148 13929 48176 13960
rect 48133 13923 48191 13929
rect 48133 13889 48145 13923
rect 48179 13920 48191 13923
rect 48317 13923 48375 13929
rect 48317 13920 48329 13923
rect 48179 13892 48329 13920
rect 48179 13889 48191 13892
rect 48133 13883 48191 13889
rect 48317 13889 48329 13892
rect 48363 13889 48375 13923
rect 48317 13883 48375 13889
rect 48409 13923 48467 13929
rect 48409 13889 48421 13923
rect 48455 13889 48467 13923
rect 48409 13883 48467 13889
rect 49053 13923 49111 13929
rect 49053 13889 49065 13923
rect 49099 13920 49111 13923
rect 49878 13920 49884 13932
rect 49099 13892 49884 13920
rect 49099 13889 49111 13892
rect 49053 13883 49111 13889
rect 47857 13855 47915 13861
rect 47857 13821 47869 13855
rect 47903 13852 47915 13855
rect 48041 13855 48099 13861
rect 48041 13852 48053 13855
rect 47903 13824 48053 13852
rect 47903 13821 47915 13824
rect 47857 13815 47915 13821
rect 48041 13821 48053 13824
rect 48087 13821 48099 13855
rect 48424 13852 48452 13883
rect 49878 13880 49884 13892
rect 49936 13880 49942 13932
rect 50985 13923 51043 13929
rect 50985 13889 50997 13923
rect 51031 13889 51043 13923
rect 50985 13883 51043 13889
rect 51169 13923 51227 13929
rect 51169 13889 51181 13923
rect 51215 13889 51227 13923
rect 51169 13883 51227 13889
rect 48498 13852 48504 13864
rect 48424 13824 48504 13852
rect 48041 13815 48099 13821
rect 48498 13812 48504 13824
rect 48556 13852 48562 13864
rect 49234 13852 49240 13864
rect 48556 13824 49240 13852
rect 48556 13812 48562 13824
rect 49234 13812 49240 13824
rect 49292 13812 49298 13864
rect 49326 13812 49332 13864
rect 49384 13812 49390 13864
rect 49142 13784 49148 13796
rect 47780 13756 49148 13784
rect 49142 13744 49148 13756
rect 49200 13744 49206 13796
rect 51000 13784 51028 13883
rect 51184 13852 51212 13883
rect 51258 13880 51264 13932
rect 51316 13880 51322 13932
rect 51374 13929 51402 13960
rect 51460 13960 52868 13988
rect 51460 13932 51488 13960
rect 52840 13942 52868 13960
rect 53004 13960 53236 13988
rect 53668 13960 54156 13988
rect 52917 13945 52975 13951
rect 52917 13942 52929 13945
rect 51353 13923 51411 13929
rect 51353 13889 51365 13923
rect 51399 13889 51411 13923
rect 51353 13883 51411 13889
rect 51442 13880 51448 13932
rect 51500 13880 51506 13932
rect 51534 13880 51540 13932
rect 51592 13880 51598 13932
rect 51810 13880 51816 13932
rect 51868 13880 51874 13932
rect 52840 13914 52929 13942
rect 51721 13855 51779 13861
rect 51721 13852 51733 13855
rect 51184 13824 51733 13852
rect 51721 13821 51733 13824
rect 51767 13821 51779 13855
rect 52840 13852 52868 13914
rect 52917 13911 52929 13914
rect 52963 13911 52975 13945
rect 52917 13905 52975 13911
rect 53004 13929 53032 13960
rect 53004 13923 53067 13929
rect 53004 13898 53021 13923
rect 53009 13889 53021 13898
rect 53055 13889 53067 13923
rect 53009 13883 53067 13889
rect 53098 13880 53104 13932
rect 53156 13880 53162 13932
rect 53208 13920 53236 13960
rect 53837 13923 53895 13929
rect 53837 13920 53849 13923
rect 53208 13892 53849 13920
rect 52914 13852 52920 13864
rect 52840 13824 52920 13852
rect 51721 13815 51779 13821
rect 52914 13812 52920 13824
rect 52972 13812 52978 13864
rect 53208 13852 53236 13892
rect 53837 13889 53849 13892
rect 53883 13920 53895 13923
rect 53926 13920 53932 13932
rect 53883 13892 53932 13920
rect 53883 13889 53895 13892
rect 53837 13883 53895 13889
rect 53926 13880 53932 13892
rect 53984 13880 53990 13932
rect 54018 13880 54024 13932
rect 54076 13880 54082 13932
rect 54128 13929 54156 13960
rect 54113 13923 54171 13929
rect 54113 13889 54125 13923
rect 54159 13889 54171 13923
rect 54113 13883 54171 13889
rect 54205 13923 54263 13929
rect 54205 13889 54217 13923
rect 54251 13889 54263 13923
rect 54389 13923 54447 13929
rect 54389 13920 54401 13923
rect 54205 13883 54263 13889
rect 54312 13892 54401 13920
rect 54220 13852 54248 13883
rect 53116 13844 53236 13852
rect 53024 13824 53236 13844
rect 53852 13824 54248 13852
rect 53024 13816 53144 13824
rect 53024 13784 53052 13816
rect 51000 13756 53052 13784
rect 53852 13728 53880 13824
rect 54113 13787 54171 13793
rect 54113 13753 54125 13787
rect 54159 13784 54171 13787
rect 54312 13784 54340 13892
rect 54389 13889 54401 13892
rect 54435 13889 54447 13923
rect 54389 13883 54447 13889
rect 54849 13923 54907 13929
rect 54849 13889 54861 13923
rect 54895 13920 54907 13923
rect 55048 13920 55076 14016
rect 54895 13892 55076 13920
rect 54895 13889 54907 13892
rect 54849 13883 54907 13889
rect 55125 13855 55183 13861
rect 55125 13821 55137 13855
rect 55171 13852 55183 13855
rect 55508 13852 55536 14016
rect 55171 13824 55536 13852
rect 55600 13852 55628 14016
rect 56704 13988 56732 14016
rect 56152 13960 56732 13988
rect 58084 13988 58112 14016
rect 58084 13960 58296 13988
rect 56152 13929 56180 13960
rect 58268 13929 58296 13960
rect 56137 13923 56195 13929
rect 56137 13889 56149 13923
rect 56183 13889 56195 13923
rect 56137 13883 56195 13889
rect 56229 13923 56287 13929
rect 56229 13889 56241 13923
rect 56275 13889 56287 13923
rect 56413 13923 56471 13929
rect 56413 13920 56425 13923
rect 56229 13883 56287 13889
rect 56336 13892 56425 13920
rect 56244 13852 56272 13883
rect 56336 13864 56364 13892
rect 56413 13889 56425 13892
rect 56459 13889 56471 13923
rect 56413 13883 56471 13889
rect 56505 13923 56563 13929
rect 56505 13889 56517 13923
rect 56551 13920 56563 13923
rect 58161 13923 58219 13929
rect 58161 13920 58173 13923
rect 56551 13892 58173 13920
rect 56551 13889 56563 13892
rect 56505 13883 56563 13889
rect 58161 13889 58173 13892
rect 58207 13889 58219 13923
rect 58161 13883 58219 13889
rect 58253 13923 58311 13929
rect 58253 13889 58265 13923
rect 58299 13889 58311 13923
rect 58253 13883 58311 13889
rect 58529 13923 58587 13929
rect 58529 13889 58541 13923
rect 58575 13920 58587 13923
rect 58912 13920 58940 14016
rect 58575 13892 58940 13920
rect 58575 13889 58587 13892
rect 58529 13883 58587 13889
rect 55600 13824 56272 13852
rect 55171 13821 55183 13824
rect 55125 13815 55183 13821
rect 54159 13756 54340 13784
rect 54159 13753 54171 13756
rect 54113 13747 54171 13753
rect 54754 13744 54760 13796
rect 54812 13784 54818 13796
rect 55493 13787 55551 13793
rect 54812 13756 55444 13784
rect 54812 13744 54818 13756
rect 53834 13676 53840 13728
rect 53892 13676 53898 13728
rect 54846 13676 54852 13728
rect 54904 13716 54910 13728
rect 54941 13719 54999 13725
rect 54941 13716 54953 13719
rect 54904 13688 54953 13716
rect 54904 13676 54910 13688
rect 54941 13685 54953 13688
rect 54987 13685 54999 13719
rect 55416 13716 55444 13756
rect 55493 13753 55505 13787
rect 55539 13784 55551 13787
rect 55600 13784 55628 13824
rect 56318 13812 56324 13864
rect 56376 13812 56382 13864
rect 56781 13855 56839 13861
rect 56781 13821 56793 13855
rect 56827 13852 56839 13855
rect 57882 13852 57888 13864
rect 56827 13824 57888 13852
rect 56827 13821 56839 13824
rect 56781 13815 56839 13821
rect 57882 13812 57888 13824
rect 57940 13812 57946 13864
rect 57974 13784 57980 13796
rect 55539 13756 55628 13784
rect 56520 13756 57980 13784
rect 55539 13753 55551 13756
rect 55493 13747 55551 13753
rect 56520 13716 56548 13756
rect 57974 13744 57980 13756
rect 58032 13744 58038 13796
rect 55416 13688 56548 13716
rect 54941 13679 54999 13685
rect 56594 13676 56600 13728
rect 56652 13676 56658 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 47578 13472 47584 13524
rect 47636 13512 47642 13524
rect 47946 13512 47952 13524
rect 47636 13484 47952 13512
rect 47636 13472 47642 13484
rect 47946 13472 47952 13484
rect 48004 13512 48010 13524
rect 48501 13515 48559 13521
rect 48501 13512 48513 13515
rect 48004 13484 48513 13512
rect 48004 13472 48010 13484
rect 48501 13481 48513 13484
rect 48547 13481 48559 13515
rect 48501 13475 48559 13481
rect 49326 13472 49332 13524
rect 49384 13512 49390 13524
rect 49421 13515 49479 13521
rect 49421 13512 49433 13515
rect 49384 13484 49433 13512
rect 49384 13472 49390 13484
rect 49421 13481 49433 13484
rect 49467 13481 49479 13515
rect 49421 13475 49479 13481
rect 51534 13472 51540 13524
rect 51592 13512 51598 13524
rect 51721 13515 51779 13521
rect 51721 13512 51733 13515
rect 51592 13484 51733 13512
rect 51592 13472 51598 13484
rect 51721 13481 51733 13484
rect 51767 13481 51779 13515
rect 51721 13475 51779 13481
rect 53834 13472 53840 13524
rect 53892 13472 53898 13524
rect 54018 13472 54024 13524
rect 54076 13512 54082 13524
rect 54573 13515 54631 13521
rect 54573 13512 54585 13515
rect 54076 13484 54585 13512
rect 54076 13472 54082 13484
rect 54573 13481 54585 13484
rect 54619 13481 54631 13515
rect 54573 13475 54631 13481
rect 54846 13472 54852 13524
rect 54904 13512 54910 13524
rect 56413 13515 56471 13521
rect 56413 13512 56425 13515
rect 54904 13484 56425 13512
rect 54904 13472 54910 13484
rect 56413 13481 56425 13484
rect 56459 13512 56471 13515
rect 56594 13512 56600 13524
rect 56459 13484 56600 13512
rect 56459 13481 56471 13484
rect 56413 13475 56471 13481
rect 56594 13472 56600 13484
rect 56652 13472 56658 13524
rect 58342 13512 58348 13524
rect 56980 13484 58348 13512
rect 47673 13447 47731 13453
rect 47673 13413 47685 13447
rect 47719 13444 47731 13447
rect 47719 13416 49096 13444
rect 47719 13413 47731 13416
rect 47673 13407 47731 13413
rect 45922 13336 45928 13388
rect 45980 13376 45986 13388
rect 46290 13376 46296 13388
rect 45980 13348 46296 13376
rect 45980 13336 45986 13348
rect 46290 13336 46296 13348
rect 46348 13336 46354 13388
rect 49068 13385 49096 13416
rect 49970 13404 49976 13456
rect 50028 13444 50034 13456
rect 50028 13416 53512 13444
rect 50028 13404 50034 13416
rect 49053 13379 49111 13385
rect 49053 13345 49065 13379
rect 49099 13345 49111 13379
rect 53484 13376 53512 13416
rect 56042 13404 56048 13456
rect 56100 13404 56106 13456
rect 56060 13376 56088 13404
rect 49053 13339 49111 13345
rect 49344 13348 53420 13376
rect 53484 13348 56088 13376
rect 2777 13311 2835 13317
rect 2777 13277 2789 13311
rect 2823 13308 2835 13311
rect 6730 13308 6736 13320
rect 2823 13280 6736 13308
rect 2823 13277 2835 13280
rect 2777 13271 2835 13277
rect 6730 13268 6736 13280
rect 6788 13268 6794 13320
rect 48314 13268 48320 13320
rect 48372 13268 48378 13320
rect 49142 13268 49148 13320
rect 49200 13308 49206 13320
rect 49344 13317 49372 13348
rect 49329 13311 49387 13317
rect 49329 13308 49341 13311
rect 49200 13280 49341 13308
rect 49200 13268 49206 13280
rect 49329 13277 49341 13280
rect 49375 13277 49387 13311
rect 49329 13271 49387 13277
rect 49513 13311 49571 13317
rect 49513 13277 49525 13311
rect 49559 13308 49571 13311
rect 49559 13280 50016 13308
rect 49559 13277 49571 13280
rect 49513 13271 49571 13277
rect 934 13200 940 13252
rect 992 13240 998 13252
rect 1581 13243 1639 13249
rect 1581 13240 1593 13243
rect 992 13212 1593 13240
rect 992 13200 998 13212
rect 1581 13209 1593 13212
rect 1627 13209 1639 13243
rect 1581 13203 1639 13209
rect 46560 13243 46618 13249
rect 46560 13209 46572 13243
rect 46606 13240 46618 13243
rect 46842 13240 46848 13252
rect 46606 13212 46848 13240
rect 46606 13209 46618 13212
rect 46560 13203 46618 13209
rect 46842 13200 46848 13212
rect 46900 13200 46906 13252
rect 49988 13184 50016 13280
rect 51442 13268 51448 13320
rect 51500 13268 51506 13320
rect 51644 13317 51672 13348
rect 53392 13320 53420 13348
rect 56594 13336 56600 13388
rect 56652 13336 56658 13388
rect 51629 13311 51687 13317
rect 51629 13277 51641 13311
rect 51675 13277 51687 13311
rect 51629 13271 51687 13277
rect 51813 13311 51871 13317
rect 51813 13277 51825 13311
rect 51859 13277 51871 13311
rect 51813 13271 51871 13277
rect 51828 13240 51856 13271
rect 52086 13268 52092 13320
rect 52144 13268 52150 13320
rect 52178 13268 52184 13320
rect 52236 13268 52242 13320
rect 53374 13268 53380 13320
rect 53432 13268 53438 13320
rect 53558 13268 53564 13320
rect 53616 13268 53622 13320
rect 53745 13311 53803 13317
rect 53745 13277 53757 13311
rect 53791 13277 53803 13311
rect 53745 13271 53803 13277
rect 51997 13243 52055 13249
rect 51997 13240 52009 13243
rect 50724 13212 52009 13240
rect 50724 13184 50752 13212
rect 51997 13209 52009 13212
rect 52043 13209 52055 13243
rect 52104 13240 52132 13268
rect 53392 13240 53420 13268
rect 53760 13240 53788 13271
rect 53926 13268 53932 13320
rect 53984 13268 53990 13320
rect 54665 13311 54723 13317
rect 54665 13277 54677 13311
rect 54711 13308 54723 13311
rect 55950 13308 55956 13320
rect 54711 13280 55956 13308
rect 54711 13277 54723 13280
rect 54665 13271 54723 13277
rect 55950 13268 55956 13280
rect 56008 13268 56014 13320
rect 56980 13317 57008 13484
rect 58342 13472 58348 13484
rect 58400 13472 58406 13524
rect 57885 13447 57943 13453
rect 57885 13413 57897 13447
rect 57931 13413 57943 13447
rect 57885 13407 57943 13413
rect 56321 13311 56379 13317
rect 56321 13277 56333 13311
rect 56367 13277 56379 13311
rect 56321 13271 56379 13277
rect 56965 13311 57023 13317
rect 56965 13277 56977 13311
rect 57011 13277 57023 13311
rect 56965 13271 57023 13277
rect 57793 13311 57851 13317
rect 57793 13277 57805 13311
rect 57839 13308 57851 13311
rect 57900 13308 57928 13407
rect 57839 13280 57928 13308
rect 58069 13311 58127 13317
rect 57839 13277 57851 13280
rect 57793 13271 57851 13277
rect 58069 13277 58081 13311
rect 58115 13277 58127 13311
rect 58069 13271 58127 13277
rect 58529 13311 58587 13317
rect 58529 13277 58541 13311
rect 58575 13308 58587 13311
rect 58894 13308 58900 13320
rect 58575 13280 58900 13308
rect 58575 13277 58587 13280
rect 58529 13271 58587 13277
rect 52104 13212 53052 13240
rect 53392 13212 53788 13240
rect 51997 13203 52055 13209
rect 47762 13132 47768 13184
rect 47820 13132 47826 13184
rect 49970 13132 49976 13184
rect 50028 13132 50034 13184
rect 50706 13132 50712 13184
rect 50764 13132 50770 13184
rect 50890 13132 50896 13184
rect 50948 13132 50954 13184
rect 52638 13132 52644 13184
rect 52696 13172 52702 13184
rect 52825 13175 52883 13181
rect 52825 13172 52837 13175
rect 52696 13144 52837 13172
rect 52696 13132 52702 13144
rect 52825 13141 52837 13144
rect 52871 13141 52883 13175
rect 52825 13135 52883 13141
rect 52914 13132 52920 13184
rect 52972 13132 52978 13184
rect 53024 13172 53052 13212
rect 54202 13200 54208 13252
rect 54260 13200 54266 13252
rect 56336 13240 56364 13271
rect 56873 13243 56931 13249
rect 56873 13240 56885 13243
rect 56336 13212 56885 13240
rect 56873 13209 56885 13212
rect 56919 13209 56931 13243
rect 58084 13240 58112 13271
rect 58894 13268 58900 13280
rect 58952 13268 58958 13320
rect 58084 13212 58756 13240
rect 56873 13203 56931 13209
rect 54220 13172 54248 13200
rect 58728 13184 58756 13212
rect 53024 13144 54248 13172
rect 56502 13132 56508 13184
rect 56560 13172 56566 13184
rect 56597 13175 56655 13181
rect 56597 13172 56609 13175
rect 56560 13144 56609 13172
rect 56560 13132 56566 13144
rect 56597 13141 56609 13144
rect 56643 13141 56655 13175
rect 56597 13135 56655 13141
rect 56686 13132 56692 13184
rect 56744 13172 56750 13184
rect 57701 13175 57759 13181
rect 57701 13172 57713 13175
rect 56744 13144 57713 13172
rect 56744 13132 56750 13144
rect 57701 13141 57713 13144
rect 57747 13141 57759 13175
rect 57701 13135 57759 13141
rect 58710 13132 58716 13184
rect 58768 13132 58774 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 46842 12928 46848 12980
rect 46900 12928 46906 12980
rect 47762 12928 47768 12980
rect 47820 12928 47826 12980
rect 47857 12971 47915 12977
rect 47857 12937 47869 12971
rect 47903 12968 47915 12971
rect 48314 12968 48320 12980
rect 47903 12940 48320 12968
rect 47903 12937 47915 12940
rect 47857 12931 47915 12937
rect 48314 12928 48320 12940
rect 48372 12928 48378 12980
rect 49970 12928 49976 12980
rect 50028 12928 50034 12980
rect 50890 12928 50896 12980
rect 50948 12928 50954 12980
rect 51169 12971 51227 12977
rect 51169 12937 51181 12971
rect 51215 12968 51227 12971
rect 51442 12968 51448 12980
rect 51215 12940 51448 12968
rect 51215 12937 51227 12940
rect 51169 12931 51227 12937
rect 51442 12928 51448 12940
rect 51500 12928 51506 12980
rect 51810 12928 51816 12980
rect 51868 12968 51874 12980
rect 52089 12971 52147 12977
rect 52089 12968 52101 12971
rect 51868 12940 52101 12968
rect 51868 12928 51874 12940
rect 52089 12937 52101 12940
rect 52135 12937 52147 12971
rect 52089 12931 52147 12937
rect 52270 12928 52276 12980
rect 52328 12928 52334 12980
rect 53558 12928 53564 12980
rect 53616 12968 53622 12980
rect 54113 12971 54171 12977
rect 54113 12968 54125 12971
rect 53616 12940 54125 12968
rect 53616 12928 53622 12940
rect 54113 12937 54125 12940
rect 54159 12937 54171 12971
rect 54113 12931 54171 12937
rect 54202 12928 54208 12980
rect 54260 12968 54266 12980
rect 54260 12940 57974 12968
rect 54260 12928 54266 12940
rect 47780 12900 47808 12928
rect 46860 12872 47808 12900
rect 46860 12773 46888 12872
rect 47026 12792 47032 12844
rect 47084 12792 47090 12844
rect 47118 12792 47124 12844
rect 47176 12792 47182 12844
rect 47670 12792 47676 12844
rect 47728 12832 47734 12844
rect 47765 12835 47823 12841
rect 47765 12832 47777 12835
rect 47728 12804 47777 12832
rect 47728 12792 47734 12804
rect 47765 12801 47777 12804
rect 47811 12801 47823 12835
rect 47765 12795 47823 12801
rect 47946 12792 47952 12844
rect 48004 12822 48010 12844
rect 48685 12835 48743 12841
rect 48004 12794 48039 12822
rect 48685 12801 48697 12835
rect 48731 12832 48743 12835
rect 49988 12832 50016 12928
rect 50614 12860 50620 12912
rect 50672 12860 50678 12912
rect 48731 12804 50016 12832
rect 48731 12801 48743 12804
rect 48685 12795 48743 12801
rect 48004 12792 48010 12794
rect 50062 12792 50068 12844
rect 50120 12792 50126 12844
rect 50341 12835 50399 12841
rect 50341 12801 50353 12835
rect 50387 12832 50399 12835
rect 50706 12832 50712 12844
rect 50387 12804 50712 12832
rect 50387 12801 50399 12804
rect 50341 12795 50399 12801
rect 50706 12792 50712 12804
rect 50764 12792 50770 12844
rect 46845 12767 46903 12773
rect 46845 12733 46857 12767
rect 46891 12733 46903 12767
rect 46845 12727 46903 12733
rect 47044 12696 47072 12792
rect 47949 12791 47961 12792
rect 47995 12791 48007 12792
rect 47949 12785 48007 12791
rect 48409 12767 48467 12773
rect 48409 12733 48421 12767
rect 48455 12764 48467 12767
rect 49145 12767 49203 12773
rect 49145 12764 49157 12767
rect 48455 12736 49157 12764
rect 48455 12733 48467 12736
rect 48409 12727 48467 12733
rect 49145 12733 49157 12736
rect 49191 12733 49203 12767
rect 49145 12727 49203 12733
rect 49694 12724 49700 12776
rect 49752 12724 49758 12776
rect 50080 12696 50108 12792
rect 50617 12767 50675 12773
rect 50617 12733 50629 12767
rect 50663 12764 50675 12767
rect 50908 12764 50936 12928
rect 51626 12900 51632 12912
rect 51092 12872 51632 12900
rect 51092 12841 51120 12872
rect 51626 12860 51632 12872
rect 51684 12860 51690 12912
rect 51077 12835 51135 12841
rect 51077 12801 51089 12835
rect 51123 12832 51135 12835
rect 51166 12832 51172 12844
rect 51123 12804 51172 12832
rect 51123 12801 51135 12804
rect 51077 12795 51135 12801
rect 51166 12792 51172 12804
rect 51224 12792 51230 12844
rect 51261 12835 51319 12841
rect 51261 12801 51273 12835
rect 51307 12832 51319 12835
rect 51828 12832 51856 12928
rect 52288 12841 52316 12928
rect 52549 12903 52607 12909
rect 52549 12869 52561 12903
rect 52595 12900 52607 12903
rect 55306 12900 55312 12912
rect 52595 12872 52684 12900
rect 52595 12869 52607 12872
rect 52549 12863 52607 12869
rect 51307 12804 51856 12832
rect 52273 12835 52331 12841
rect 51307 12801 51319 12804
rect 51261 12795 51319 12801
rect 52273 12801 52285 12835
rect 52319 12801 52331 12835
rect 52656 12832 52684 12872
rect 53852 12872 55312 12900
rect 53852 12844 53880 12872
rect 55306 12860 55312 12872
rect 55364 12900 55370 12912
rect 56502 12909 56508 12912
rect 56485 12903 56508 12909
rect 55364 12872 56272 12900
rect 55364 12860 55370 12872
rect 52989 12835 53047 12841
rect 52989 12832 53001 12835
rect 52656 12804 53001 12832
rect 52273 12795 52331 12801
rect 52989 12801 53001 12804
rect 53035 12801 53047 12835
rect 52989 12795 53047 12801
rect 53834 12792 53840 12844
rect 53892 12792 53898 12844
rect 53926 12792 53932 12844
rect 53984 12832 53990 12844
rect 54205 12835 54263 12841
rect 54205 12832 54217 12835
rect 53984 12804 54217 12832
rect 53984 12792 53990 12804
rect 54205 12801 54217 12804
rect 54251 12832 54263 12835
rect 54665 12835 54723 12841
rect 54665 12832 54677 12835
rect 54251 12804 54677 12832
rect 54251 12801 54263 12804
rect 54205 12795 54263 12801
rect 54665 12801 54677 12804
rect 54711 12801 54723 12835
rect 54665 12795 54723 12801
rect 54754 12792 54760 12844
rect 54812 12792 54818 12844
rect 56244 12841 56272 12872
rect 56485 12869 56497 12903
rect 56485 12863 56508 12869
rect 56502 12860 56508 12863
rect 56560 12860 56566 12912
rect 56229 12835 56287 12841
rect 56229 12801 56241 12835
rect 56275 12801 56287 12835
rect 57946 12832 57974 12940
rect 58526 12928 58532 12980
rect 58584 12928 58590 12980
rect 58066 12832 58072 12844
rect 57946 12804 58072 12832
rect 56229 12795 56287 12801
rect 58066 12792 58072 12804
rect 58124 12792 58130 12844
rect 50663 12736 50936 12764
rect 50663 12733 50675 12736
rect 50617 12727 50675 12733
rect 51534 12724 51540 12776
rect 51592 12724 51598 12776
rect 52549 12767 52607 12773
rect 52012 12756 52316 12764
rect 52012 12736 52500 12756
rect 51074 12696 51080 12708
rect 47044 12668 48636 12696
rect 50080 12668 51080 12696
rect 48498 12588 48504 12640
rect 48556 12588 48562 12640
rect 48608 12637 48636 12668
rect 51074 12656 51080 12668
rect 51132 12656 51138 12708
rect 48593 12631 48651 12637
rect 48593 12597 48605 12631
rect 48639 12628 48651 12631
rect 50433 12631 50491 12637
rect 50433 12628 50445 12631
rect 48639 12600 50445 12628
rect 48639 12597 48651 12600
rect 48593 12591 48651 12597
rect 50433 12597 50445 12600
rect 50479 12628 50491 12631
rect 52012 12628 52040 12736
rect 52288 12728 52500 12736
rect 50479 12600 52040 12628
rect 52365 12631 52423 12637
rect 50479 12597 50491 12600
rect 50433 12591 50491 12597
rect 52365 12597 52377 12631
rect 52411 12628 52423 12631
rect 52472 12628 52500 12728
rect 52549 12733 52561 12767
rect 52595 12764 52607 12767
rect 52638 12764 52644 12776
rect 52595 12736 52644 12764
rect 52595 12733 52607 12736
rect 52549 12727 52607 12733
rect 52638 12724 52644 12736
rect 52696 12724 52702 12776
rect 52730 12724 52736 12776
rect 52788 12724 52794 12776
rect 54297 12767 54355 12773
rect 54297 12733 54309 12767
rect 54343 12733 54355 12767
rect 54297 12727 54355 12733
rect 54481 12767 54539 12773
rect 54481 12733 54493 12767
rect 54527 12764 54539 12767
rect 55033 12767 55091 12773
rect 55033 12764 55045 12767
rect 54527 12736 55045 12764
rect 54527 12733 54539 12736
rect 54481 12727 54539 12733
rect 55033 12733 55045 12736
rect 55079 12733 55091 12767
rect 55033 12727 55091 12733
rect 55677 12767 55735 12773
rect 55677 12733 55689 12767
rect 55723 12764 55735 12767
rect 56134 12764 56140 12776
rect 55723 12736 56140 12764
rect 55723 12733 55735 12736
rect 55677 12727 55735 12733
rect 54312 12696 54340 12727
rect 56134 12724 56140 12736
rect 56192 12724 56198 12776
rect 57885 12767 57943 12773
rect 57885 12733 57897 12767
rect 57931 12733 57943 12767
rect 57885 12727 57943 12733
rect 54846 12696 54852 12708
rect 54312 12668 54852 12696
rect 54312 12628 54340 12668
rect 54846 12656 54852 12668
rect 54904 12656 54910 12708
rect 57609 12699 57667 12705
rect 57609 12665 57621 12699
rect 57655 12696 57667 12699
rect 57900 12696 57928 12727
rect 57655 12668 57928 12696
rect 57655 12665 57667 12668
rect 57609 12659 57667 12665
rect 58342 12656 58348 12708
rect 58400 12656 58406 12708
rect 52411 12600 54340 12628
rect 52411 12597 52423 12600
rect 52365 12591 52423 12597
rect 54386 12588 54392 12640
rect 54444 12588 54450 12640
rect 54478 12588 54484 12640
rect 54536 12628 54542 12640
rect 58360 12628 58388 12656
rect 54536 12600 58388 12628
rect 54536 12588 54542 12600
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 49694 12384 49700 12436
rect 49752 12424 49758 12436
rect 49789 12427 49847 12433
rect 49789 12424 49801 12427
rect 49752 12396 49801 12424
rect 49752 12384 49758 12396
rect 49789 12393 49801 12396
rect 49835 12393 49847 12427
rect 49789 12387 49847 12393
rect 51534 12384 51540 12436
rect 51592 12424 51598 12436
rect 51629 12427 51687 12433
rect 51629 12424 51641 12427
rect 51592 12396 51641 12424
rect 51592 12384 51598 12396
rect 51629 12393 51641 12396
rect 51675 12393 51687 12427
rect 51629 12387 51687 12393
rect 52086 12384 52092 12436
rect 52144 12384 52150 12436
rect 55950 12384 55956 12436
rect 56008 12384 56014 12436
rect 56134 12384 56140 12436
rect 56192 12384 56198 12436
rect 56594 12384 56600 12436
rect 56652 12424 56658 12436
rect 56781 12427 56839 12433
rect 56781 12424 56793 12427
rect 56652 12396 56793 12424
rect 56652 12384 56658 12396
rect 56781 12393 56793 12396
rect 56827 12393 56839 12427
rect 56781 12387 56839 12393
rect 55125 12359 55183 12365
rect 55125 12325 55137 12359
rect 55171 12325 55183 12359
rect 55125 12319 55183 12325
rect 46382 12248 46388 12300
rect 46440 12288 46446 12300
rect 48225 12291 48283 12297
rect 48225 12288 48237 12291
rect 46440 12260 48237 12288
rect 46440 12248 46446 12260
rect 48225 12257 48237 12260
rect 48271 12257 48283 12291
rect 52730 12288 52736 12300
rect 48225 12251 48283 12257
rect 51920 12260 52736 12288
rect 48498 12229 48504 12232
rect 48492 12220 48504 12229
rect 48459 12192 48504 12220
rect 48492 12183 48504 12192
rect 48498 12180 48504 12183
rect 48556 12180 48562 12232
rect 49697 12223 49755 12229
rect 49697 12189 49709 12223
rect 49743 12220 49755 12223
rect 49743 12192 49832 12220
rect 49743 12189 49755 12192
rect 49697 12183 49755 12189
rect 49602 12044 49608 12096
rect 49660 12044 49666 12096
rect 49804 12084 49832 12192
rect 49878 12180 49884 12232
rect 49936 12180 49942 12232
rect 50249 12223 50307 12229
rect 50249 12189 50261 12223
rect 50295 12220 50307 12223
rect 50982 12220 50988 12232
rect 50295 12192 50988 12220
rect 50295 12189 50307 12192
rect 50249 12183 50307 12189
rect 50982 12180 50988 12192
rect 51040 12220 51046 12232
rect 51920 12220 51948 12260
rect 52730 12248 52736 12260
rect 52788 12288 52794 12300
rect 55140 12288 55168 12319
rect 55309 12291 55367 12297
rect 55309 12288 55321 12291
rect 52788 12260 53604 12288
rect 55140 12260 55321 12288
rect 52788 12248 52794 12260
rect 51040 12192 51948 12220
rect 51997 12223 52055 12229
rect 51040 12180 51046 12192
rect 51997 12189 52009 12223
rect 52043 12220 52055 12223
rect 52086 12220 52092 12232
rect 52043 12192 52092 12220
rect 52043 12189 52055 12192
rect 51997 12183 52055 12189
rect 52086 12180 52092 12192
rect 52144 12180 52150 12232
rect 52181 12223 52239 12229
rect 52181 12189 52193 12223
rect 52227 12220 52239 12223
rect 52914 12220 52920 12232
rect 52227 12192 52920 12220
rect 52227 12189 52239 12192
rect 52181 12183 52239 12189
rect 52914 12180 52920 12192
rect 52972 12180 52978 12232
rect 53576 12220 53604 12260
rect 55309 12257 55321 12260
rect 55355 12257 55367 12291
rect 55309 12251 55367 12257
rect 53745 12223 53803 12229
rect 53745 12220 53757 12223
rect 53576 12192 53757 12220
rect 53745 12189 53757 12192
rect 53791 12220 53803 12223
rect 53834 12220 53840 12232
rect 53791 12192 53840 12220
rect 53791 12189 53803 12192
rect 53745 12183 53803 12189
rect 53834 12180 53840 12192
rect 53892 12180 53898 12232
rect 54012 12223 54070 12229
rect 54012 12189 54024 12223
rect 54058 12220 54070 12223
rect 54386 12220 54392 12232
rect 54058 12192 54392 12220
rect 54058 12189 54070 12192
rect 54012 12183 54070 12189
rect 54386 12180 54392 12192
rect 54444 12180 54450 12232
rect 55968 12220 55996 12384
rect 56042 12316 56048 12368
rect 56100 12356 56106 12368
rect 58253 12359 58311 12365
rect 58253 12356 58265 12359
rect 56100 12328 58265 12356
rect 56100 12316 56106 12328
rect 58253 12325 58265 12328
rect 58299 12325 58311 12359
rect 58253 12319 58311 12325
rect 57425 12291 57483 12297
rect 57425 12257 57437 12291
rect 57471 12288 57483 12291
rect 57609 12291 57667 12297
rect 57609 12288 57621 12291
rect 57471 12260 57621 12288
rect 57471 12257 57483 12260
rect 57425 12251 57483 12257
rect 57609 12257 57621 12260
rect 57655 12257 57667 12291
rect 57609 12251 57667 12257
rect 57716 12260 58296 12288
rect 56045 12223 56103 12229
rect 56045 12220 56057 12223
rect 55968 12192 56057 12220
rect 56045 12189 56057 12192
rect 56091 12189 56103 12223
rect 56045 12183 56103 12189
rect 56229 12223 56287 12229
rect 56229 12189 56241 12223
rect 56275 12220 56287 12223
rect 56318 12220 56324 12232
rect 56275 12192 56324 12220
rect 56275 12189 56287 12192
rect 56229 12183 56287 12189
rect 50522 12161 50528 12164
rect 50516 12152 50528 12161
rect 50483 12124 50528 12152
rect 50516 12115 50528 12124
rect 50522 12112 50528 12115
rect 50580 12112 50586 12164
rect 50632 12124 51074 12152
rect 50632 12084 50660 12124
rect 49804 12056 50660 12084
rect 51046 12084 51074 12124
rect 51626 12084 51632 12096
rect 51046 12056 51632 12084
rect 51626 12044 51632 12056
rect 51684 12084 51690 12096
rect 52086 12084 52092 12096
rect 51684 12056 52092 12084
rect 51684 12044 51690 12056
rect 52086 12044 52092 12056
rect 52144 12084 52150 12096
rect 56244 12084 56272 12183
rect 56318 12180 56324 12192
rect 56376 12220 56382 12232
rect 57716 12229 57744 12260
rect 58268 12232 58296 12260
rect 57517 12223 57575 12229
rect 57517 12220 57529 12223
rect 56376 12192 57529 12220
rect 56376 12180 56382 12192
rect 57517 12189 57529 12192
rect 57563 12189 57575 12223
rect 57517 12183 57575 12189
rect 57701 12223 57759 12229
rect 57701 12189 57713 12223
rect 57747 12189 57759 12223
rect 57701 12183 57759 12189
rect 57885 12223 57943 12229
rect 57885 12189 57897 12223
rect 57931 12189 57943 12223
rect 58161 12223 58219 12229
rect 58161 12220 58173 12223
rect 57885 12183 57943 12189
rect 58084 12192 58173 12220
rect 57900 12152 57928 12183
rect 57974 12152 57980 12164
rect 57900 12124 57980 12152
rect 57974 12112 57980 12124
rect 58032 12112 58038 12164
rect 58084 12093 58112 12192
rect 58161 12189 58173 12192
rect 58207 12189 58219 12223
rect 58161 12183 58219 12189
rect 58250 12180 58256 12232
rect 58308 12180 58314 12232
rect 52144 12056 56272 12084
rect 58069 12087 58127 12093
rect 52144 12044 52150 12056
rect 58069 12053 58081 12087
rect 58115 12053 58127 12087
rect 58069 12047 58127 12053
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 49602 11840 49608 11892
rect 49660 11840 49666 11892
rect 49878 11840 49884 11892
rect 49936 11880 49942 11892
rect 50341 11883 50399 11889
rect 50341 11880 50353 11883
rect 49936 11852 50353 11880
rect 49936 11840 49942 11852
rect 50341 11849 50353 11852
rect 50387 11849 50399 11883
rect 50341 11843 50399 11849
rect 58069 11883 58127 11889
rect 58069 11849 58081 11883
rect 58115 11849 58127 11883
rect 58069 11843 58127 11849
rect 2682 11704 2688 11756
rect 2740 11704 2746 11756
rect 49620 11744 49648 11840
rect 49697 11747 49755 11753
rect 49697 11744 49709 11747
rect 49620 11716 49709 11744
rect 49697 11713 49709 11716
rect 49743 11713 49755 11747
rect 49697 11707 49755 11713
rect 57885 11747 57943 11753
rect 57885 11713 57897 11747
rect 57931 11713 57943 11747
rect 58084 11744 58112 11843
rect 58161 11747 58219 11753
rect 58161 11744 58173 11747
rect 58084 11716 58173 11744
rect 57885 11707 57943 11713
rect 58161 11713 58173 11716
rect 58207 11713 58219 11747
rect 58161 11707 58219 11713
rect 934 11636 940 11688
rect 992 11676 998 11688
rect 1581 11679 1639 11685
rect 1581 11676 1593 11679
rect 992 11648 1593 11676
rect 992 11636 998 11648
rect 1581 11645 1593 11648
rect 1627 11645 1639 11679
rect 1581 11639 1639 11645
rect 52362 11636 52368 11688
rect 52420 11636 52426 11688
rect 57900 11676 57928 11707
rect 57900 11648 58664 11676
rect 52380 11608 52408 11636
rect 58253 11611 58311 11617
rect 58253 11608 58265 11611
rect 52380 11580 58265 11608
rect 58253 11577 58265 11580
rect 58299 11577 58311 11611
rect 58253 11571 58311 11577
rect 58636 11552 58664 11648
rect 58618 11500 58624 11552
rect 58676 11500 58682 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 48774 10752 48780 10804
rect 48832 10792 48838 10804
rect 49237 10795 49295 10801
rect 49237 10792 49249 10795
rect 48832 10764 49249 10792
rect 48832 10752 48838 10764
rect 49237 10761 49249 10764
rect 49283 10761 49295 10795
rect 49237 10755 49295 10761
rect 49329 10659 49387 10665
rect 49329 10625 49341 10659
rect 49375 10656 49387 10659
rect 58529 10659 58587 10665
rect 49375 10628 51074 10656
rect 49375 10625 49387 10628
rect 49329 10619 49387 10625
rect 51046 10520 51074 10628
rect 58529 10625 58541 10659
rect 58575 10656 58587 10659
rect 58575 10628 58940 10656
rect 58575 10625 58587 10628
rect 58529 10619 58587 10625
rect 58912 10532 58940 10628
rect 58345 10523 58403 10529
rect 58345 10520 58357 10523
rect 51046 10492 58357 10520
rect 58345 10489 58357 10492
rect 58391 10489 58403 10523
rect 58345 10483 58403 10489
rect 58894 10480 58900 10532
rect 58952 10480 58958 10532
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 57974 10208 57980 10260
rect 58032 10248 58038 10260
rect 58345 10251 58403 10257
rect 58345 10248 58357 10251
rect 58032 10220 58357 10248
rect 58032 10208 58038 10220
rect 58345 10217 58357 10220
rect 58391 10217 58403 10251
rect 58345 10211 58403 10217
rect 2685 10047 2743 10053
rect 2685 10013 2697 10047
rect 2731 10044 2743 10047
rect 10226 10044 10232 10056
rect 2731 10016 10232 10044
rect 2731 10013 2743 10016
rect 2685 10007 2743 10013
rect 10226 10004 10232 10016
rect 10284 10004 10290 10056
rect 58529 10047 58587 10053
rect 58529 10013 58541 10047
rect 58575 10044 58587 10047
rect 58575 10016 58940 10044
rect 58575 10013 58587 10016
rect 58529 10007 58587 10013
rect 1578 9936 1584 9988
rect 1636 9936 1642 9988
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 58912 9716 58940 10016
rect 58894 9664 58900 9716
rect 58952 9664 58958 9716
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 58342 9120 58348 9172
rect 58400 9120 58406 9172
rect 58529 8959 58587 8965
rect 58529 8925 58541 8959
rect 58575 8925 58587 8959
rect 58529 8919 58587 8925
rect 58544 8888 58572 8919
rect 58894 8888 58900 8900
rect 58544 8860 58900 8888
rect 58894 8848 58900 8860
rect 58952 8848 58958 8900
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 58066 8576 58072 8628
rect 58124 8616 58130 8628
rect 58345 8619 58403 8625
rect 58345 8616 58357 8619
rect 58124 8588 58357 8616
rect 58124 8576 58130 8588
rect 58345 8585 58357 8588
rect 58391 8585 58403 8619
rect 58345 8579 58403 8585
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8480 2743 8483
rect 9306 8480 9312 8492
rect 2731 8452 9312 8480
rect 2731 8449 2743 8452
rect 2685 8443 2743 8449
rect 9306 8440 9312 8452
rect 9364 8440 9370 8492
rect 58529 8483 58587 8489
rect 58529 8449 58541 8483
rect 58575 8480 58587 8483
rect 58575 8452 58940 8480
rect 58575 8449 58587 8452
rect 58529 8443 58587 8449
rect 1578 8372 1584 8424
rect 1636 8372 1642 8424
rect 58912 8356 58940 8452
rect 58894 8304 58900 8356
rect 58952 8304 58958 8356
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 58529 7395 58587 7401
rect 58529 7361 58541 7395
rect 58575 7392 58587 7395
rect 58575 7364 58940 7392
rect 58575 7361 58587 7364
rect 58529 7355 58587 7361
rect 58912 7268 58940 7364
rect 58894 7216 58900 7268
rect 58952 7216 58958 7268
rect 49234 7148 49240 7200
rect 49292 7188 49298 7200
rect 58345 7191 58403 7197
rect 58345 7188 58357 7191
rect 49292 7160 58357 7188
rect 49292 7148 49298 7160
rect 58345 7157 58357 7160
rect 58391 7157 58403 7191
rect 58345 7151 58403 7157
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 2682 6740 2688 6792
rect 2740 6740 2746 6792
rect 934 6672 940 6724
rect 992 6712 998 6724
rect 1581 6715 1639 6721
rect 1581 6712 1593 6715
rect 992 6684 1593 6712
rect 992 6672 998 6684
rect 1581 6681 1593 6684
rect 1627 6681 1639 6715
rect 1581 6675 1639 6681
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 2685 5219 2743 5225
rect 2685 5185 2697 5219
rect 2731 5216 2743 5219
rect 4614 5216 4620 5228
rect 2731 5188 4620 5216
rect 2731 5185 2743 5188
rect 2685 5179 2743 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 934 5108 940 5160
rect 992 5148 998 5160
rect 1581 5151 1639 5157
rect 1581 5148 1593 5151
rect 992 5120 1593 5148
rect 992 5108 998 5120
rect 1581 5117 1593 5120
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 2685 3519 2743 3525
rect 2685 3485 2697 3519
rect 2731 3516 2743 3519
rect 9030 3516 9036 3528
rect 2731 3488 9036 3516
rect 2731 3485 2743 3488
rect 2685 3479 2743 3485
rect 9030 3476 9036 3488
rect 9088 3476 9094 3528
rect 934 3408 940 3460
rect 992 3448 998 3460
rect 1581 3451 1639 3457
rect 1581 3448 1593 3451
rect 992 3420 1593 3448
rect 992 3408 998 3420
rect 1581 3417 1593 3420
rect 1627 3417 1639 3451
rect 1581 3411 1639 3417
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 12802 2592 12808 2644
rect 12860 2592 12866 2644
rect 15378 2592 15384 2644
rect 15436 2592 15442 2644
rect 42610 2592 42616 2644
rect 42668 2592 42674 2644
rect 49786 2592 49792 2644
rect 49844 2632 49850 2644
rect 56137 2635 56195 2641
rect 56137 2632 56149 2635
rect 49844 2604 56149 2632
rect 49844 2592 49850 2604
rect 56137 2601 56149 2604
rect 56183 2601 56195 2635
rect 56137 2595 56195 2601
rect 9217 2567 9275 2573
rect 9217 2533 9229 2567
rect 9263 2564 9275 2567
rect 15396 2564 15424 2592
rect 29273 2567 29331 2573
rect 29273 2564 29285 2567
rect 9263 2536 15424 2564
rect 28920 2536 29285 2564
rect 9263 2533 9275 2536
rect 9217 2527 9275 2533
rect 3605 2431 3663 2437
rect 3605 2397 3617 2431
rect 3651 2428 3663 2431
rect 8757 2431 8815 2437
rect 3651 2400 4108 2428
rect 3651 2397 3663 2400
rect 3605 2391 3663 2397
rect 2590 2320 2596 2372
rect 2648 2320 2654 2372
rect 4080 2304 4108 2400
rect 8757 2397 8769 2431
rect 8803 2428 8815 2431
rect 9232 2428 9260 2527
rect 11790 2456 11796 2508
rect 11848 2496 11854 2508
rect 22833 2499 22891 2505
rect 22833 2496 22845 2499
rect 11848 2468 22845 2496
rect 11848 2456 11854 2468
rect 22833 2465 22845 2468
rect 22879 2465 22891 2499
rect 22833 2459 22891 2465
rect 8803 2400 9260 2428
rect 8803 2397 8815 2400
rect 8757 2391 8815 2397
rect 12618 2388 12624 2440
rect 12676 2388 12682 2440
rect 17586 2388 17592 2440
rect 17644 2388 17650 2440
rect 22554 2388 22560 2440
rect 22612 2388 22618 2440
rect 28920 2437 28948 2536
rect 29273 2533 29285 2536
rect 29319 2564 29331 2567
rect 29319 2536 35894 2564
rect 29319 2533 29331 2536
rect 29273 2527 29331 2533
rect 32493 2499 32551 2505
rect 32493 2496 32505 2499
rect 29012 2468 32505 2496
rect 28905 2431 28963 2437
rect 26206 2400 27844 2428
rect 7558 2320 7564 2372
rect 7616 2320 7622 2372
rect 9214 2320 9220 2372
rect 9272 2360 9278 2372
rect 26206 2360 26234 2400
rect 9272 2332 26234 2360
rect 9272 2320 9278 2332
rect 27706 2320 27712 2372
rect 27764 2320 27770 2372
rect 27816 2360 27844 2400
rect 28905 2397 28917 2431
rect 28951 2397 28963 2431
rect 28905 2391 28963 2397
rect 29012 2360 29040 2468
rect 32493 2465 32505 2468
rect 32539 2465 32551 2499
rect 35866 2496 35894 2536
rect 45646 2496 45652 2508
rect 35866 2468 45652 2496
rect 32493 2459 32551 2465
rect 45646 2456 45652 2468
rect 45704 2456 45710 2508
rect 47670 2456 47676 2508
rect 47728 2496 47734 2508
rect 48041 2499 48099 2505
rect 48041 2496 48053 2499
rect 47728 2468 48053 2496
rect 47728 2456 47734 2468
rect 48041 2465 48053 2468
rect 48087 2465 48099 2499
rect 48041 2459 48099 2465
rect 27816 2332 29040 2360
rect 29104 2400 35894 2428
rect 4062 2252 4068 2304
rect 4120 2252 4126 2304
rect 12434 2252 12440 2304
rect 12492 2292 12498 2304
rect 29104 2292 29132 2400
rect 32398 2320 32404 2372
rect 32456 2360 32462 2372
rect 32677 2363 32735 2369
rect 32677 2360 32689 2363
rect 32456 2332 32689 2360
rect 32456 2320 32462 2332
rect 32677 2329 32689 2332
rect 32723 2329 32735 2363
rect 32677 2323 32735 2329
rect 12492 2264 29132 2292
rect 35866 2292 35894 2400
rect 38654 2388 38660 2440
rect 38712 2428 38718 2440
rect 39117 2431 39175 2437
rect 39117 2428 39129 2431
rect 38712 2400 39129 2428
rect 38712 2388 38718 2400
rect 39117 2397 39129 2400
rect 39163 2397 39175 2431
rect 39117 2391 39175 2397
rect 42426 2388 42432 2440
rect 42484 2388 42490 2440
rect 47210 2388 47216 2440
rect 47268 2428 47274 2440
rect 47581 2431 47639 2437
rect 47581 2428 47593 2431
rect 47268 2400 47593 2428
rect 47268 2388 47274 2400
rect 47581 2397 47593 2400
rect 47627 2397 47639 2431
rect 47581 2391 47639 2397
rect 52454 2388 52460 2440
rect 52512 2428 52518 2440
rect 52733 2431 52791 2437
rect 52733 2428 52745 2431
rect 52512 2400 52745 2428
rect 52512 2388 52518 2400
rect 52733 2397 52745 2400
rect 52779 2397 52791 2431
rect 56152 2428 56180 2595
rect 56321 2431 56379 2437
rect 56321 2428 56333 2431
rect 56152 2400 56333 2428
rect 52733 2391 52791 2397
rect 56321 2397 56333 2400
rect 56367 2397 56379 2431
rect 56321 2391 56379 2397
rect 37366 2320 37372 2372
rect 37424 2360 37430 2372
rect 37645 2363 37703 2369
rect 37645 2360 37657 2363
rect 37424 2332 37657 2360
rect 37424 2320 37430 2332
rect 37645 2329 37657 2332
rect 37691 2329 37703 2363
rect 37645 2323 37703 2329
rect 57238 2320 57244 2372
rect 57296 2320 57302 2372
rect 52917 2295 52975 2301
rect 52917 2292 52929 2295
rect 35866 2264 52929 2292
rect 12492 2252 12498 2264
rect 52917 2261 52929 2264
rect 52963 2261 52975 2295
rect 52917 2255 52975 2261
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 4062 1980 4068 2032
rect 4120 2020 4126 2032
rect 42242 2020 42248 2032
rect 4120 1992 42248 2020
rect 4120 1980 4126 1992
rect 42242 1980 42248 1992
rect 42300 1980 42306 2032
<< via1 >>
rect 19574 57638 19626 57690
rect 19638 57638 19690 57690
rect 19702 57638 19754 57690
rect 19766 57638 19818 57690
rect 19830 57638 19882 57690
rect 50294 57638 50346 57690
rect 50358 57638 50410 57690
rect 50422 57638 50474 57690
rect 50486 57638 50538 57690
rect 50550 57638 50602 57690
rect 44916 57468 44968 57520
rect 940 57332 992 57384
rect 46480 57332 46532 57384
rect 3056 57239 3108 57248
rect 3056 57205 3065 57239
rect 3065 57205 3099 57239
rect 3099 57205 3108 57239
rect 3056 57196 3108 57205
rect 4214 57094 4266 57146
rect 4278 57094 4330 57146
rect 4342 57094 4394 57146
rect 4406 57094 4458 57146
rect 4470 57094 4522 57146
rect 34934 57094 34986 57146
rect 34998 57094 35050 57146
rect 35062 57094 35114 57146
rect 35126 57094 35178 57146
rect 35190 57094 35242 57146
rect 19574 56550 19626 56602
rect 19638 56550 19690 56602
rect 19702 56550 19754 56602
rect 19766 56550 19818 56602
rect 19830 56550 19882 56602
rect 50294 56550 50346 56602
rect 50358 56550 50410 56602
rect 50422 56550 50474 56602
rect 50486 56550 50538 56602
rect 50550 56550 50602 56602
rect 4214 56006 4266 56058
rect 4278 56006 4330 56058
rect 4342 56006 4394 56058
rect 4406 56006 4458 56058
rect 4470 56006 4522 56058
rect 34934 56006 34986 56058
rect 34998 56006 35050 56058
rect 35062 56006 35114 56058
rect 35126 56006 35178 56058
rect 35190 56006 35242 56058
rect 940 55632 992 55684
rect 15844 55564 15896 55616
rect 19574 55462 19626 55514
rect 19638 55462 19690 55514
rect 19702 55462 19754 55514
rect 19766 55462 19818 55514
rect 19830 55462 19882 55514
rect 50294 55462 50346 55514
rect 50358 55462 50410 55514
rect 50422 55462 50474 55514
rect 50486 55462 50538 55514
rect 50550 55462 50602 55514
rect 4214 54918 4266 54970
rect 4278 54918 4330 54970
rect 4342 54918 4394 54970
rect 4406 54918 4458 54970
rect 4470 54918 4522 54970
rect 34934 54918 34986 54970
rect 34998 54918 35050 54970
rect 35062 54918 35114 54970
rect 35126 54918 35178 54970
rect 35190 54918 35242 54970
rect 19574 54374 19626 54426
rect 19638 54374 19690 54426
rect 19702 54374 19754 54426
rect 19766 54374 19818 54426
rect 19830 54374 19882 54426
rect 50294 54374 50346 54426
rect 50358 54374 50410 54426
rect 50422 54374 50474 54426
rect 50486 54374 50538 54426
rect 50550 54374 50602 54426
rect 1584 54111 1636 54120
rect 1584 54077 1593 54111
rect 1593 54077 1627 54111
rect 1627 54077 1636 54111
rect 1584 54068 1636 54077
rect 2872 53932 2924 53984
rect 4214 53830 4266 53882
rect 4278 53830 4330 53882
rect 4342 53830 4394 53882
rect 4406 53830 4458 53882
rect 4470 53830 4522 53882
rect 34934 53830 34986 53882
rect 34998 53830 35050 53882
rect 35062 53830 35114 53882
rect 35126 53830 35178 53882
rect 35190 53830 35242 53882
rect 19574 53286 19626 53338
rect 19638 53286 19690 53338
rect 19702 53286 19754 53338
rect 19766 53286 19818 53338
rect 19830 53286 19882 53338
rect 50294 53286 50346 53338
rect 50358 53286 50410 53338
rect 50422 53286 50474 53338
rect 50486 53286 50538 53338
rect 50550 53286 50602 53338
rect 58900 53048 58952 53100
rect 58992 52844 59044 52896
rect 4214 52742 4266 52794
rect 4278 52742 4330 52794
rect 4342 52742 4394 52794
rect 4406 52742 4458 52794
rect 4470 52742 4522 52794
rect 34934 52742 34986 52794
rect 34998 52742 35050 52794
rect 35062 52742 35114 52794
rect 35126 52742 35178 52794
rect 35190 52742 35242 52794
rect 58624 52640 58676 52692
rect 1584 52479 1636 52488
rect 1584 52445 1593 52479
rect 1593 52445 1627 52479
rect 1627 52445 1636 52479
rect 1584 52436 1636 52445
rect 5540 52436 5592 52488
rect 58900 52368 58952 52420
rect 19574 52198 19626 52250
rect 19638 52198 19690 52250
rect 19702 52198 19754 52250
rect 19766 52198 19818 52250
rect 19830 52198 19882 52250
rect 50294 52198 50346 52250
rect 50358 52198 50410 52250
rect 50422 52198 50474 52250
rect 50486 52198 50538 52250
rect 50550 52198 50602 52250
rect 4214 51654 4266 51706
rect 4278 51654 4330 51706
rect 4342 51654 4394 51706
rect 4406 51654 4458 51706
rect 4470 51654 4522 51706
rect 34934 51654 34986 51706
rect 34998 51654 35050 51706
rect 35062 51654 35114 51706
rect 35126 51654 35178 51706
rect 35190 51654 35242 51706
rect 58900 51280 58952 51332
rect 58716 51212 58768 51264
rect 19574 51110 19626 51162
rect 19638 51110 19690 51162
rect 19702 51110 19754 51162
rect 19766 51110 19818 51162
rect 19830 51110 19882 51162
rect 50294 51110 50346 51162
rect 50358 51110 50410 51162
rect 50422 51110 50474 51162
rect 50486 51110 50538 51162
rect 50550 51110 50602 51162
rect 2688 50915 2740 50924
rect 2688 50881 2697 50915
rect 2697 50881 2731 50915
rect 2731 50881 2740 50915
rect 2688 50872 2740 50881
rect 940 50804 992 50856
rect 4214 50566 4266 50618
rect 4278 50566 4330 50618
rect 4342 50566 4394 50618
rect 4406 50566 4458 50618
rect 4470 50566 4522 50618
rect 34934 50566 34986 50618
rect 34998 50566 35050 50618
rect 35062 50566 35114 50618
rect 35126 50566 35178 50618
rect 35190 50566 35242 50618
rect 19574 50022 19626 50074
rect 19638 50022 19690 50074
rect 19702 50022 19754 50074
rect 19766 50022 19818 50074
rect 19830 50022 19882 50074
rect 50294 50022 50346 50074
rect 50358 50022 50410 50074
rect 50422 50022 50474 50074
rect 50486 50022 50538 50074
rect 50550 50022 50602 50074
rect 58808 49716 58860 49768
rect 58900 49716 58952 49768
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 2228 49172 2280 49224
rect 940 49104 992 49156
rect 58348 49079 58400 49088
rect 58348 49045 58357 49079
rect 58357 49045 58391 49079
rect 58391 49045 58400 49079
rect 58348 49036 58400 49045
rect 58900 49036 58952 49088
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 50294 48934 50346 48986
rect 50358 48934 50410 48986
rect 50422 48934 50474 48986
rect 50486 48934 50538 48986
rect 50550 48934 50602 48986
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 58900 48016 58952 48068
rect 57796 47948 57848 48000
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 50294 47846 50346 47898
rect 50358 47846 50410 47898
rect 50422 47846 50474 47898
rect 50486 47846 50538 47898
rect 50550 47846 50602 47898
rect 2596 47651 2648 47660
rect 2596 47617 2605 47651
rect 2605 47617 2639 47651
rect 2639 47617 2648 47651
rect 2596 47608 2648 47617
rect 58900 47608 58952 47660
rect 940 47540 992 47592
rect 59084 47404 59136 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 50294 46758 50346 46810
rect 50358 46758 50410 46810
rect 50422 46758 50474 46810
rect 50486 46758 50538 46810
rect 50550 46758 50602 46810
rect 58900 46384 58952 46436
rect 58348 46359 58400 46368
rect 58348 46325 58357 46359
rect 58357 46325 58391 46359
rect 58391 46325 58400 46359
rect 58348 46316 58400 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 6552 45908 6604 45960
rect 57888 45908 57940 45960
rect 1584 45883 1636 45892
rect 1584 45849 1593 45883
rect 1593 45849 1627 45883
rect 1627 45849 1636 45883
rect 1584 45840 1636 45849
rect 58348 45815 58400 45824
rect 58348 45781 58357 45815
rect 58357 45781 58391 45815
rect 58391 45781 58400 45815
rect 58348 45772 58400 45781
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 50294 45670 50346 45722
rect 50358 45670 50410 45722
rect 50422 45670 50474 45722
rect 50486 45670 50538 45722
rect 50550 45670 50602 45722
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 58992 44752 59044 44804
rect 57520 44684 57572 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 50294 44582 50346 44634
rect 50358 44582 50410 44634
rect 50422 44582 50474 44634
rect 50486 44582 50538 44634
rect 50550 44582 50602 44634
rect 3792 44344 3844 44396
rect 1584 44319 1636 44328
rect 1584 44285 1593 44319
rect 1593 44285 1627 44319
rect 1627 44285 1636 44319
rect 1584 44276 1636 44285
rect 57980 44140 58032 44192
rect 58992 44140 59044 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 58072 43979 58124 43988
rect 58072 43945 58081 43979
rect 58081 43945 58115 43979
rect 58115 43945 58124 43979
rect 58072 43936 58124 43945
rect 58348 43800 58400 43852
rect 57520 43664 57572 43716
rect 57980 43596 58032 43648
rect 58256 43596 58308 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 50294 43494 50346 43546
rect 50358 43494 50410 43546
rect 50422 43494 50474 43546
rect 50486 43494 50538 43546
rect 50550 43494 50602 43546
rect 58072 43392 58124 43444
rect 58164 43392 58216 43444
rect 57796 43324 57848 43376
rect 59084 43256 59136 43308
rect 57428 43231 57480 43240
rect 57428 43197 57437 43231
rect 57437 43197 57471 43231
rect 57471 43197 57480 43231
rect 57428 43188 57480 43197
rect 58440 43188 58492 43240
rect 56692 43095 56744 43104
rect 56692 43061 56701 43095
rect 56701 43061 56735 43095
rect 56735 43061 56744 43095
rect 56692 43052 56744 43061
rect 56784 43095 56836 43104
rect 56784 43061 56793 43095
rect 56793 43061 56827 43095
rect 56827 43061 56836 43095
rect 56784 43052 56836 43061
rect 58808 43120 58860 43172
rect 59176 43120 59228 43172
rect 58532 43052 58584 43104
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 58072 42891 58124 42900
rect 58072 42857 58081 42891
rect 58081 42857 58115 42891
rect 58115 42857 58124 42891
rect 58072 42848 58124 42857
rect 58808 42848 58860 42900
rect 56692 42712 56744 42764
rect 57060 42712 57112 42764
rect 57428 42712 57480 42764
rect 58164 42712 58216 42764
rect 7564 42644 7616 42696
rect 57520 42644 57572 42696
rect 58348 42644 58400 42696
rect 58992 42644 59044 42696
rect 940 42576 992 42628
rect 55680 42576 55732 42628
rect 57796 42576 57848 42628
rect 56876 42508 56928 42560
rect 58072 42508 58124 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 50294 42406 50346 42458
rect 50358 42406 50410 42458
rect 50422 42406 50474 42458
rect 50486 42406 50538 42458
rect 50550 42406 50602 42458
rect 57980 42304 58032 42356
rect 59084 42304 59136 42356
rect 56968 42007 57020 42016
rect 56968 41973 56977 42007
rect 56977 41973 57011 42007
rect 57011 41973 57020 42007
rect 56968 41964 57020 41973
rect 57060 41964 57112 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 58808 41488 58860 41540
rect 58164 41420 58216 41472
rect 58348 41463 58400 41472
rect 58348 41429 58357 41463
rect 58357 41429 58391 41463
rect 58391 41429 58400 41463
rect 58348 41420 58400 41429
rect 58992 41420 59044 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 50294 41318 50346 41370
rect 50358 41318 50410 41370
rect 50422 41318 50474 41370
rect 50486 41318 50538 41370
rect 50550 41318 50602 41370
rect 1400 41123 1452 41132
rect 1400 41089 1409 41123
rect 1409 41089 1443 41123
rect 1443 41089 1452 41123
rect 1400 41080 1452 41089
rect 57980 41080 58032 41132
rect 1216 41012 1268 41064
rect 58164 41216 58216 41268
rect 58256 41123 58308 41132
rect 58256 41089 58265 41123
rect 58265 41089 58299 41123
rect 58299 41089 58308 41123
rect 58256 41080 58308 41089
rect 58440 41123 58492 41132
rect 58440 41089 58449 41123
rect 58449 41089 58483 41123
rect 58483 41089 58492 41123
rect 58440 41080 58492 41089
rect 58164 41055 58216 41064
rect 58164 41021 58173 41055
rect 58173 41021 58207 41055
rect 58207 41021 58216 41055
rect 58164 41012 58216 41021
rect 58808 40944 58860 40996
rect 58072 40919 58124 40928
rect 58072 40885 58081 40919
rect 58081 40885 58115 40919
rect 58115 40885 58124 40919
rect 58072 40876 58124 40885
rect 58256 40919 58308 40928
rect 58256 40885 58265 40919
rect 58265 40885 58299 40919
rect 58299 40885 58308 40919
rect 58256 40876 58308 40885
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 58072 40672 58124 40724
rect 58256 40672 58308 40724
rect 2688 40511 2740 40520
rect 2688 40477 2697 40511
rect 2697 40477 2731 40511
rect 2731 40477 2740 40511
rect 2688 40468 2740 40477
rect 47308 40400 47360 40452
rect 58532 40468 58584 40520
rect 2964 40332 3016 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 50294 40230 50346 40282
rect 50358 40230 50410 40282
rect 50422 40230 50474 40282
rect 50486 40230 50538 40282
rect 50550 40230 50602 40282
rect 2688 40128 2740 40180
rect 1400 39992 1452 40044
rect 3884 40060 3936 40112
rect 8300 40060 8352 40112
rect 57980 40171 58032 40180
rect 57980 40137 57989 40171
rect 57989 40137 58023 40171
rect 58023 40137 58032 40171
rect 57980 40128 58032 40137
rect 57888 40060 57940 40112
rect 58348 40103 58400 40112
rect 58348 40069 58357 40103
rect 58357 40069 58391 40103
rect 58391 40069 58400 40103
rect 58348 40060 58400 40069
rect 7564 40035 7616 40044
rect 7564 40001 7573 40035
rect 7573 40001 7607 40035
rect 7607 40001 7616 40035
rect 7564 39992 7616 40001
rect 8392 39992 8444 40044
rect 3516 39967 3568 39976
rect 3516 39933 3525 39967
rect 3525 39933 3559 39967
rect 3559 39933 3568 39967
rect 3516 39924 3568 39933
rect 1952 39831 2004 39840
rect 1952 39797 1961 39831
rect 1961 39797 1995 39831
rect 1995 39797 2004 39831
rect 1952 39788 2004 39797
rect 3240 39788 3292 39840
rect 9864 39967 9916 39976
rect 9864 39933 9873 39967
rect 9873 39933 9907 39967
rect 9907 39933 9916 39967
rect 9864 39924 9916 39933
rect 10140 39967 10192 39976
rect 10140 39933 10149 39967
rect 10149 39933 10183 39967
rect 10183 39933 10192 39967
rect 10140 39924 10192 39933
rect 57796 39856 57848 39908
rect 11704 39831 11756 39840
rect 11704 39797 11713 39831
rect 11713 39797 11747 39831
rect 11747 39797 11756 39831
rect 11704 39788 11756 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 1400 39627 1452 39636
rect 1400 39593 1409 39627
rect 1409 39593 1443 39627
rect 1443 39593 1452 39627
rect 1400 39584 1452 39593
rect 3516 39584 3568 39636
rect 9864 39584 9916 39636
rect 58072 39584 58124 39636
rect 3792 39448 3844 39500
rect 6552 39491 6604 39500
rect 6552 39457 6561 39491
rect 6561 39457 6595 39491
rect 6595 39457 6604 39491
rect 6552 39448 6604 39457
rect 57060 39448 57112 39500
rect 2412 39312 2464 39364
rect 2964 39312 3016 39364
rect 3240 39423 3292 39432
rect 3240 39389 3249 39423
rect 3249 39389 3283 39423
rect 3283 39389 3292 39423
rect 3240 39380 3292 39389
rect 4620 39423 4672 39432
rect 4620 39389 4629 39423
rect 4629 39389 4663 39423
rect 4663 39389 4672 39423
rect 4620 39380 4672 39389
rect 3240 39244 3292 39296
rect 3332 39244 3384 39296
rect 4068 39287 4120 39296
rect 4068 39253 4077 39287
rect 4077 39253 4111 39287
rect 4111 39253 4120 39287
rect 4068 39244 4120 39253
rect 4804 39287 4856 39296
rect 4804 39253 4813 39287
rect 4813 39253 4847 39287
rect 4847 39253 4856 39287
rect 4804 39244 4856 39253
rect 7196 39287 7248 39296
rect 7196 39253 7205 39287
rect 7205 39253 7239 39287
rect 7239 39253 7248 39287
rect 7196 39244 7248 39253
rect 7748 39423 7800 39432
rect 7748 39389 7757 39423
rect 7757 39389 7791 39423
rect 7791 39389 7800 39423
rect 7748 39380 7800 39389
rect 8668 39423 8720 39432
rect 8668 39389 8677 39423
rect 8677 39389 8711 39423
rect 8711 39389 8720 39423
rect 8668 39380 8720 39389
rect 9128 39244 9180 39296
rect 57888 39423 57940 39432
rect 57888 39389 57897 39423
rect 57897 39389 57931 39423
rect 57931 39389 57940 39423
rect 57888 39380 57940 39389
rect 58164 39380 58216 39432
rect 58348 39423 58400 39432
rect 58348 39389 58357 39423
rect 58357 39389 58391 39423
rect 58391 39389 58400 39423
rect 58348 39380 58400 39389
rect 57336 39244 57388 39296
rect 57612 39244 57664 39296
rect 58256 39244 58308 39296
rect 58532 39244 58584 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 50294 39142 50346 39194
rect 50358 39142 50410 39194
rect 50422 39142 50474 39194
rect 50486 39142 50538 39194
rect 50550 39142 50602 39194
rect 2596 39040 2648 39092
rect 3792 39083 3844 39092
rect 3792 39049 3801 39083
rect 3801 39049 3835 39083
rect 3835 39049 3844 39083
rect 3792 39040 3844 39049
rect 940 38904 992 38956
rect 3700 38836 3752 38888
rect 2412 38768 2464 38820
rect 6552 39040 6604 39092
rect 8208 39040 8260 39092
rect 8300 39040 8352 39092
rect 8668 39040 8720 39092
rect 58072 39040 58124 39092
rect 8484 38947 8536 38956
rect 8484 38913 8493 38947
rect 8493 38913 8527 38947
rect 8527 38913 8536 38947
rect 8484 38904 8536 38913
rect 57980 38904 58032 38956
rect 5264 38879 5316 38888
rect 5264 38845 5273 38879
rect 5273 38845 5307 38879
rect 5307 38845 5316 38879
rect 5264 38836 5316 38845
rect 5540 38879 5592 38888
rect 5540 38845 5549 38879
rect 5549 38845 5583 38879
rect 5583 38845 5592 38879
rect 5540 38836 5592 38845
rect 7932 38879 7984 38888
rect 7932 38845 7941 38879
rect 7941 38845 7975 38879
rect 7975 38845 7984 38879
rect 7932 38836 7984 38845
rect 3516 38743 3568 38752
rect 3516 38709 3525 38743
rect 3525 38709 3559 38743
rect 3559 38709 3568 38743
rect 3516 38700 3568 38709
rect 8760 38836 8812 38888
rect 10232 38700 10284 38752
rect 57336 38700 57388 38752
rect 58256 38768 58308 38820
rect 58164 38700 58216 38752
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 1952 38539 2004 38548
rect 1952 38505 1961 38539
rect 1961 38505 1995 38539
rect 1995 38505 2004 38539
rect 1952 38496 2004 38505
rect 2688 38496 2740 38548
rect 4068 38496 4120 38548
rect 4620 38496 4672 38548
rect 5264 38496 5316 38548
rect 7932 38496 7984 38548
rect 8392 38496 8444 38548
rect 1860 38335 1912 38344
rect 1860 38301 1869 38335
rect 1869 38301 1903 38335
rect 1903 38301 1912 38335
rect 1860 38292 1912 38301
rect 2688 38292 2740 38344
rect 3424 38292 3476 38344
rect 3792 38335 3844 38344
rect 3792 38301 3801 38335
rect 3801 38301 3835 38335
rect 3835 38301 3844 38335
rect 3792 38292 3844 38301
rect 7748 38428 7800 38480
rect 4252 38335 4304 38344
rect 4252 38301 4261 38335
rect 4261 38301 4295 38335
rect 4295 38301 4304 38335
rect 4252 38292 4304 38301
rect 2504 38224 2556 38276
rect 2872 38199 2924 38208
rect 2872 38165 2881 38199
rect 2881 38165 2915 38199
rect 2915 38165 2924 38199
rect 2872 38156 2924 38165
rect 7472 38360 7524 38412
rect 57244 38428 57296 38480
rect 4804 38292 4856 38344
rect 5632 38335 5684 38344
rect 5632 38301 5641 38335
rect 5641 38301 5675 38335
rect 5675 38301 5684 38335
rect 5632 38292 5684 38301
rect 7748 38335 7800 38344
rect 7748 38301 7757 38335
rect 7757 38301 7791 38335
rect 7791 38301 7800 38335
rect 7748 38292 7800 38301
rect 8668 38335 8720 38344
rect 8668 38301 8677 38335
rect 8677 38301 8711 38335
rect 8711 38301 8720 38335
rect 8668 38292 8720 38301
rect 8760 38292 8812 38344
rect 10508 38360 10560 38412
rect 58808 38428 58860 38480
rect 58256 38403 58308 38412
rect 58256 38369 58265 38403
rect 58265 38369 58299 38403
rect 58299 38369 58308 38403
rect 58256 38360 58308 38369
rect 9496 38292 9548 38344
rect 10232 38224 10284 38276
rect 57980 38267 58032 38276
rect 9036 38199 9088 38208
rect 9036 38165 9045 38199
rect 9045 38165 9079 38199
rect 9079 38165 9088 38199
rect 9036 38156 9088 38165
rect 57336 38156 57388 38208
rect 57980 38233 57989 38267
rect 57989 38233 58023 38267
rect 58023 38233 58032 38267
rect 57980 38224 58032 38233
rect 58348 38224 58400 38276
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 50294 38054 50346 38106
rect 50358 38054 50410 38106
rect 50422 38054 50474 38106
rect 50486 38054 50538 38106
rect 50550 38054 50602 38106
rect 2596 37952 2648 38004
rect 2872 37952 2924 38004
rect 2412 37884 2464 37936
rect 3424 37995 3476 38004
rect 3424 37961 3433 37995
rect 3433 37961 3467 37995
rect 3467 37961 3476 37995
rect 3424 37952 3476 37961
rect 3516 37952 3568 38004
rect 7196 37952 7248 38004
rect 7472 37995 7524 38004
rect 7472 37961 7481 37995
rect 7481 37961 7515 37995
rect 7515 37961 7524 37995
rect 7472 37952 7524 37961
rect 8668 37952 8720 38004
rect 9036 37952 9088 38004
rect 58440 37995 58492 38004
rect 58440 37961 58449 37995
rect 58449 37961 58483 37995
rect 58483 37961 58492 37995
rect 58440 37952 58492 37961
rect 3332 37859 3384 37868
rect 3332 37825 3341 37859
rect 3341 37825 3375 37859
rect 3375 37825 3384 37859
rect 3332 37816 3384 37825
rect 4252 37816 4304 37868
rect 2964 37748 3016 37800
rect 3240 37791 3292 37800
rect 3240 37757 3249 37791
rect 3249 37757 3283 37791
rect 3283 37757 3292 37791
rect 3240 37748 3292 37757
rect 4620 37791 4672 37800
rect 4620 37757 4629 37791
rect 4629 37757 4663 37791
rect 4663 37757 4672 37791
rect 4620 37748 4672 37757
rect 5724 37816 5776 37868
rect 8392 37859 8444 37868
rect 8392 37825 8393 37859
rect 8393 37825 8427 37859
rect 8427 37825 8444 37859
rect 8392 37816 8444 37825
rect 59176 37884 59228 37936
rect 8668 37680 8720 37732
rect 4068 37655 4120 37664
rect 4068 37621 4077 37655
rect 4077 37621 4111 37655
rect 4111 37621 4120 37655
rect 4068 37612 4120 37621
rect 7288 37655 7340 37664
rect 7288 37621 7297 37655
rect 7297 37621 7331 37655
rect 7331 37621 7340 37655
rect 7288 37612 7340 37621
rect 56784 37612 56836 37664
rect 58256 37859 58308 37868
rect 58256 37825 58265 37859
rect 58265 37825 58299 37859
rect 58299 37825 58308 37859
rect 58256 37816 58308 37825
rect 58164 37655 58216 37664
rect 58164 37621 58173 37655
rect 58173 37621 58207 37655
rect 58207 37621 58216 37655
rect 58164 37612 58216 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 5724 37408 5776 37460
rect 7288 37408 7340 37460
rect 8668 37451 8720 37460
rect 8668 37417 8677 37451
rect 8677 37417 8711 37451
rect 8711 37417 8720 37451
rect 8668 37408 8720 37417
rect 58256 37408 58308 37460
rect 3332 37272 3384 37324
rect 1584 37247 1636 37256
rect 1584 37213 1593 37247
rect 1593 37213 1627 37247
rect 1627 37213 1636 37247
rect 1584 37204 1636 37213
rect 2780 37247 2832 37256
rect 2780 37213 2789 37247
rect 2789 37213 2823 37247
rect 2823 37213 2832 37247
rect 2780 37204 2832 37213
rect 3700 37272 3752 37324
rect 7656 37272 7708 37324
rect 3976 37136 4028 37188
rect 6092 37136 6144 37188
rect 4620 37068 4672 37120
rect 5356 37068 5408 37120
rect 5540 37068 5592 37120
rect 5724 37068 5776 37120
rect 8392 37247 8444 37256
rect 8392 37213 8401 37247
rect 8401 37213 8435 37247
rect 8435 37213 8444 37247
rect 58900 37272 58952 37324
rect 8392 37204 8444 37213
rect 7472 37111 7524 37120
rect 7472 37077 7481 37111
rect 7481 37077 7515 37111
rect 7515 37077 7524 37111
rect 7472 37068 7524 37077
rect 8760 37068 8812 37120
rect 8944 37111 8996 37120
rect 8944 37077 8953 37111
rect 8953 37077 8987 37111
rect 8987 37077 8996 37111
rect 8944 37068 8996 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 7472 36864 7524 36916
rect 7656 36907 7708 36916
rect 7656 36873 7665 36907
rect 7665 36873 7699 36907
rect 7699 36873 7708 36907
rect 7656 36864 7708 36873
rect 58256 36864 58308 36916
rect 2412 36796 2464 36848
rect 5356 36796 5408 36848
rect 3608 36703 3660 36712
rect 3608 36669 3617 36703
rect 3617 36669 3651 36703
rect 3651 36669 3660 36703
rect 3608 36660 3660 36669
rect 3700 36660 3752 36712
rect 5724 36771 5776 36780
rect 5724 36737 5733 36771
rect 5733 36737 5767 36771
rect 5767 36737 5776 36771
rect 5724 36728 5776 36737
rect 6092 36728 6144 36780
rect 3332 36592 3384 36644
rect 8668 36796 8720 36848
rect 9496 36796 9548 36848
rect 10508 36771 10560 36780
rect 10508 36737 10517 36771
rect 10517 36737 10551 36771
rect 10551 36737 10560 36771
rect 10508 36728 10560 36737
rect 8392 36703 8444 36712
rect 8392 36669 8401 36703
rect 8401 36669 8435 36703
rect 8435 36669 8444 36703
rect 8392 36660 8444 36669
rect 10232 36703 10284 36712
rect 10232 36669 10241 36703
rect 10241 36669 10275 36703
rect 10275 36669 10284 36703
rect 10232 36660 10284 36669
rect 7012 36592 7064 36644
rect 58900 36592 58952 36644
rect 2688 36524 2740 36576
rect 2872 36524 2924 36576
rect 7288 36524 7340 36576
rect 8208 36524 8260 36576
rect 57704 36567 57756 36576
rect 57704 36533 57713 36567
rect 57713 36533 57747 36567
rect 57747 36533 57756 36567
rect 57704 36524 57756 36533
rect 57980 36567 58032 36576
rect 57980 36533 57989 36567
rect 57989 36533 58023 36567
rect 58023 36533 58032 36567
rect 57980 36524 58032 36533
rect 58164 36524 58216 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 2780 36320 2832 36372
rect 3608 36320 3660 36372
rect 3976 36363 4028 36372
rect 3976 36329 3985 36363
rect 3985 36329 4019 36363
rect 4019 36329 4028 36363
rect 3976 36320 4028 36329
rect 4068 36320 4120 36372
rect 8208 36320 8260 36372
rect 8392 36320 8444 36372
rect 8944 36320 8996 36372
rect 10232 36320 10284 36372
rect 57980 36320 58032 36372
rect 58532 36320 58584 36372
rect 3240 36252 3292 36304
rect 2872 36227 2924 36236
rect 2872 36193 2881 36227
rect 2881 36193 2915 36227
rect 2915 36193 2924 36227
rect 2872 36184 2924 36193
rect 3424 36159 3476 36168
rect 3424 36125 3433 36159
rect 3433 36125 3467 36159
rect 3467 36125 3476 36159
rect 3424 36116 3476 36125
rect 2412 36048 2464 36100
rect 3148 36048 3200 36100
rect 3976 36116 4028 36168
rect 4528 36159 4580 36168
rect 4528 36125 4537 36159
rect 4537 36125 4571 36159
rect 4571 36125 4580 36159
rect 4528 36116 4580 36125
rect 7288 36116 7340 36168
rect 8392 36116 8444 36168
rect 8760 36184 8812 36236
rect 57520 36295 57572 36304
rect 57520 36261 57529 36295
rect 57529 36261 57563 36295
rect 57563 36261 57572 36295
rect 57520 36252 57572 36261
rect 4620 36048 4672 36100
rect 2228 35980 2280 36032
rect 6460 36048 6512 36100
rect 58440 36048 58492 36100
rect 4988 35980 5040 36032
rect 8484 35980 8536 36032
rect 58348 36023 58400 36032
rect 58348 35989 58357 36023
rect 58357 35989 58391 36023
rect 58391 35989 58400 36023
rect 58348 35980 58400 35989
rect 58900 35980 58952 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 3424 35776 3476 35828
rect 4528 35776 4580 35828
rect 6184 35819 6236 35828
rect 6184 35785 6193 35819
rect 6193 35785 6227 35819
rect 6227 35785 6236 35819
rect 6184 35776 6236 35785
rect 6460 35819 6512 35828
rect 6460 35785 6469 35819
rect 6469 35785 6503 35819
rect 6503 35785 6512 35819
rect 6460 35776 6512 35785
rect 940 35640 992 35692
rect 4988 35708 5040 35760
rect 6092 35708 6144 35760
rect 58348 35708 58400 35760
rect 2872 35683 2924 35692
rect 2872 35649 2881 35683
rect 2881 35649 2915 35683
rect 2915 35649 2924 35683
rect 2872 35640 2924 35649
rect 4068 35683 4120 35692
rect 4068 35649 4077 35683
rect 4077 35649 4111 35683
rect 4111 35649 4120 35683
rect 4068 35640 4120 35649
rect 3148 35572 3200 35624
rect 10508 35640 10560 35692
rect 17132 35640 17184 35692
rect 58072 35683 58124 35692
rect 58072 35649 58081 35683
rect 58081 35649 58115 35683
rect 58115 35649 58124 35683
rect 58072 35640 58124 35649
rect 2688 35436 2740 35488
rect 3424 35436 3476 35488
rect 3976 35436 4028 35488
rect 5724 35572 5776 35624
rect 8208 35615 8260 35624
rect 8208 35581 8217 35615
rect 8217 35581 8251 35615
rect 8251 35581 8260 35615
rect 8208 35572 8260 35581
rect 8852 35615 8904 35624
rect 8852 35581 8861 35615
rect 8861 35581 8895 35615
rect 8895 35581 8904 35615
rect 8852 35572 8904 35581
rect 58440 35683 58492 35692
rect 58440 35649 58449 35683
rect 58449 35649 58483 35683
rect 58483 35649 58492 35683
rect 58440 35640 58492 35649
rect 4712 35436 4764 35488
rect 56416 35436 56468 35488
rect 57704 35436 57756 35488
rect 57888 35479 57940 35488
rect 57888 35445 57897 35479
rect 57897 35445 57931 35479
rect 57931 35445 57940 35479
rect 57888 35436 57940 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 3332 35232 3384 35284
rect 3884 35275 3936 35284
rect 3884 35241 3893 35275
rect 3893 35241 3927 35275
rect 3927 35241 3936 35275
rect 3884 35232 3936 35241
rect 4712 35275 4764 35284
rect 4712 35241 4721 35275
rect 4721 35241 4755 35275
rect 4755 35241 4764 35275
rect 4712 35232 4764 35241
rect 6184 35232 6236 35284
rect 8852 35232 8904 35284
rect 2596 35028 2648 35080
rect 4988 35028 5040 35080
rect 7288 35207 7340 35216
rect 7288 35173 7297 35207
rect 7297 35173 7331 35207
rect 7331 35173 7340 35207
rect 7288 35164 7340 35173
rect 56048 35164 56100 35216
rect 3700 34960 3752 35012
rect 3056 34935 3108 34944
rect 3056 34901 3065 34935
rect 3065 34901 3099 34935
rect 3099 34901 3108 34935
rect 3056 34892 3108 34901
rect 5172 34892 5224 34944
rect 6644 35028 6696 35080
rect 8484 35071 8536 35080
rect 8484 35037 8493 35071
rect 8493 35037 8527 35071
rect 8527 35037 8536 35071
rect 8484 35028 8536 35037
rect 8300 34960 8352 35012
rect 8760 35028 8812 35080
rect 9128 34960 9180 35012
rect 55312 34892 55364 34944
rect 55864 35071 55916 35080
rect 55864 35037 55873 35071
rect 55873 35037 55907 35071
rect 55907 35037 55916 35071
rect 55864 35028 55916 35037
rect 56140 35071 56192 35080
rect 56140 35037 56149 35071
rect 56149 35037 56183 35071
rect 56183 35037 56192 35071
rect 56140 35028 56192 35037
rect 56968 35028 57020 35080
rect 57060 35071 57112 35080
rect 57060 35037 57069 35071
rect 57069 35037 57103 35071
rect 57103 35037 57112 35071
rect 57060 35028 57112 35037
rect 57244 35071 57296 35080
rect 57244 35037 57253 35071
rect 57253 35037 57287 35071
rect 57287 35037 57296 35071
rect 57244 35028 57296 35037
rect 57704 35096 57756 35148
rect 56416 34892 56468 34944
rect 58900 34960 58952 35012
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 4068 34688 4120 34740
rect 2412 34620 2464 34672
rect 2596 34620 2648 34672
rect 56140 34688 56192 34740
rect 56692 34688 56744 34740
rect 3884 34552 3936 34604
rect 3148 34527 3200 34536
rect 3148 34493 3157 34527
rect 3157 34493 3191 34527
rect 3191 34493 3200 34527
rect 3148 34484 3200 34493
rect 3424 34484 3476 34536
rect 6000 34552 6052 34604
rect 49700 34552 49752 34604
rect 9864 34484 9916 34536
rect 50804 34527 50856 34536
rect 50804 34493 50813 34527
rect 50813 34493 50847 34527
rect 50847 34493 50856 34527
rect 50804 34484 50856 34493
rect 51448 34484 51500 34536
rect 4620 34416 4672 34468
rect 55496 34552 55548 34604
rect 56048 34620 56100 34672
rect 56232 34620 56284 34672
rect 55864 34595 55916 34604
rect 55864 34561 55873 34595
rect 55873 34561 55907 34595
rect 55907 34561 55916 34595
rect 55864 34552 55916 34561
rect 56692 34595 56744 34604
rect 56692 34561 56701 34595
rect 56701 34561 56735 34595
rect 56735 34561 56744 34595
rect 56692 34552 56744 34561
rect 56876 34595 56928 34604
rect 56876 34561 56885 34595
rect 56885 34561 56919 34595
rect 56919 34561 56928 34595
rect 56876 34552 56928 34561
rect 57520 34552 57572 34604
rect 51172 34348 51224 34400
rect 52184 34348 52236 34400
rect 56324 34391 56376 34400
rect 56324 34357 56333 34391
rect 56333 34357 56367 34391
rect 56367 34357 56376 34391
rect 56324 34348 56376 34357
rect 56508 34416 56560 34468
rect 57980 34484 58032 34536
rect 58900 34484 58952 34536
rect 58348 34391 58400 34400
rect 58348 34357 58357 34391
rect 58357 34357 58391 34391
rect 58391 34357 58400 34391
rect 58348 34348 58400 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 3424 34144 3476 34196
rect 6000 34144 6052 34196
rect 6552 34144 6604 34196
rect 50804 34187 50856 34196
rect 50804 34153 50813 34187
rect 50813 34153 50847 34187
rect 50847 34153 50856 34187
rect 50804 34144 50856 34153
rect 52644 34144 52696 34196
rect 56416 34144 56468 34196
rect 57980 34187 58032 34196
rect 57980 34153 57989 34187
rect 57989 34153 58023 34187
rect 58023 34153 58032 34187
rect 57980 34144 58032 34153
rect 58348 34144 58400 34196
rect 940 34008 992 34060
rect 57796 34008 57848 34060
rect 2596 33983 2648 33992
rect 2596 33949 2605 33983
rect 2605 33949 2639 33983
rect 2639 33949 2648 33983
rect 2596 33940 2648 33949
rect 2872 33983 2924 33992
rect 2872 33949 2881 33983
rect 2881 33949 2915 33983
rect 2915 33949 2924 33983
rect 2872 33940 2924 33949
rect 3056 33940 3108 33992
rect 5172 33940 5224 33992
rect 3332 33872 3384 33924
rect 4804 33804 4856 33856
rect 9312 33983 9364 33992
rect 9312 33949 9321 33983
rect 9321 33949 9355 33983
rect 9355 33949 9364 33983
rect 9312 33940 9364 33949
rect 41604 33983 41656 33992
rect 41604 33949 41613 33983
rect 41613 33949 41647 33983
rect 41647 33949 41656 33983
rect 41604 33940 41656 33949
rect 5908 33915 5960 33924
rect 5908 33881 5942 33915
rect 5942 33881 5960 33915
rect 5908 33872 5960 33881
rect 9404 33872 9456 33924
rect 41880 33915 41932 33924
rect 41880 33881 41889 33915
rect 41889 33881 41923 33915
rect 41923 33881 41932 33915
rect 41880 33872 41932 33881
rect 6736 33804 6788 33856
rect 9772 33804 9824 33856
rect 9864 33804 9916 33856
rect 42616 33804 42668 33856
rect 45652 33983 45704 33992
rect 45652 33949 45661 33983
rect 45661 33949 45695 33983
rect 45695 33949 45704 33983
rect 45652 33940 45704 33949
rect 50160 33983 50212 33992
rect 50160 33949 50169 33983
rect 50169 33949 50203 33983
rect 50203 33949 50212 33983
rect 50160 33940 50212 33949
rect 57060 33940 57112 33992
rect 57612 33940 57664 33992
rect 57888 33940 57940 33992
rect 43260 33804 43312 33856
rect 44180 33915 44232 33924
rect 44180 33881 44189 33915
rect 44189 33881 44223 33915
rect 44223 33881 44232 33915
rect 44180 33872 44232 33881
rect 51264 33872 51316 33924
rect 57980 33872 58032 33924
rect 58440 33872 58492 33924
rect 45468 33847 45520 33856
rect 45468 33813 45477 33847
rect 45477 33813 45511 33847
rect 45511 33813 45520 33847
rect 45468 33804 45520 33813
rect 46388 33847 46440 33856
rect 46388 33813 46397 33847
rect 46397 33813 46431 33847
rect 46431 33813 46440 33847
rect 46388 33804 46440 33813
rect 51540 33804 51592 33856
rect 56600 33804 56652 33856
rect 57520 33804 57572 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 4804 33600 4856 33652
rect 4988 33643 5040 33652
rect 4988 33609 4997 33643
rect 4997 33609 5031 33643
rect 5031 33609 5040 33643
rect 4988 33600 5040 33609
rect 5264 33575 5316 33584
rect 5264 33541 5273 33575
rect 5273 33541 5307 33575
rect 5307 33541 5316 33575
rect 5264 33532 5316 33541
rect 5908 33643 5960 33652
rect 5908 33609 5923 33643
rect 5923 33609 5957 33643
rect 5957 33609 5960 33643
rect 5908 33600 5960 33609
rect 6552 33600 6604 33652
rect 6644 33600 6696 33652
rect 6460 33532 6512 33584
rect 4988 33396 5040 33448
rect 6000 33507 6052 33516
rect 6000 33473 6009 33507
rect 6009 33473 6043 33507
rect 6043 33473 6052 33507
rect 6000 33464 6052 33473
rect 6368 33507 6420 33516
rect 6368 33473 6377 33507
rect 6377 33473 6411 33507
rect 6411 33473 6420 33507
rect 6368 33464 6420 33473
rect 9312 33600 9364 33652
rect 6736 33507 6788 33516
rect 6736 33473 6745 33507
rect 6745 33473 6779 33507
rect 6779 33473 6788 33507
rect 6736 33464 6788 33473
rect 7472 33532 7524 33584
rect 7748 33532 7800 33584
rect 9036 33532 9088 33584
rect 7564 33507 7616 33516
rect 7564 33473 7598 33507
rect 7598 33473 7616 33507
rect 7564 33464 7616 33473
rect 7840 33464 7892 33516
rect 9312 33507 9364 33516
rect 9312 33473 9321 33507
rect 9321 33473 9355 33507
rect 9355 33473 9364 33507
rect 9312 33464 9364 33473
rect 9864 33600 9916 33652
rect 41880 33600 41932 33652
rect 43260 33532 43312 33584
rect 45652 33600 45704 33652
rect 6368 33328 6420 33380
rect 9404 33328 9456 33380
rect 5540 33260 5592 33312
rect 6000 33260 6052 33312
rect 7104 33303 7156 33312
rect 7104 33269 7113 33303
rect 7113 33269 7147 33303
rect 7147 33269 7156 33303
rect 7104 33260 7156 33269
rect 42892 33464 42944 33516
rect 44640 33532 44692 33584
rect 49516 33600 49568 33652
rect 49240 33532 49292 33584
rect 50160 33643 50212 33652
rect 50160 33609 50169 33643
rect 50169 33609 50203 33643
rect 50203 33609 50212 33643
rect 50160 33600 50212 33609
rect 50896 33532 50948 33584
rect 10324 33371 10376 33380
rect 10324 33337 10333 33371
rect 10333 33337 10367 33371
rect 10367 33337 10376 33371
rect 10324 33328 10376 33337
rect 43260 33396 43312 33448
rect 46388 33464 46440 33516
rect 46480 33507 46532 33516
rect 46480 33473 46489 33507
rect 46489 33473 46523 33507
rect 46523 33473 46532 33507
rect 46480 33464 46532 33473
rect 46020 33439 46072 33448
rect 46020 33405 46029 33439
rect 46029 33405 46063 33439
rect 46063 33405 46072 33439
rect 46020 33396 46072 33405
rect 47400 33464 47452 33516
rect 47860 33439 47912 33448
rect 47860 33405 47869 33439
rect 47869 33405 47903 33439
rect 47903 33405 47912 33439
rect 47860 33396 47912 33405
rect 49792 33464 49844 33516
rect 51172 33532 51224 33584
rect 50804 33439 50856 33448
rect 50804 33405 50813 33439
rect 50813 33405 50847 33439
rect 50847 33405 50856 33439
rect 50804 33396 50856 33405
rect 51264 33507 51316 33516
rect 51264 33473 51273 33507
rect 51273 33473 51307 33507
rect 51307 33473 51316 33507
rect 51264 33464 51316 33473
rect 51540 33464 51592 33516
rect 52644 33600 52696 33652
rect 55680 33643 55732 33652
rect 55680 33609 55689 33643
rect 55689 33609 55723 33643
rect 55723 33609 55732 33643
rect 55680 33600 55732 33609
rect 56600 33600 56652 33652
rect 57336 33600 57388 33652
rect 58164 33600 58216 33652
rect 52184 33507 52236 33516
rect 52184 33473 52193 33507
rect 52193 33473 52227 33507
rect 52227 33473 52236 33507
rect 52184 33464 52236 33473
rect 55496 33507 55548 33516
rect 55496 33473 55505 33507
rect 55505 33473 55539 33507
rect 55539 33473 55548 33507
rect 55496 33464 55548 33473
rect 56600 33464 56652 33516
rect 43812 33328 43864 33380
rect 50436 33328 50488 33380
rect 57796 33464 57848 33516
rect 57520 33439 57572 33448
rect 57520 33405 57529 33439
rect 57529 33405 57563 33439
rect 57563 33405 57572 33439
rect 57520 33396 57572 33405
rect 57704 33396 57756 33448
rect 9772 33260 9824 33312
rect 10416 33260 10468 33312
rect 44824 33260 44876 33312
rect 50896 33303 50948 33312
rect 50896 33269 50905 33303
rect 50905 33269 50939 33303
rect 50939 33269 50948 33303
rect 50896 33260 50948 33269
rect 50988 33260 51040 33312
rect 58900 33328 58952 33380
rect 52644 33260 52696 33312
rect 55496 33303 55548 33312
rect 55496 33269 55505 33303
rect 55505 33269 55539 33303
rect 55539 33269 55548 33303
rect 55496 33260 55548 33269
rect 56968 33303 57020 33312
rect 56968 33269 56977 33303
rect 56977 33269 57011 33303
rect 57011 33269 57020 33303
rect 56968 33260 57020 33269
rect 57336 33260 57388 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 7564 33056 7616 33108
rect 38384 33056 38436 33108
rect 44088 33056 44140 33108
rect 44272 33056 44324 33108
rect 43260 32988 43312 33040
rect 46020 33056 46072 33108
rect 46112 33056 46164 33108
rect 46480 33056 46532 33108
rect 47860 33056 47912 33108
rect 6460 32920 6512 32972
rect 6828 32920 6880 32972
rect 940 32784 992 32836
rect 1400 32716 1452 32768
rect 7104 32852 7156 32904
rect 41604 32920 41656 32972
rect 7840 32852 7892 32904
rect 40592 32827 40644 32836
rect 40592 32793 40601 32827
rect 40601 32793 40635 32827
rect 40635 32793 40644 32827
rect 40592 32784 40644 32793
rect 3516 32759 3568 32768
rect 3516 32725 3525 32759
rect 3525 32725 3559 32759
rect 3559 32725 3568 32759
rect 3516 32716 3568 32725
rect 4804 32716 4856 32768
rect 6368 32716 6420 32768
rect 7288 32759 7340 32768
rect 7288 32725 7297 32759
rect 7297 32725 7331 32759
rect 7331 32725 7340 32759
rect 7288 32716 7340 32725
rect 7380 32716 7432 32768
rect 41420 32716 41472 32768
rect 42616 32852 42668 32904
rect 42708 32895 42760 32904
rect 42708 32861 42717 32895
rect 42717 32861 42751 32895
rect 42751 32861 42760 32895
rect 42708 32852 42760 32861
rect 42892 32852 42944 32904
rect 43260 32852 43312 32904
rect 43536 32895 43588 32904
rect 43536 32861 43545 32895
rect 43545 32861 43579 32895
rect 43579 32861 43588 32895
rect 43536 32852 43588 32861
rect 43720 32852 43772 32904
rect 55588 33056 55640 33108
rect 56600 33056 56652 33108
rect 57704 33056 57756 33108
rect 50804 32988 50856 33040
rect 56508 32988 56560 33040
rect 44640 32895 44692 32904
rect 44640 32861 44649 32895
rect 44649 32861 44683 32895
rect 44683 32861 44692 32895
rect 44640 32852 44692 32861
rect 44824 32852 44876 32904
rect 42800 32784 42852 32836
rect 43812 32784 43864 32836
rect 44456 32784 44508 32836
rect 47676 32852 47728 32904
rect 48320 32852 48372 32904
rect 49240 32895 49292 32904
rect 49240 32861 49249 32895
rect 49249 32861 49283 32895
rect 49283 32861 49292 32895
rect 49240 32852 49292 32861
rect 50436 32852 50488 32904
rect 50988 32852 51040 32904
rect 48964 32784 49016 32836
rect 56416 32852 56468 32904
rect 56968 32852 57020 32904
rect 57336 32852 57388 32904
rect 57888 32988 57940 33040
rect 58900 32784 58952 32836
rect 42156 32759 42208 32768
rect 42156 32725 42165 32759
rect 42165 32725 42199 32759
rect 42199 32725 42208 32759
rect 42156 32716 42208 32725
rect 43076 32716 43128 32768
rect 43536 32716 43588 32768
rect 44732 32716 44784 32768
rect 49884 32759 49936 32768
rect 49884 32725 49893 32759
rect 49893 32725 49927 32759
rect 49927 32725 49936 32759
rect 49884 32716 49936 32725
rect 51264 32759 51316 32768
rect 51264 32725 51273 32759
rect 51273 32725 51307 32759
rect 51307 32725 51316 32759
rect 51264 32716 51316 32725
rect 51540 32716 51592 32768
rect 52736 32716 52788 32768
rect 56784 32716 56836 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 1400 32555 1452 32564
rect 1400 32521 1409 32555
rect 1409 32521 1443 32555
rect 1443 32521 1452 32555
rect 1400 32512 1452 32521
rect 2872 32512 2924 32564
rect 2412 32444 2464 32496
rect 7288 32512 7340 32564
rect 7472 32512 7524 32564
rect 8576 32555 8628 32564
rect 8576 32521 8585 32555
rect 8585 32521 8619 32555
rect 8619 32521 8628 32555
rect 8576 32512 8628 32521
rect 9312 32512 9364 32564
rect 38384 32555 38436 32564
rect 38384 32521 38393 32555
rect 38393 32521 38427 32555
rect 38427 32521 38436 32555
rect 38384 32512 38436 32521
rect 40592 32512 40644 32564
rect 42156 32512 42208 32564
rect 42708 32512 42760 32564
rect 42800 32512 42852 32564
rect 42892 32555 42944 32564
rect 42892 32521 42901 32555
rect 42901 32521 42935 32555
rect 42935 32521 42944 32555
rect 42892 32512 42944 32521
rect 2872 32351 2924 32360
rect 2872 32317 2881 32351
rect 2881 32317 2915 32351
rect 2915 32317 2924 32351
rect 2872 32308 2924 32317
rect 3148 32351 3200 32360
rect 3148 32317 3157 32351
rect 3157 32317 3191 32351
rect 3191 32317 3200 32351
rect 3148 32308 3200 32317
rect 2504 32172 2556 32224
rect 3792 32351 3844 32360
rect 3792 32317 3801 32351
rect 3801 32317 3835 32351
rect 3835 32317 3844 32351
rect 3792 32308 3844 32317
rect 3884 32308 3936 32360
rect 4804 32376 4856 32428
rect 10324 32444 10376 32496
rect 12440 32444 12492 32496
rect 3424 32240 3476 32292
rect 4068 32172 4120 32224
rect 4620 32215 4672 32224
rect 4620 32181 4629 32215
rect 4629 32181 4663 32215
rect 4663 32181 4672 32215
rect 4620 32172 4672 32181
rect 4988 32172 5040 32224
rect 7840 32172 7892 32224
rect 8852 32376 8904 32428
rect 39028 32419 39080 32428
rect 39028 32385 39037 32419
rect 39037 32385 39071 32419
rect 39071 32385 39080 32419
rect 39028 32376 39080 32385
rect 39212 32419 39264 32428
rect 39212 32385 39221 32419
rect 39221 32385 39255 32419
rect 39255 32385 39264 32419
rect 39212 32376 39264 32385
rect 10232 32351 10284 32360
rect 10232 32317 10241 32351
rect 10241 32317 10275 32351
rect 10275 32317 10284 32351
rect 10232 32308 10284 32317
rect 39488 32419 39540 32428
rect 39488 32385 39497 32419
rect 39497 32385 39531 32419
rect 39531 32385 39540 32419
rect 39488 32376 39540 32385
rect 43720 32444 43772 32496
rect 43812 32444 43864 32496
rect 44272 32512 44324 32564
rect 40592 32351 40644 32360
rect 40592 32317 40601 32351
rect 40601 32317 40635 32351
rect 40635 32317 40644 32351
rect 40592 32308 40644 32317
rect 42064 32308 42116 32360
rect 42892 32419 42944 32428
rect 42892 32385 42901 32419
rect 42901 32385 42935 32419
rect 42935 32385 42944 32419
rect 42892 32376 42944 32385
rect 43076 32419 43128 32428
rect 43076 32385 43085 32419
rect 43085 32385 43119 32419
rect 43119 32385 43128 32419
rect 43076 32376 43128 32385
rect 44548 32487 44600 32496
rect 44548 32453 44557 32487
rect 44557 32453 44591 32487
rect 44591 32453 44600 32487
rect 44548 32444 44600 32453
rect 44916 32512 44968 32564
rect 43628 32308 43680 32360
rect 44180 32308 44232 32360
rect 44916 32376 44968 32428
rect 45652 32512 45704 32564
rect 52736 32512 52788 32564
rect 46664 32444 46716 32496
rect 45468 32376 45520 32428
rect 47400 32419 47452 32428
rect 47400 32385 47409 32419
rect 47409 32385 47443 32419
rect 47443 32385 47452 32419
rect 47400 32376 47452 32385
rect 47676 32376 47728 32428
rect 49884 32444 49936 32496
rect 49240 32376 49292 32428
rect 55128 32512 55180 32564
rect 53748 32444 53800 32496
rect 53196 32376 53248 32428
rect 44456 32283 44508 32292
rect 44456 32249 44465 32283
rect 44465 32249 44499 32283
rect 44499 32249 44508 32283
rect 44456 32240 44508 32249
rect 45560 32308 45612 32360
rect 46664 32308 46716 32360
rect 47032 32351 47084 32360
rect 47032 32317 47041 32351
rect 47041 32317 47075 32351
rect 47075 32317 47084 32351
rect 47032 32308 47084 32317
rect 12348 32172 12400 32224
rect 39304 32172 39356 32224
rect 39396 32215 39448 32224
rect 39396 32181 39405 32215
rect 39405 32181 39439 32215
rect 39439 32181 39448 32215
rect 39396 32172 39448 32181
rect 41236 32215 41288 32224
rect 41236 32181 41245 32215
rect 41245 32181 41279 32215
rect 41279 32181 41288 32215
rect 41236 32172 41288 32181
rect 44640 32172 44692 32224
rect 44732 32215 44784 32224
rect 44732 32181 44741 32215
rect 44741 32181 44775 32215
rect 44775 32181 44784 32215
rect 44732 32172 44784 32181
rect 46204 32240 46256 32292
rect 45560 32172 45612 32224
rect 54392 32351 54444 32360
rect 54392 32317 54401 32351
rect 54401 32317 54435 32351
rect 54435 32317 54444 32351
rect 54392 32308 54444 32317
rect 55588 32351 55640 32360
rect 55588 32317 55597 32351
rect 55597 32317 55631 32351
rect 55631 32317 55640 32351
rect 55588 32308 55640 32317
rect 49056 32172 49108 32224
rect 49516 32172 49568 32224
rect 55496 32240 55548 32292
rect 53104 32215 53156 32224
rect 53104 32181 53113 32215
rect 53113 32181 53147 32215
rect 53147 32181 53156 32215
rect 53104 32172 53156 32181
rect 55036 32215 55088 32224
rect 55036 32181 55045 32215
rect 55045 32181 55079 32215
rect 55079 32181 55088 32215
rect 55036 32172 55088 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2872 31968 2924 32020
rect 3424 31968 3476 32020
rect 3516 31968 3568 32020
rect 4620 31968 4672 32020
rect 4988 32011 5040 32020
rect 4988 31977 4997 32011
rect 4997 31977 5031 32011
rect 5031 31977 5040 32011
rect 4988 31968 5040 31977
rect 6368 31968 6420 32020
rect 6920 31968 6972 32020
rect 7840 31968 7892 32020
rect 2504 31832 2556 31884
rect 3332 31764 3384 31816
rect 4988 31832 5040 31884
rect 4896 31764 4948 31816
rect 5264 31764 5316 31816
rect 10232 31968 10284 32020
rect 37740 31900 37792 31952
rect 6460 31764 6512 31816
rect 38844 31875 38896 31884
rect 38844 31841 38853 31875
rect 38853 31841 38887 31875
rect 38887 31841 38896 31875
rect 38844 31832 38896 31841
rect 4344 31696 4396 31748
rect 5356 31696 5408 31748
rect 6276 31696 6328 31748
rect 7196 31696 7248 31748
rect 10600 31764 10652 31816
rect 36268 31807 36320 31816
rect 36268 31773 36277 31807
rect 36277 31773 36311 31807
rect 36311 31773 36320 31807
rect 36268 31764 36320 31773
rect 38384 31764 38436 31816
rect 39396 31968 39448 32020
rect 40592 31968 40644 32020
rect 42064 32011 42116 32020
rect 42064 31977 42073 32011
rect 42073 31977 42107 32011
rect 42107 31977 42116 32011
rect 42064 31968 42116 31977
rect 43076 31968 43128 32020
rect 40040 31832 40092 31884
rect 41236 31832 41288 31884
rect 41604 31875 41656 31884
rect 41604 31841 41613 31875
rect 41613 31841 41647 31875
rect 41647 31841 41656 31875
rect 41604 31832 41656 31841
rect 43352 31900 43404 31952
rect 10416 31696 10468 31748
rect 13452 31696 13504 31748
rect 36728 31739 36780 31748
rect 36728 31705 36737 31739
rect 36737 31705 36771 31739
rect 36771 31705 36780 31739
rect 36728 31696 36780 31705
rect 39948 31764 40000 31816
rect 3516 31671 3568 31680
rect 3516 31637 3525 31671
rect 3525 31637 3559 31671
rect 3559 31637 3568 31671
rect 3516 31628 3568 31637
rect 4068 31628 4120 31680
rect 10140 31628 10192 31680
rect 11704 31628 11756 31680
rect 38476 31628 38528 31680
rect 38660 31671 38712 31680
rect 38660 31637 38669 31671
rect 38669 31637 38703 31671
rect 38703 31637 38712 31671
rect 39396 31739 39448 31748
rect 39396 31705 39405 31739
rect 39405 31705 39439 31739
rect 39439 31705 39448 31739
rect 39396 31696 39448 31705
rect 41420 31696 41472 31748
rect 43628 31807 43680 31816
rect 43628 31773 43637 31807
rect 43637 31773 43671 31807
rect 43671 31773 43680 31807
rect 43628 31764 43680 31773
rect 44180 31900 44232 31952
rect 44640 31968 44692 32020
rect 47032 31968 47084 32020
rect 47124 31968 47176 32020
rect 48596 31968 48648 32020
rect 44548 31900 44600 31952
rect 38660 31628 38712 31637
rect 42892 31628 42944 31680
rect 44640 31764 44692 31816
rect 45652 31807 45704 31816
rect 45652 31773 45661 31807
rect 45661 31773 45695 31807
rect 45695 31773 45704 31807
rect 45652 31764 45704 31773
rect 46756 31807 46808 31816
rect 46756 31773 46765 31807
rect 46765 31773 46799 31807
rect 46799 31773 46808 31807
rect 46756 31764 46808 31773
rect 47308 31807 47360 31816
rect 44364 31696 44416 31748
rect 45192 31696 45244 31748
rect 47308 31773 47317 31807
rect 47317 31773 47351 31807
rect 47351 31773 47360 31807
rect 47308 31764 47360 31773
rect 48320 31900 48372 31952
rect 49056 31900 49108 31952
rect 48964 31875 49016 31884
rect 48964 31841 48973 31875
rect 48973 31841 49007 31875
rect 49007 31841 49016 31875
rect 48964 31832 49016 31841
rect 51080 31968 51132 32020
rect 54392 31968 54444 32020
rect 55588 31968 55640 32020
rect 50896 31900 50948 31952
rect 52552 31900 52604 31952
rect 47676 31696 47728 31748
rect 49516 31807 49568 31816
rect 49516 31773 49525 31807
rect 49525 31773 49559 31807
rect 49559 31773 49568 31807
rect 49516 31764 49568 31773
rect 49792 31807 49844 31816
rect 49792 31773 49801 31807
rect 49801 31773 49835 31807
rect 49835 31773 49844 31807
rect 49792 31764 49844 31773
rect 51448 31764 51500 31816
rect 52092 31807 52144 31816
rect 52092 31773 52101 31807
rect 52101 31773 52135 31807
rect 52135 31773 52144 31807
rect 52092 31764 52144 31773
rect 52460 31832 52512 31884
rect 53012 31696 53064 31748
rect 55128 31807 55180 31816
rect 55128 31773 55137 31807
rect 55137 31773 55171 31807
rect 55171 31773 55180 31807
rect 55128 31764 55180 31773
rect 56508 31764 56560 31816
rect 58900 31764 58952 31816
rect 55220 31696 55272 31748
rect 56876 31696 56928 31748
rect 46940 31628 46992 31680
rect 47032 31628 47084 31680
rect 47216 31628 47268 31680
rect 48964 31628 49016 31680
rect 49240 31671 49292 31680
rect 49240 31637 49249 31671
rect 49249 31637 49283 31671
rect 49283 31637 49292 31671
rect 49240 31628 49292 31637
rect 54852 31628 54904 31680
rect 56692 31671 56744 31680
rect 56692 31637 56701 31671
rect 56701 31637 56735 31671
rect 56735 31637 56744 31671
rect 56692 31628 56744 31637
rect 58164 31671 58216 31680
rect 58164 31637 58173 31671
rect 58173 31637 58207 31671
rect 58207 31637 58216 31671
rect 58164 31628 58216 31637
rect 58348 31671 58400 31680
rect 58348 31637 58357 31671
rect 58357 31637 58391 31671
rect 58391 31637 58400 31671
rect 58348 31628 58400 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 4896 31467 4948 31476
rect 4896 31433 4905 31467
rect 4905 31433 4939 31467
rect 4939 31433 4948 31467
rect 4896 31424 4948 31433
rect 5632 31424 5684 31476
rect 8392 31424 8444 31476
rect 2688 31331 2740 31340
rect 2688 31297 2697 31331
rect 2697 31297 2731 31331
rect 2731 31297 2740 31331
rect 2688 31288 2740 31297
rect 3884 31331 3936 31340
rect 3884 31297 3893 31331
rect 3893 31297 3927 31331
rect 3927 31297 3936 31331
rect 3884 31288 3936 31297
rect 4988 31356 5040 31408
rect 9036 31356 9088 31408
rect 36728 31424 36780 31476
rect 38660 31424 38712 31476
rect 38844 31424 38896 31476
rect 39488 31424 39540 31476
rect 10048 31356 10100 31408
rect 4160 31331 4212 31340
rect 4160 31297 4169 31331
rect 4169 31297 4203 31331
rect 4203 31297 4212 31331
rect 4160 31288 4212 31297
rect 4344 31331 4396 31340
rect 4344 31297 4353 31331
rect 4353 31297 4387 31331
rect 4387 31297 4396 31331
rect 4344 31288 4396 31297
rect 5172 31288 5224 31340
rect 940 31220 992 31272
rect 3700 31263 3752 31272
rect 3700 31229 3709 31263
rect 3709 31229 3743 31263
rect 3743 31229 3752 31263
rect 3700 31220 3752 31229
rect 3792 31220 3844 31272
rect 6092 31288 6144 31340
rect 6276 31288 6328 31340
rect 5816 31220 5868 31272
rect 6920 31331 6972 31340
rect 6920 31297 6929 31331
rect 6929 31297 6963 31331
rect 6963 31297 6972 31331
rect 6920 31288 6972 31297
rect 7104 31288 7156 31340
rect 8484 31331 8536 31340
rect 8484 31297 8493 31331
rect 8493 31297 8527 31331
rect 8527 31297 8536 31331
rect 8484 31288 8536 31297
rect 8760 31331 8812 31340
rect 8760 31297 8769 31331
rect 8769 31297 8803 31331
rect 8803 31297 8812 31331
rect 8760 31288 8812 31297
rect 10968 31288 11020 31340
rect 11520 31288 11572 31340
rect 12532 31288 12584 31340
rect 37740 31288 37792 31340
rect 38200 31331 38252 31340
rect 38200 31297 38209 31331
rect 38209 31297 38243 31331
rect 38243 31297 38252 31331
rect 38200 31288 38252 31297
rect 38476 31331 38528 31340
rect 38476 31297 38485 31331
rect 38485 31297 38519 31331
rect 38519 31297 38528 31331
rect 38476 31288 38528 31297
rect 38660 31288 38712 31340
rect 39028 31288 39080 31340
rect 39396 31331 39448 31340
rect 39396 31297 39405 31331
rect 39405 31297 39439 31331
rect 39439 31297 39448 31331
rect 39396 31288 39448 31297
rect 40224 31331 40276 31340
rect 40224 31297 40233 31331
rect 40233 31297 40267 31331
rect 40267 31297 40276 31331
rect 40224 31288 40276 31297
rect 5908 31152 5960 31204
rect 6368 31152 6420 31204
rect 8852 31152 8904 31204
rect 13452 31263 13504 31272
rect 13452 31229 13461 31263
rect 13461 31229 13495 31263
rect 13495 31229 13504 31263
rect 13452 31220 13504 31229
rect 15844 31220 15896 31272
rect 39120 31152 39172 31204
rect 39396 31152 39448 31204
rect 45560 31424 45612 31476
rect 45192 31288 45244 31340
rect 41604 31220 41656 31272
rect 42524 31220 42576 31272
rect 44088 31263 44140 31272
rect 44088 31229 44097 31263
rect 44097 31229 44131 31263
rect 44131 31229 44140 31263
rect 44088 31220 44140 31229
rect 43168 31152 43220 31204
rect 3148 31127 3200 31136
rect 3148 31093 3157 31127
rect 3157 31093 3191 31127
rect 3191 31093 3200 31127
rect 3148 31084 3200 31093
rect 3424 31084 3476 31136
rect 4620 31084 4672 31136
rect 7196 31127 7248 31136
rect 7196 31093 7205 31127
rect 7205 31093 7239 31127
rect 7239 31093 7248 31127
rect 7196 31084 7248 31093
rect 8484 31084 8536 31136
rect 8760 31084 8812 31136
rect 8944 31084 8996 31136
rect 9680 31084 9732 31136
rect 40132 31084 40184 31136
rect 47032 31424 47084 31476
rect 47124 31424 47176 31476
rect 49240 31424 49292 31476
rect 52460 31467 52512 31476
rect 52460 31433 52469 31467
rect 52469 31433 52503 31467
rect 52503 31433 52512 31467
rect 52460 31424 52512 31433
rect 53012 31424 53064 31476
rect 55220 31424 55272 31476
rect 56876 31424 56928 31476
rect 46204 31356 46256 31408
rect 45836 31263 45888 31272
rect 45836 31229 45845 31263
rect 45845 31229 45879 31263
rect 45879 31229 45888 31263
rect 45836 31220 45888 31229
rect 46756 31220 46808 31272
rect 48320 31331 48372 31340
rect 48320 31297 48329 31331
rect 48329 31297 48363 31331
rect 48363 31297 48372 31331
rect 48320 31288 48372 31297
rect 51080 31331 51132 31340
rect 51080 31297 51089 31331
rect 51089 31297 51123 31331
rect 51123 31297 51132 31331
rect 51080 31288 51132 31297
rect 52920 31356 52972 31408
rect 53748 31356 53800 31408
rect 54852 31356 54904 31408
rect 48872 31263 48924 31272
rect 48872 31229 48881 31263
rect 48881 31229 48915 31263
rect 48915 31229 48924 31263
rect 48872 31220 48924 31229
rect 51816 31263 51868 31272
rect 51816 31229 51825 31263
rect 51825 31229 51859 31263
rect 51859 31229 51868 31263
rect 51816 31220 51868 31229
rect 53104 31263 53156 31272
rect 53104 31229 53113 31263
rect 53113 31229 53147 31263
rect 53147 31229 53156 31263
rect 53104 31220 53156 31229
rect 55128 31288 55180 31340
rect 56968 31356 57020 31408
rect 54944 31263 54996 31272
rect 54944 31229 54953 31263
rect 54953 31229 54987 31263
rect 54987 31229 54996 31263
rect 54944 31220 54996 31229
rect 57336 31288 57388 31340
rect 58164 31288 58216 31340
rect 56692 31220 56744 31272
rect 45744 31084 45796 31136
rect 45928 31127 45980 31136
rect 45928 31093 45937 31127
rect 45937 31093 45971 31127
rect 45971 31093 45980 31127
rect 45928 31084 45980 31093
rect 47124 31084 47176 31136
rect 48412 31084 48464 31136
rect 48504 31084 48556 31136
rect 48688 31127 48740 31136
rect 48688 31093 48697 31127
rect 48697 31093 48731 31127
rect 48731 31093 48740 31127
rect 48688 31084 48740 31093
rect 48780 31127 48832 31136
rect 48780 31093 48789 31127
rect 48789 31093 48823 31127
rect 48823 31093 48832 31127
rect 48780 31084 48832 31093
rect 49516 31084 49568 31136
rect 51356 31084 51408 31136
rect 51724 31127 51776 31136
rect 51724 31093 51733 31127
rect 51733 31093 51767 31127
rect 51767 31093 51776 31127
rect 51724 31084 51776 31093
rect 52552 31084 52604 31136
rect 54484 31127 54536 31136
rect 54484 31093 54493 31127
rect 54493 31093 54527 31127
rect 54527 31093 54536 31127
rect 54484 31084 54536 31093
rect 54852 31152 54904 31204
rect 56140 31084 56192 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 3148 30880 3200 30932
rect 3700 30880 3752 30932
rect 7012 30880 7064 30932
rect 8300 30880 8352 30932
rect 9220 30880 9272 30932
rect 10140 30880 10192 30932
rect 38200 30880 38252 30932
rect 38660 30923 38712 30932
rect 38660 30889 38669 30923
rect 38669 30889 38703 30923
rect 38703 30889 38712 30923
rect 38660 30880 38712 30889
rect 39948 30923 40000 30932
rect 39948 30889 39957 30923
rect 39957 30889 39991 30923
rect 39991 30889 40000 30923
rect 39948 30880 40000 30889
rect 44088 30880 44140 30932
rect 9680 30812 9732 30864
rect 11704 30812 11756 30864
rect 3148 30787 3200 30796
rect 3148 30753 3157 30787
rect 3157 30753 3191 30787
rect 3191 30753 3200 30787
rect 3148 30744 3200 30753
rect 3424 30744 3476 30796
rect 4620 30744 4672 30796
rect 8208 30744 8260 30796
rect 3332 30719 3384 30728
rect 3332 30685 3341 30719
rect 3341 30685 3375 30719
rect 3375 30685 3384 30719
rect 3332 30676 3384 30685
rect 3884 30676 3936 30728
rect 2412 30608 2464 30660
rect 5080 30608 5132 30660
rect 2688 30540 2740 30592
rect 5816 30676 5868 30728
rect 6368 30676 6420 30728
rect 7472 30676 7524 30728
rect 8944 30719 8996 30728
rect 8944 30685 8953 30719
rect 8953 30685 8987 30719
rect 8987 30685 8996 30719
rect 8944 30676 8996 30685
rect 39580 30744 39632 30796
rect 41328 30787 41380 30796
rect 41328 30753 41337 30787
rect 41337 30753 41371 30787
rect 41371 30753 41380 30787
rect 41328 30744 41380 30753
rect 41972 30744 42024 30796
rect 9772 30608 9824 30660
rect 38844 30676 38896 30728
rect 40040 30719 40092 30728
rect 40040 30685 40049 30719
rect 40049 30685 40083 30719
rect 40083 30685 40092 30719
rect 40040 30676 40092 30685
rect 40132 30719 40184 30728
rect 40132 30685 40141 30719
rect 40141 30685 40175 30719
rect 40175 30685 40184 30719
rect 40132 30676 40184 30685
rect 42984 30719 43036 30728
rect 42984 30685 42993 30719
rect 42993 30685 43027 30719
rect 43027 30685 43036 30719
rect 42984 30676 43036 30685
rect 43168 30676 43220 30728
rect 43720 30719 43772 30728
rect 43720 30685 43729 30719
rect 43729 30685 43763 30719
rect 43763 30685 43772 30719
rect 43720 30676 43772 30685
rect 45928 30880 45980 30932
rect 48504 30923 48556 30932
rect 48504 30889 48513 30923
rect 48513 30889 48547 30923
rect 48547 30889 48556 30923
rect 48504 30880 48556 30889
rect 48780 30880 48832 30932
rect 45744 30855 45796 30864
rect 45744 30821 45753 30855
rect 45753 30821 45787 30855
rect 45787 30821 45796 30855
rect 45744 30812 45796 30821
rect 45836 30744 45888 30796
rect 10048 30608 10100 30660
rect 13728 30608 13780 30660
rect 5448 30540 5500 30592
rect 6184 30583 6236 30592
rect 6184 30549 6193 30583
rect 6193 30549 6227 30583
rect 6227 30549 6236 30583
rect 6184 30540 6236 30549
rect 6368 30540 6420 30592
rect 6736 30540 6788 30592
rect 9312 30540 9364 30592
rect 9864 30583 9916 30592
rect 9864 30549 9873 30583
rect 9873 30549 9907 30583
rect 9907 30549 9916 30583
rect 9864 30540 9916 30549
rect 9956 30540 10008 30592
rect 10324 30583 10376 30592
rect 10324 30549 10333 30583
rect 10333 30549 10367 30583
rect 10367 30549 10376 30583
rect 10324 30540 10376 30549
rect 10600 30540 10652 30592
rect 12900 30540 12952 30592
rect 17132 30608 17184 30660
rect 38292 30651 38344 30660
rect 38292 30617 38301 30651
rect 38301 30617 38335 30651
rect 38335 30617 38344 30651
rect 38292 30608 38344 30617
rect 42800 30608 42852 30660
rect 45560 30719 45612 30728
rect 45560 30685 45569 30719
rect 45569 30685 45603 30719
rect 45603 30685 45612 30719
rect 45560 30676 45612 30685
rect 45652 30676 45704 30728
rect 47400 30744 47452 30796
rect 51816 30880 51868 30932
rect 54484 30880 54536 30932
rect 56968 30880 57020 30932
rect 57336 30880 57388 30932
rect 51724 30744 51776 30796
rect 36268 30540 36320 30592
rect 43076 30583 43128 30592
rect 43076 30549 43085 30583
rect 43085 30549 43119 30583
rect 43119 30549 43128 30583
rect 43076 30540 43128 30549
rect 45744 30651 45796 30660
rect 45744 30617 45753 30651
rect 45753 30617 45787 30651
rect 45787 30617 45796 30651
rect 45744 30608 45796 30617
rect 47216 30608 47268 30660
rect 51172 30608 51224 30660
rect 53104 30719 53156 30728
rect 53104 30685 53113 30719
rect 53113 30685 53147 30719
rect 53147 30685 53156 30719
rect 53104 30676 53156 30685
rect 58624 30744 58676 30796
rect 51816 30608 51868 30660
rect 58348 30719 58400 30728
rect 58348 30685 58357 30719
rect 58357 30685 58391 30719
rect 58391 30685 58400 30719
rect 58348 30676 58400 30685
rect 46664 30540 46716 30592
rect 47308 30540 47360 30592
rect 50160 30540 50212 30592
rect 51632 30540 51684 30592
rect 53472 30583 53524 30592
rect 53472 30549 53481 30583
rect 53481 30549 53515 30583
rect 53515 30549 53524 30583
rect 53472 30540 53524 30549
rect 54300 30583 54352 30592
rect 54300 30549 54309 30583
rect 54309 30549 54343 30583
rect 54343 30549 54352 30583
rect 54300 30540 54352 30549
rect 57244 30583 57296 30592
rect 57244 30549 57253 30583
rect 57253 30549 57287 30583
rect 57287 30549 57296 30583
rect 57244 30540 57296 30549
rect 57612 30540 57664 30592
rect 58072 30583 58124 30592
rect 58072 30549 58081 30583
rect 58081 30549 58115 30583
rect 58115 30549 58124 30583
rect 58072 30540 58124 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 4068 30336 4120 30388
rect 3148 30268 3200 30320
rect 5908 30336 5960 30388
rect 9864 30336 9916 30388
rect 10324 30336 10376 30388
rect 2688 30243 2740 30252
rect 2688 30209 2697 30243
rect 2697 30209 2731 30243
rect 2731 30209 2740 30243
rect 2688 30200 2740 30209
rect 4068 30200 4120 30252
rect 3700 30175 3752 30184
rect 3700 30141 3709 30175
rect 3709 30141 3743 30175
rect 3743 30141 3752 30175
rect 3700 30132 3752 30141
rect 3332 30064 3384 30116
rect 5172 30200 5224 30252
rect 5356 30243 5408 30252
rect 5356 30209 5365 30243
rect 5365 30209 5399 30243
rect 5399 30209 5408 30243
rect 5356 30200 5408 30209
rect 5540 30243 5592 30252
rect 5540 30209 5549 30243
rect 5549 30209 5583 30243
rect 5583 30209 5592 30243
rect 5540 30200 5592 30209
rect 6828 30268 6880 30320
rect 5632 30064 5684 30116
rect 3608 30039 3660 30048
rect 3608 30005 3617 30039
rect 3617 30005 3651 30039
rect 3651 30005 3660 30039
rect 3608 29996 3660 30005
rect 4896 29996 4948 30048
rect 6184 30200 6236 30252
rect 6644 30243 6696 30252
rect 6644 30209 6678 30243
rect 6678 30209 6696 30243
rect 6644 30200 6696 30209
rect 10600 30268 10652 30320
rect 10692 30200 10744 30252
rect 11060 30336 11112 30388
rect 10968 30268 11020 30320
rect 12624 30268 12676 30320
rect 40040 30336 40092 30388
rect 43076 30336 43128 30388
rect 43720 30379 43772 30388
rect 43720 30345 43729 30379
rect 43729 30345 43763 30379
rect 43763 30345 43772 30379
rect 43720 30336 43772 30345
rect 45744 30336 45796 30388
rect 46572 30336 46624 30388
rect 10876 30233 10928 30242
rect 10876 30199 10885 30233
rect 10885 30199 10919 30233
rect 10919 30199 10928 30233
rect 10876 30190 10928 30199
rect 41420 30268 41472 30320
rect 10416 30107 10468 30116
rect 10416 30073 10425 30107
rect 10425 30073 10459 30107
rect 10459 30073 10468 30107
rect 10416 30064 10468 30073
rect 39212 30243 39264 30252
rect 39212 30209 39221 30243
rect 39221 30209 39255 30243
rect 39255 30209 39264 30243
rect 39212 30200 39264 30209
rect 39396 30243 39448 30252
rect 39396 30209 39405 30243
rect 39405 30209 39439 30243
rect 39439 30209 39448 30243
rect 39396 30200 39448 30209
rect 39488 30200 39540 30252
rect 40408 30200 40460 30252
rect 42800 30200 42852 30252
rect 43352 30243 43404 30252
rect 43352 30209 43361 30243
rect 43361 30209 43395 30243
rect 43395 30209 43404 30243
rect 43352 30200 43404 30209
rect 47308 30268 47360 30320
rect 11520 30175 11572 30184
rect 11520 30141 11529 30175
rect 11529 30141 11563 30175
rect 11563 30141 11572 30175
rect 11520 30132 11572 30141
rect 15384 30132 15436 30184
rect 7472 29996 7524 30048
rect 9220 29996 9272 30048
rect 31024 30064 31076 30116
rect 11060 29996 11112 30048
rect 37372 30064 37424 30116
rect 38292 30064 38344 30116
rect 38660 29996 38712 30048
rect 38936 29996 38988 30048
rect 39764 29996 39816 30048
rect 41972 30132 42024 30184
rect 42524 30132 42576 30184
rect 43996 30132 44048 30184
rect 44180 30243 44232 30252
rect 44180 30209 44189 30243
rect 44189 30209 44223 30243
rect 44223 30209 44232 30243
rect 44180 30200 44232 30209
rect 43444 29996 43496 30048
rect 43536 30039 43588 30048
rect 43536 30005 43545 30039
rect 43545 30005 43579 30039
rect 43579 30005 43588 30039
rect 43536 29996 43588 30005
rect 45100 30039 45152 30048
rect 45100 30005 45109 30039
rect 45109 30005 45143 30039
rect 45143 30005 45152 30039
rect 48412 30243 48464 30252
rect 48412 30209 48421 30243
rect 48421 30209 48455 30243
rect 48455 30209 48464 30243
rect 48412 30200 48464 30209
rect 48964 30268 49016 30320
rect 49608 30336 49660 30388
rect 50160 30268 50212 30320
rect 51724 30336 51776 30388
rect 53472 30336 53524 30388
rect 45744 30132 45796 30184
rect 47032 30175 47084 30184
rect 47032 30141 47041 30175
rect 47041 30141 47075 30175
rect 47075 30141 47084 30175
rect 47032 30132 47084 30141
rect 46020 30064 46072 30116
rect 45100 29996 45152 30005
rect 45744 29996 45796 30048
rect 47860 30039 47912 30048
rect 47860 30005 47869 30039
rect 47869 30005 47903 30039
rect 47903 30005 47912 30039
rect 47860 29996 47912 30005
rect 51632 30249 51684 30252
rect 51632 30215 51641 30249
rect 51641 30215 51675 30249
rect 51675 30215 51684 30249
rect 51632 30200 51684 30215
rect 51816 30132 51868 30184
rect 52092 30243 52144 30252
rect 52092 30209 52101 30243
rect 52101 30209 52135 30243
rect 52135 30209 52144 30243
rect 52092 30200 52144 30209
rect 52920 30243 52972 30252
rect 52920 30209 52929 30243
rect 52929 30209 52963 30243
rect 52963 30209 52972 30243
rect 52920 30200 52972 30209
rect 53196 30200 53248 30252
rect 53564 30268 53616 30320
rect 57796 30336 57848 30388
rect 54300 30243 54352 30252
rect 54300 30209 54309 30243
rect 54309 30209 54343 30243
rect 54343 30209 54352 30243
rect 54300 30200 54352 30209
rect 54668 30200 54720 30252
rect 54852 30268 54904 30320
rect 55220 30243 55272 30252
rect 55220 30209 55229 30243
rect 55229 30209 55263 30243
rect 55263 30209 55272 30243
rect 55220 30200 55272 30209
rect 57520 30243 57572 30252
rect 57520 30209 57529 30243
rect 57529 30209 57563 30243
rect 57563 30209 57572 30243
rect 57520 30200 57572 30209
rect 54576 30132 54628 30184
rect 58072 30200 58124 30252
rect 58532 30200 58584 30252
rect 52092 30064 52144 30116
rect 58624 30064 58676 30116
rect 51908 29996 51960 30048
rect 52000 29996 52052 30048
rect 52184 29996 52236 30048
rect 53380 30039 53432 30048
rect 53380 30005 53389 30039
rect 53389 30005 53423 30039
rect 53423 30005 53432 30039
rect 53380 29996 53432 30005
rect 54392 30039 54444 30048
rect 54392 30005 54401 30039
rect 54401 30005 54435 30039
rect 54435 30005 54444 30039
rect 54392 29996 54444 30005
rect 54668 29996 54720 30048
rect 55864 30039 55916 30048
rect 55864 30005 55873 30039
rect 55873 30005 55907 30039
rect 55907 30005 55916 30039
rect 55864 29996 55916 30005
rect 58072 30039 58124 30048
rect 58072 30005 58081 30039
rect 58081 30005 58115 30039
rect 58115 30005 58124 30039
rect 58072 29996 58124 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 3608 29792 3660 29844
rect 3700 29792 3752 29844
rect 4068 29792 4120 29844
rect 5080 29792 5132 29844
rect 5908 29792 5960 29844
rect 6644 29792 6696 29844
rect 6736 29792 6788 29844
rect 15844 29835 15896 29844
rect 15844 29801 15853 29835
rect 15853 29801 15887 29835
rect 15887 29801 15896 29835
rect 15844 29792 15896 29801
rect 5172 29724 5224 29776
rect 940 29520 992 29572
rect 1400 29452 1452 29504
rect 4896 29656 4948 29708
rect 6736 29656 6788 29708
rect 9128 29699 9180 29708
rect 9128 29665 9137 29699
rect 9137 29665 9171 29699
rect 9171 29665 9180 29699
rect 9128 29656 9180 29665
rect 4804 29520 4856 29572
rect 2964 29495 3016 29504
rect 2964 29461 2973 29495
rect 2973 29461 3007 29495
rect 3007 29461 3016 29495
rect 2964 29452 3016 29461
rect 3148 29452 3200 29504
rect 5816 29520 5868 29572
rect 6552 29563 6604 29572
rect 6552 29529 6561 29563
rect 6561 29529 6595 29563
rect 6595 29529 6604 29563
rect 6552 29520 6604 29529
rect 8944 29588 8996 29640
rect 10232 29724 10284 29776
rect 15016 29724 15068 29776
rect 31024 29792 31076 29844
rect 39948 29792 40000 29844
rect 41328 29792 41380 29844
rect 9772 29588 9824 29640
rect 9956 29520 10008 29572
rect 10876 29588 10928 29640
rect 15844 29656 15896 29708
rect 38660 29724 38712 29776
rect 43536 29792 43588 29844
rect 44180 29792 44232 29844
rect 11888 29631 11940 29640
rect 11888 29597 11897 29631
rect 11897 29597 11931 29631
rect 11931 29597 11940 29631
rect 11888 29588 11940 29597
rect 11612 29520 11664 29572
rect 12440 29563 12492 29572
rect 12440 29529 12449 29563
rect 12449 29529 12483 29563
rect 12483 29529 12492 29563
rect 36268 29656 36320 29708
rect 37188 29656 37240 29708
rect 39396 29656 39448 29708
rect 39580 29699 39632 29708
rect 39580 29665 39589 29699
rect 39589 29665 39623 29699
rect 39623 29665 39632 29699
rect 39580 29656 39632 29665
rect 40040 29656 40092 29708
rect 39764 29588 39816 29640
rect 41972 29631 42024 29640
rect 41972 29597 41981 29631
rect 41981 29597 42015 29631
rect 42015 29597 42024 29631
rect 41972 29588 42024 29597
rect 43444 29724 43496 29776
rect 47032 29792 47084 29844
rect 47124 29792 47176 29844
rect 51816 29792 51868 29844
rect 52092 29792 52144 29844
rect 53196 29792 53248 29844
rect 53380 29792 53432 29844
rect 55220 29792 55272 29844
rect 56508 29792 56560 29844
rect 45652 29656 45704 29708
rect 42524 29588 42576 29640
rect 12440 29520 12492 29529
rect 37648 29563 37700 29572
rect 37648 29529 37657 29563
rect 37657 29529 37691 29563
rect 37691 29529 37700 29563
rect 37648 29520 37700 29529
rect 40960 29520 41012 29572
rect 41420 29520 41472 29572
rect 6736 29495 6788 29504
rect 6736 29461 6745 29495
rect 6745 29461 6779 29495
rect 6779 29461 6788 29495
rect 6736 29452 6788 29461
rect 6920 29452 6972 29504
rect 7472 29452 7524 29504
rect 11152 29452 11204 29504
rect 15384 29495 15436 29504
rect 15384 29461 15393 29495
rect 15393 29461 15427 29495
rect 15427 29461 15436 29495
rect 15384 29452 15436 29461
rect 37464 29452 37516 29504
rect 38936 29452 38988 29504
rect 39488 29452 39540 29504
rect 39580 29452 39632 29504
rect 40040 29452 40092 29504
rect 43996 29588 44048 29640
rect 44824 29588 44876 29640
rect 43628 29520 43680 29572
rect 44548 29520 44600 29572
rect 43536 29452 43588 29504
rect 46572 29588 46624 29640
rect 50160 29767 50212 29776
rect 50160 29733 50169 29767
rect 50169 29733 50203 29767
rect 50203 29733 50212 29767
rect 50160 29724 50212 29733
rect 52000 29724 52052 29776
rect 47400 29656 47452 29708
rect 47860 29656 47912 29708
rect 48964 29656 49016 29708
rect 50620 29656 50672 29708
rect 47308 29588 47360 29640
rect 49976 29588 50028 29640
rect 51080 29631 51132 29640
rect 51080 29597 51089 29631
rect 51089 29597 51123 29631
rect 51123 29597 51132 29631
rect 51080 29588 51132 29597
rect 51448 29631 51500 29640
rect 51448 29597 51457 29631
rect 51457 29597 51491 29631
rect 51491 29597 51500 29631
rect 51448 29588 51500 29597
rect 51816 29588 51868 29640
rect 51356 29563 51408 29572
rect 51356 29529 51365 29563
rect 51365 29529 51399 29563
rect 51399 29529 51408 29563
rect 51356 29520 51408 29529
rect 51540 29520 51592 29572
rect 46572 29452 46624 29504
rect 46848 29452 46900 29504
rect 49240 29495 49292 29504
rect 49240 29461 49249 29495
rect 49249 29461 49283 29495
rect 49283 29461 49292 29495
rect 49240 29452 49292 29461
rect 49424 29452 49476 29504
rect 52184 29631 52236 29640
rect 52184 29597 52193 29631
rect 52193 29597 52227 29631
rect 52227 29597 52236 29631
rect 52184 29588 52236 29597
rect 52460 29631 52512 29640
rect 52460 29597 52469 29631
rect 52469 29597 52503 29631
rect 52503 29597 52512 29631
rect 52460 29588 52512 29597
rect 54392 29656 54444 29708
rect 55036 29656 55088 29708
rect 57520 29835 57572 29844
rect 57520 29801 57529 29835
rect 57529 29801 57563 29835
rect 57563 29801 57572 29835
rect 57520 29792 57572 29801
rect 58716 29724 58768 29776
rect 53564 29631 53616 29640
rect 53564 29597 53573 29631
rect 53573 29597 53607 29631
rect 53607 29597 53616 29631
rect 53564 29588 53616 29597
rect 55128 29631 55180 29640
rect 55128 29597 55137 29631
rect 55137 29597 55171 29631
rect 55171 29597 55180 29631
rect 55128 29588 55180 29597
rect 56968 29631 57020 29640
rect 53840 29520 53892 29572
rect 56968 29597 56977 29631
rect 56977 29597 57011 29631
rect 57011 29597 57020 29631
rect 56968 29588 57020 29597
rect 56048 29520 56100 29572
rect 57244 29588 57296 29640
rect 52276 29495 52328 29504
rect 52276 29461 52285 29495
rect 52285 29461 52319 29495
rect 52319 29461 52328 29495
rect 52276 29452 52328 29461
rect 53012 29452 53064 29504
rect 53564 29452 53616 29504
rect 55312 29495 55364 29504
rect 55312 29461 55321 29495
rect 55321 29461 55355 29495
rect 55355 29461 55364 29495
rect 55312 29452 55364 29461
rect 55404 29452 55456 29504
rect 57060 29495 57112 29504
rect 57060 29461 57069 29495
rect 57069 29461 57103 29495
rect 57103 29461 57112 29495
rect 57060 29452 57112 29461
rect 57796 29588 57848 29640
rect 57612 29520 57664 29572
rect 58532 29452 58584 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 1400 29291 1452 29300
rect 1400 29257 1409 29291
rect 1409 29257 1443 29291
rect 1443 29257 1452 29291
rect 1400 29248 1452 29257
rect 2412 29180 2464 29232
rect 2964 29180 3016 29232
rect 3240 29112 3292 29164
rect 5448 29248 5500 29300
rect 6460 29248 6512 29300
rect 6736 29248 6788 29300
rect 8944 29291 8996 29300
rect 8944 29257 8953 29291
rect 8953 29257 8987 29291
rect 8987 29257 8996 29291
rect 8944 29248 8996 29257
rect 4712 29223 4764 29232
rect 4712 29189 4746 29223
rect 4746 29189 4764 29223
rect 4712 29180 4764 29189
rect 6276 29180 6328 29232
rect 4988 29112 5040 29164
rect 5908 29112 5960 29164
rect 6920 29180 6972 29232
rect 9956 29180 10008 29232
rect 10968 29223 11020 29232
rect 10968 29189 10977 29223
rect 10977 29189 11011 29223
rect 11011 29189 11020 29223
rect 10968 29180 11020 29189
rect 11060 29180 11112 29232
rect 11612 29291 11664 29300
rect 11612 29257 11621 29291
rect 11621 29257 11655 29291
rect 11655 29257 11664 29291
rect 11612 29248 11664 29257
rect 15016 29248 15068 29300
rect 11428 29180 11480 29232
rect 10508 29155 10560 29164
rect 10508 29121 10517 29155
rect 10517 29121 10551 29155
rect 10551 29121 10560 29155
rect 10508 29112 10560 29121
rect 10600 29155 10652 29164
rect 10600 29121 10609 29155
rect 10609 29121 10643 29155
rect 10643 29121 10652 29155
rect 10600 29112 10652 29121
rect 10692 29112 10744 29164
rect 4252 29044 4304 29096
rect 5632 29044 5684 29096
rect 6828 29044 6880 29096
rect 7196 28976 7248 29028
rect 11060 29044 11112 29096
rect 37188 29248 37240 29300
rect 37648 29180 37700 29232
rect 37372 29155 37424 29164
rect 37372 29121 37381 29155
rect 37381 29121 37415 29155
rect 37415 29121 37424 29155
rect 37372 29112 37424 29121
rect 39212 29155 39264 29164
rect 39212 29121 39221 29155
rect 39221 29121 39255 29155
rect 39255 29121 39264 29155
rect 39212 29112 39264 29121
rect 3608 28908 3660 28960
rect 4620 28908 4672 28960
rect 9312 28908 9364 28960
rect 11520 28976 11572 29028
rect 37832 29044 37884 29096
rect 37464 29019 37516 29028
rect 37464 28985 37473 29019
rect 37473 28985 37507 29019
rect 37507 28985 37516 29019
rect 37464 28976 37516 28985
rect 39028 29087 39080 29096
rect 39028 29053 39037 29087
rect 39037 29053 39071 29087
rect 39071 29053 39080 29087
rect 39028 29044 39080 29053
rect 38660 28976 38712 29028
rect 40132 29248 40184 29300
rect 45100 29248 45152 29300
rect 45652 29248 45704 29300
rect 46848 29248 46900 29300
rect 48688 29248 48740 29300
rect 49240 29248 49292 29300
rect 52460 29248 52512 29300
rect 52552 29248 52604 29300
rect 53012 29291 53064 29300
rect 53012 29257 53021 29291
rect 53021 29257 53055 29291
rect 53055 29257 53064 29291
rect 53012 29248 53064 29257
rect 40960 29180 41012 29232
rect 43536 29223 43588 29232
rect 43536 29189 43545 29223
rect 43545 29189 43579 29223
rect 43579 29189 43588 29223
rect 43536 29180 43588 29189
rect 42800 29044 42852 29096
rect 39488 28976 39540 29028
rect 44088 29019 44140 29028
rect 44088 28985 44097 29019
rect 44097 28985 44131 29019
rect 44131 28985 44140 29019
rect 49148 29155 49200 29164
rect 49148 29121 49157 29155
rect 49157 29121 49191 29155
rect 49191 29121 49200 29155
rect 49148 29112 49200 29121
rect 51356 29180 51408 29232
rect 44732 29044 44784 29096
rect 46112 29044 46164 29096
rect 48228 29044 48280 29096
rect 44088 28976 44140 28985
rect 49792 28976 49844 29028
rect 13360 28951 13412 28960
rect 13360 28917 13369 28951
rect 13369 28917 13403 28951
rect 13403 28917 13412 28951
rect 13360 28908 13412 28917
rect 38016 28908 38068 28960
rect 40684 28908 40736 28960
rect 42248 28908 42300 28960
rect 45560 28908 45612 28960
rect 47124 28908 47176 28960
rect 51540 29112 51592 29164
rect 51816 29155 51868 29164
rect 51816 29121 51825 29155
rect 51825 29121 51859 29155
rect 51859 29121 51868 29155
rect 51816 29112 51868 29121
rect 52644 29112 52696 29164
rect 53104 29112 53156 29164
rect 53472 29112 53524 29164
rect 53840 29248 53892 29300
rect 55128 29248 55180 29300
rect 55312 29248 55364 29300
rect 55864 29248 55916 29300
rect 56048 29248 56100 29300
rect 56968 29248 57020 29300
rect 57060 29248 57112 29300
rect 58072 29248 58124 29300
rect 52000 29044 52052 29096
rect 54576 29044 54628 29096
rect 52552 29019 52604 29028
rect 52552 28985 52561 29019
rect 52561 28985 52595 29019
rect 52595 28985 52604 29019
rect 55404 29044 55456 29096
rect 56140 29155 56192 29164
rect 56140 29121 56149 29155
rect 56149 29121 56183 29155
rect 56183 29121 56192 29155
rect 56140 29112 56192 29121
rect 56416 29112 56468 29164
rect 57244 29155 57296 29164
rect 57244 29121 57253 29155
rect 57253 29121 57287 29155
rect 57287 29121 57296 29155
rect 57244 29112 57296 29121
rect 57428 29155 57480 29164
rect 57428 29121 57437 29155
rect 57437 29121 57471 29155
rect 57471 29121 57480 29155
rect 57428 29112 57480 29121
rect 52552 28976 52604 28985
rect 56692 28976 56744 29028
rect 53656 28951 53708 28960
rect 53656 28917 53665 28951
rect 53665 28917 53699 28951
rect 53699 28917 53708 28951
rect 53656 28908 53708 28917
rect 55864 28908 55916 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 2044 28704 2096 28756
rect 4068 28704 4120 28756
rect 4712 28704 4764 28756
rect 4896 28704 4948 28756
rect 5816 28704 5868 28756
rect 5908 28747 5960 28756
rect 5908 28713 5917 28747
rect 5917 28713 5951 28747
rect 5951 28713 5960 28747
rect 5908 28704 5960 28713
rect 6092 28704 6144 28756
rect 6736 28704 6788 28756
rect 6828 28704 6880 28756
rect 7288 28704 7340 28756
rect 6552 28679 6604 28688
rect 4804 28568 4856 28620
rect 5448 28568 5500 28620
rect 3608 28500 3660 28552
rect 3700 28500 3752 28552
rect 4068 28500 4120 28552
rect 4160 28543 4212 28552
rect 4160 28509 4169 28543
rect 4169 28509 4203 28543
rect 4203 28509 4212 28543
rect 4160 28500 4212 28509
rect 3792 28432 3844 28484
rect 4620 28500 4672 28552
rect 6552 28645 6561 28679
rect 6561 28645 6595 28679
rect 6595 28645 6604 28679
rect 6552 28636 6604 28645
rect 10508 28704 10560 28756
rect 10600 28747 10652 28756
rect 10600 28713 10609 28747
rect 10609 28713 10643 28747
rect 10643 28713 10652 28747
rect 10600 28704 10652 28713
rect 11244 28747 11296 28756
rect 11244 28713 11253 28747
rect 11253 28713 11287 28747
rect 11287 28713 11296 28747
rect 11244 28704 11296 28713
rect 11888 28704 11940 28756
rect 36268 28704 36320 28756
rect 9864 28636 9916 28688
rect 4896 28432 4948 28484
rect 4988 28432 5040 28484
rect 6920 28500 6972 28552
rect 7196 28500 7248 28552
rect 8392 28432 8444 28484
rect 9956 28500 10008 28552
rect 12532 28568 12584 28620
rect 37464 28704 37516 28756
rect 38384 28704 38436 28756
rect 39028 28704 39080 28756
rect 40684 28704 40736 28756
rect 42800 28747 42852 28756
rect 42800 28713 42809 28747
rect 42809 28713 42843 28747
rect 42843 28713 42852 28747
rect 42800 28704 42852 28713
rect 44640 28704 44692 28756
rect 46112 28704 46164 28756
rect 48136 28704 48188 28756
rect 48320 28704 48372 28756
rect 38016 28636 38068 28688
rect 11060 28500 11112 28552
rect 11336 28543 11388 28552
rect 11336 28509 11345 28543
rect 11345 28509 11379 28543
rect 11379 28509 11388 28543
rect 11336 28500 11388 28509
rect 42248 28611 42300 28620
rect 42248 28577 42257 28611
rect 42257 28577 42291 28611
rect 42291 28577 42300 28611
rect 42248 28568 42300 28577
rect 42800 28568 42852 28620
rect 12992 28500 13044 28552
rect 38568 28543 38620 28552
rect 38568 28509 38577 28543
rect 38577 28509 38611 28543
rect 38611 28509 38620 28543
rect 38568 28500 38620 28509
rect 37464 28432 37516 28484
rect 4712 28364 4764 28416
rect 5356 28364 5408 28416
rect 5540 28364 5592 28416
rect 9128 28364 9180 28416
rect 9312 28364 9364 28416
rect 13360 28364 13412 28416
rect 38660 28432 38712 28484
rect 42524 28500 42576 28552
rect 45192 28636 45244 28688
rect 49148 28704 49200 28756
rect 45652 28611 45704 28620
rect 45652 28577 45661 28611
rect 45661 28577 45695 28611
rect 45695 28577 45704 28611
rect 45652 28568 45704 28577
rect 46572 28568 46624 28620
rect 48320 28568 48372 28620
rect 43260 28475 43312 28484
rect 43260 28441 43269 28475
rect 43269 28441 43303 28475
rect 43303 28441 43312 28475
rect 43260 28432 43312 28441
rect 45192 28543 45244 28552
rect 45192 28509 45201 28543
rect 45201 28509 45235 28543
rect 45235 28509 45244 28543
rect 45192 28500 45244 28509
rect 45560 28500 45612 28552
rect 50160 28704 50212 28756
rect 51540 28747 51592 28756
rect 51540 28713 51549 28747
rect 51549 28713 51583 28747
rect 51583 28713 51592 28747
rect 51540 28704 51592 28713
rect 51816 28704 51868 28756
rect 57152 28747 57204 28756
rect 57152 28713 57161 28747
rect 57161 28713 57195 28747
rect 57195 28713 57204 28747
rect 57152 28704 57204 28713
rect 57428 28704 57480 28756
rect 49884 28636 49936 28688
rect 50252 28568 50304 28620
rect 50620 28543 50672 28552
rect 50620 28509 50629 28543
rect 50629 28509 50663 28543
rect 50663 28509 50672 28543
rect 50620 28500 50672 28509
rect 55220 28636 55272 28688
rect 38476 28407 38528 28416
rect 38476 28373 38485 28407
rect 38485 28373 38519 28407
rect 38519 28373 38528 28407
rect 38476 28364 38528 28373
rect 39304 28364 39356 28416
rect 43076 28364 43128 28416
rect 46572 28432 46624 28484
rect 48044 28432 48096 28484
rect 48228 28364 48280 28416
rect 49148 28364 49200 28416
rect 49700 28475 49752 28484
rect 49700 28441 49709 28475
rect 49709 28441 49743 28475
rect 49743 28441 49752 28475
rect 49700 28432 49752 28441
rect 50712 28432 50764 28484
rect 49976 28364 50028 28416
rect 50068 28364 50120 28416
rect 51724 28500 51776 28552
rect 51540 28364 51592 28416
rect 51724 28364 51776 28416
rect 52000 28500 52052 28552
rect 52184 28500 52236 28552
rect 52552 28500 52604 28552
rect 53656 28500 53708 28552
rect 55864 28500 55916 28552
rect 56416 28500 56468 28552
rect 57612 28543 57664 28552
rect 57612 28509 57621 28543
rect 57621 28509 57655 28543
rect 57655 28509 57664 28543
rect 57612 28500 57664 28509
rect 57704 28543 57756 28552
rect 57704 28509 57713 28543
rect 57713 28509 57747 28543
rect 57747 28509 57756 28543
rect 57704 28500 57756 28509
rect 57796 28500 57848 28552
rect 58348 28543 58400 28552
rect 58348 28509 58357 28543
rect 58357 28509 58391 28543
rect 58391 28509 58400 28543
rect 58348 28500 58400 28509
rect 53196 28364 53248 28416
rect 53288 28407 53340 28416
rect 53288 28373 53297 28407
rect 53297 28373 53331 28407
rect 53331 28373 53340 28407
rect 53288 28364 53340 28373
rect 56600 28364 56652 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 3976 28203 4028 28212
rect 3976 28169 3985 28203
rect 3985 28169 4019 28203
rect 4019 28169 4028 28203
rect 3976 28160 4028 28169
rect 4068 28160 4120 28212
rect 6368 28160 6420 28212
rect 7104 28160 7156 28212
rect 2688 28067 2740 28076
rect 2688 28033 2697 28067
rect 2697 28033 2731 28067
rect 2731 28033 2740 28067
rect 2688 28024 2740 28033
rect 1584 27999 1636 28008
rect 1584 27965 1593 27999
rect 1593 27965 1627 27999
rect 1627 27965 1636 27999
rect 1584 27956 1636 27965
rect 3424 27999 3476 28008
rect 3424 27965 3433 27999
rect 3433 27965 3467 27999
rect 3467 27965 3476 27999
rect 3424 27956 3476 27965
rect 4804 28024 4856 28076
rect 8392 28092 8444 28144
rect 8760 28160 8812 28212
rect 9128 28203 9180 28212
rect 9128 28169 9137 28203
rect 9137 28169 9171 28203
rect 9171 28169 9180 28203
rect 9128 28160 9180 28169
rect 10232 28203 10284 28212
rect 10232 28169 10241 28203
rect 10241 28169 10275 28203
rect 10275 28169 10284 28203
rect 10232 28160 10284 28169
rect 38476 28160 38528 28212
rect 38568 28160 38620 28212
rect 39212 28160 39264 28212
rect 40040 28160 40092 28212
rect 8484 28067 8536 28076
rect 8484 28033 8493 28067
rect 8493 28033 8527 28067
rect 8527 28033 8536 28067
rect 8484 28024 8536 28033
rect 11336 28092 11388 28144
rect 9864 28024 9916 28076
rect 13084 28024 13136 28076
rect 4988 27956 5040 28008
rect 8668 27999 8720 28008
rect 4160 27888 4212 27940
rect 8668 27965 8677 27999
rect 8677 27965 8711 27999
rect 8711 27965 8720 27999
rect 8668 27956 8720 27965
rect 8944 27956 8996 28008
rect 10140 27956 10192 28008
rect 11060 27956 11112 28008
rect 12900 27999 12952 28008
rect 12900 27965 12909 27999
rect 12909 27965 12943 27999
rect 12943 27965 12952 27999
rect 12900 27956 12952 27965
rect 38108 28067 38160 28076
rect 38108 28033 38117 28067
rect 38117 28033 38151 28067
rect 38151 28033 38160 28067
rect 38108 28024 38160 28033
rect 43260 28160 43312 28212
rect 43628 28203 43680 28212
rect 40040 28067 40092 28076
rect 40040 28033 40049 28067
rect 40049 28033 40083 28067
rect 40083 28033 40092 28067
rect 40040 28024 40092 28033
rect 43628 28169 43637 28203
rect 43637 28169 43671 28203
rect 43671 28169 43680 28203
rect 43628 28160 43680 28169
rect 44640 28160 44692 28212
rect 45192 28160 45244 28212
rect 49056 28160 49108 28212
rect 49700 28203 49752 28212
rect 49700 28169 49709 28203
rect 49709 28169 49743 28203
rect 49743 28169 49752 28203
rect 49700 28160 49752 28169
rect 50160 28160 50212 28212
rect 53840 28160 53892 28212
rect 57704 28160 57756 28212
rect 58808 28160 58860 28212
rect 39672 27999 39724 28008
rect 39672 27965 39681 27999
rect 39681 27965 39715 27999
rect 39715 27965 39724 27999
rect 39672 27956 39724 27965
rect 40224 28024 40276 28076
rect 40408 28067 40460 28076
rect 40408 28033 40417 28067
rect 40417 28033 40451 28067
rect 40451 28033 40460 28067
rect 40408 28024 40460 28033
rect 40684 28024 40736 28076
rect 41328 28067 41380 28076
rect 41328 28033 41337 28067
rect 41337 28033 41371 28067
rect 41371 28033 41380 28067
rect 41328 28024 41380 28033
rect 41972 28067 42024 28076
rect 41972 28033 41981 28067
rect 41981 28033 42015 28067
rect 42015 28033 42024 28067
rect 41972 28024 42024 28033
rect 40316 27956 40368 28008
rect 2780 27820 2832 27872
rect 4620 27820 4672 27872
rect 5356 27863 5408 27872
rect 5356 27829 5365 27863
rect 5365 27829 5399 27863
rect 5399 27829 5408 27863
rect 5356 27820 5408 27829
rect 6092 27820 6144 27872
rect 7656 27820 7708 27872
rect 10324 27820 10376 27872
rect 11244 27820 11296 27872
rect 37924 27820 37976 27872
rect 40224 27820 40276 27872
rect 40408 27820 40460 27872
rect 43444 28067 43496 28076
rect 43444 28033 43453 28067
rect 43453 28033 43487 28067
rect 43487 28033 43496 28067
rect 43444 28024 43496 28033
rect 46388 28092 46440 28144
rect 47124 28092 47176 28144
rect 43628 27956 43680 28008
rect 47216 28067 47268 28076
rect 47216 28033 47225 28067
rect 47225 28033 47259 28067
rect 47259 28033 47268 28067
rect 47216 28024 47268 28033
rect 44640 27999 44692 28008
rect 44640 27965 44649 27999
rect 44649 27965 44683 27999
rect 44683 27965 44692 27999
rect 44640 27956 44692 27965
rect 47124 27999 47176 28008
rect 47124 27965 47133 27999
rect 47133 27965 47167 27999
rect 47167 27965 47176 27999
rect 47124 27956 47176 27965
rect 47584 28024 47636 28076
rect 47860 28067 47912 28076
rect 47860 28033 47869 28067
rect 47869 28033 47903 28067
rect 47903 28033 47912 28067
rect 47860 28024 47912 28033
rect 49240 28024 49292 28076
rect 51908 28092 51960 28144
rect 50160 28067 50212 28076
rect 47768 27888 47820 27940
rect 47952 27888 48004 27940
rect 48228 27956 48280 28008
rect 49424 27956 49476 28008
rect 50160 28033 50169 28067
rect 50169 28033 50203 28067
rect 50203 28033 50212 28067
rect 50160 28024 50212 28033
rect 51172 28024 51224 28076
rect 52368 28067 52420 28076
rect 52368 28033 52377 28067
rect 52377 28033 52411 28067
rect 52411 28033 52420 28067
rect 52368 28024 52420 28033
rect 52552 28067 52604 28076
rect 52552 28033 52561 28067
rect 52561 28033 52595 28067
rect 52595 28033 52604 28067
rect 52552 28024 52604 28033
rect 54024 28024 54076 28076
rect 56508 28092 56560 28144
rect 56784 28092 56836 28144
rect 56416 28067 56468 28076
rect 56416 28033 56450 28067
rect 56450 28033 56468 28067
rect 52920 27956 52972 28008
rect 55680 27999 55732 28008
rect 55680 27965 55689 27999
rect 55689 27965 55723 27999
rect 55723 27965 55732 27999
rect 55680 27956 55732 27965
rect 56416 28024 56468 28033
rect 48136 27820 48188 27872
rect 48228 27820 48280 27872
rect 49976 27820 50028 27872
rect 51632 27863 51684 27872
rect 51632 27829 51641 27863
rect 51641 27829 51675 27863
rect 51675 27829 51684 27863
rect 51632 27820 51684 27829
rect 55036 27820 55088 27872
rect 55864 27863 55916 27872
rect 55864 27829 55873 27863
rect 55873 27829 55907 27863
rect 55907 27829 55916 27863
rect 55864 27820 55916 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3424 27616 3476 27668
rect 3240 27548 3292 27600
rect 3240 27455 3292 27464
rect 3240 27421 3249 27455
rect 3249 27421 3283 27455
rect 3283 27421 3292 27455
rect 3240 27412 3292 27421
rect 3424 27455 3476 27464
rect 3424 27421 3433 27455
rect 3433 27421 3467 27455
rect 3467 27421 3476 27455
rect 3424 27412 3476 27421
rect 4620 27616 4672 27668
rect 10968 27659 11020 27668
rect 10968 27625 10977 27659
rect 10977 27625 11011 27659
rect 11011 27625 11020 27659
rect 10968 27616 11020 27625
rect 11336 27616 11388 27668
rect 6828 27480 6880 27532
rect 8392 27480 8444 27532
rect 8852 27480 8904 27532
rect 10416 27480 10468 27532
rect 5632 27412 5684 27464
rect 6460 27455 6512 27464
rect 6460 27421 6469 27455
rect 6469 27421 6503 27455
rect 6503 27421 6512 27455
rect 6460 27412 6512 27421
rect 6552 27412 6604 27464
rect 7472 27455 7524 27464
rect 7472 27421 7481 27455
rect 7481 27421 7515 27455
rect 7515 27421 7524 27455
rect 7472 27412 7524 27421
rect 10232 27412 10284 27464
rect 12348 27455 12400 27464
rect 12348 27421 12357 27455
rect 12357 27421 12391 27455
rect 12391 27421 12400 27455
rect 12348 27412 12400 27421
rect 2412 27344 2464 27396
rect 2872 27387 2924 27396
rect 2872 27353 2881 27387
rect 2881 27353 2915 27387
rect 2915 27353 2924 27387
rect 2872 27344 2924 27353
rect 4160 27344 4212 27396
rect 5264 27344 5316 27396
rect 7656 27387 7708 27396
rect 7656 27353 7665 27387
rect 7665 27353 7699 27387
rect 7699 27353 7708 27387
rect 7656 27344 7708 27353
rect 2688 27276 2740 27328
rect 4804 27276 4856 27328
rect 5172 27276 5224 27328
rect 6276 27319 6328 27328
rect 6276 27285 6285 27319
rect 6285 27285 6319 27319
rect 6319 27285 6328 27319
rect 6276 27276 6328 27285
rect 6736 27276 6788 27328
rect 11244 27344 11296 27396
rect 11336 27344 11388 27396
rect 8208 27276 8260 27328
rect 11980 27276 12032 27328
rect 12624 27455 12676 27464
rect 12624 27421 12633 27455
rect 12633 27421 12667 27455
rect 12667 27421 12676 27455
rect 12624 27412 12676 27421
rect 12808 27455 12860 27464
rect 12808 27421 12817 27455
rect 12817 27421 12851 27455
rect 12851 27421 12860 27455
rect 12808 27412 12860 27421
rect 12900 27412 12952 27464
rect 13176 27455 13228 27464
rect 13176 27421 13185 27455
rect 13185 27421 13219 27455
rect 13219 27421 13228 27455
rect 13176 27412 13228 27421
rect 39672 27616 39724 27668
rect 40040 27616 40092 27668
rect 40316 27616 40368 27668
rect 42984 27616 43036 27668
rect 43444 27616 43496 27668
rect 43720 27616 43772 27668
rect 13360 27276 13412 27328
rect 25320 27387 25372 27396
rect 25320 27353 25329 27387
rect 25329 27353 25363 27387
rect 25363 27353 25372 27387
rect 25320 27344 25372 27353
rect 37924 27455 37976 27464
rect 37924 27421 37933 27455
rect 37933 27421 37967 27455
rect 37967 27421 37976 27455
rect 37924 27412 37976 27421
rect 38016 27455 38068 27464
rect 38016 27421 38025 27455
rect 38025 27421 38059 27455
rect 38059 27421 38068 27455
rect 38016 27412 38068 27421
rect 38476 27412 38528 27464
rect 38660 27455 38712 27464
rect 38660 27421 38669 27455
rect 38669 27421 38703 27455
rect 38703 27421 38712 27455
rect 38660 27412 38712 27421
rect 39212 27480 39264 27532
rect 40500 27480 40552 27532
rect 39396 27412 39448 27464
rect 39856 27412 39908 27464
rect 40224 27412 40276 27464
rect 40684 27412 40736 27464
rect 43904 27480 43956 27532
rect 46388 27616 46440 27668
rect 47952 27616 48004 27668
rect 52920 27616 52972 27668
rect 53196 27659 53248 27668
rect 53196 27625 53205 27659
rect 53205 27625 53239 27659
rect 53239 27625 53248 27659
rect 53196 27616 53248 27625
rect 54024 27616 54076 27668
rect 55680 27616 55732 27668
rect 56416 27659 56468 27668
rect 56416 27625 56425 27659
rect 56425 27625 56459 27659
rect 56459 27625 56468 27659
rect 56416 27616 56468 27625
rect 58348 27659 58400 27668
rect 58348 27625 58357 27659
rect 58357 27625 58391 27659
rect 58391 27625 58400 27659
rect 58348 27616 58400 27625
rect 44916 27548 44968 27600
rect 45836 27548 45888 27600
rect 46020 27548 46072 27600
rect 50620 27591 50672 27600
rect 38660 27276 38712 27328
rect 39212 27319 39264 27328
rect 39212 27285 39221 27319
rect 39221 27285 39255 27319
rect 39255 27285 39264 27319
rect 39212 27276 39264 27285
rect 39304 27276 39356 27328
rect 42156 27319 42208 27328
rect 42156 27285 42165 27319
rect 42165 27285 42199 27319
rect 42199 27285 42208 27319
rect 42156 27276 42208 27285
rect 42892 27319 42944 27328
rect 42892 27285 42901 27319
rect 42901 27285 42935 27319
rect 42935 27285 42944 27319
rect 42892 27276 42944 27285
rect 43536 27276 43588 27328
rect 44824 27412 44876 27464
rect 45652 27412 45704 27464
rect 45928 27455 45980 27464
rect 45928 27421 45937 27455
rect 45937 27421 45971 27455
rect 45971 27421 45980 27455
rect 45928 27412 45980 27421
rect 46480 27455 46532 27464
rect 45284 27344 45336 27396
rect 44732 27319 44784 27328
rect 44732 27285 44741 27319
rect 44741 27285 44775 27319
rect 44775 27285 44784 27319
rect 44732 27276 44784 27285
rect 45744 27276 45796 27328
rect 46480 27421 46489 27455
rect 46489 27421 46523 27455
rect 46523 27421 46532 27455
rect 46480 27412 46532 27421
rect 47768 27412 47820 27464
rect 48136 27412 48188 27464
rect 48320 27455 48372 27464
rect 48320 27421 48329 27455
rect 48329 27421 48363 27455
rect 48363 27421 48372 27455
rect 48320 27412 48372 27421
rect 48596 27412 48648 27464
rect 49056 27412 49108 27464
rect 50620 27557 50629 27591
rect 50629 27557 50663 27591
rect 50663 27557 50672 27591
rect 50620 27548 50672 27557
rect 56784 27548 56836 27600
rect 56140 27480 56192 27532
rect 49700 27344 49752 27396
rect 49976 27412 50028 27464
rect 50988 27455 51040 27464
rect 50988 27421 50997 27455
rect 50997 27421 51031 27455
rect 51031 27421 51040 27455
rect 50988 27412 51040 27421
rect 51908 27412 51960 27464
rect 51448 27387 51500 27396
rect 51448 27353 51482 27387
rect 51482 27353 51500 27387
rect 51448 27344 51500 27353
rect 53840 27412 53892 27464
rect 48688 27319 48740 27328
rect 48688 27285 48697 27319
rect 48697 27285 48731 27319
rect 48731 27285 48740 27319
rect 48688 27276 48740 27285
rect 48780 27276 48832 27328
rect 49240 27276 49292 27328
rect 50896 27276 50948 27328
rect 53012 27276 53064 27328
rect 53840 27276 53892 27328
rect 54852 27455 54904 27464
rect 54852 27421 54861 27455
rect 54861 27421 54895 27455
rect 54895 27421 54904 27455
rect 54852 27412 54904 27421
rect 55036 27455 55088 27464
rect 55036 27421 55045 27455
rect 55045 27421 55079 27455
rect 55079 27421 55088 27455
rect 55036 27412 55088 27421
rect 55864 27412 55916 27464
rect 56416 27412 56468 27464
rect 56600 27455 56652 27464
rect 56600 27421 56609 27455
rect 56609 27421 56643 27455
rect 56643 27421 56652 27455
rect 56600 27412 56652 27421
rect 56876 27480 56928 27532
rect 54944 27276 54996 27328
rect 56140 27276 56192 27328
rect 56324 27276 56376 27328
rect 57704 27412 57756 27464
rect 58900 27412 58952 27464
rect 58716 27344 58768 27396
rect 58164 27319 58216 27328
rect 58164 27285 58173 27319
rect 58173 27285 58207 27319
rect 58207 27285 58216 27319
rect 58164 27276 58216 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 2872 27072 2924 27124
rect 3424 27072 3476 27124
rect 4160 27072 4212 27124
rect 4712 27072 4764 27124
rect 2780 26911 2832 26920
rect 2780 26877 2789 26911
rect 2789 26877 2823 26911
rect 2823 26877 2832 26911
rect 2780 26868 2832 26877
rect 2688 26800 2740 26852
rect 3792 26800 3844 26852
rect 4988 26979 5040 26988
rect 4988 26945 4997 26979
rect 4997 26945 5031 26979
rect 5031 26945 5040 26979
rect 4988 26936 5040 26945
rect 5172 27004 5224 27056
rect 6276 27004 6328 27056
rect 6368 27004 6420 27056
rect 5632 26936 5684 26988
rect 6092 26936 6144 26988
rect 4620 26868 4672 26920
rect 7196 26979 7248 26988
rect 7196 26945 7205 26979
rect 7205 26945 7239 26979
rect 7239 26945 7248 26979
rect 7196 26936 7248 26945
rect 7472 27004 7524 27056
rect 9956 27072 10008 27124
rect 11336 27115 11388 27124
rect 11336 27081 11345 27115
rect 11345 27081 11379 27115
rect 11379 27081 11388 27115
rect 11336 27072 11388 27081
rect 12808 27115 12860 27124
rect 12808 27081 12817 27115
rect 12817 27081 12851 27115
rect 12851 27081 12860 27115
rect 12808 27072 12860 27081
rect 38016 27072 38068 27124
rect 38568 27072 38620 27124
rect 42892 27072 42944 27124
rect 42984 27072 43036 27124
rect 43076 27115 43128 27124
rect 43076 27081 43085 27115
rect 43085 27081 43119 27115
rect 43119 27081 43128 27115
rect 43076 27072 43128 27081
rect 7840 26979 7892 26988
rect 7840 26945 7874 26979
rect 7874 26945 7892 26979
rect 7840 26936 7892 26945
rect 8208 26936 8260 26988
rect 9772 26936 9824 26988
rect 10416 26979 10468 26988
rect 10416 26945 10425 26979
rect 10425 26945 10459 26979
rect 10459 26945 10468 26979
rect 10416 26936 10468 26945
rect 11520 26936 11572 26988
rect 11704 26936 11756 26988
rect 5080 26800 5132 26852
rect 3332 26732 3384 26784
rect 5816 26775 5868 26784
rect 5816 26741 5825 26775
rect 5825 26741 5859 26775
rect 5859 26741 5868 26775
rect 5816 26732 5868 26741
rect 6184 26732 6236 26784
rect 6552 26775 6604 26784
rect 6552 26741 6561 26775
rect 6561 26741 6595 26775
rect 6595 26741 6604 26775
rect 6552 26732 6604 26741
rect 7104 26775 7156 26784
rect 7104 26741 7113 26775
rect 7113 26741 7147 26775
rect 7147 26741 7156 26775
rect 7104 26732 7156 26741
rect 25320 27004 25372 27056
rect 38108 27004 38160 27056
rect 39396 27004 39448 27056
rect 42156 27004 42208 27056
rect 43352 27047 43404 27056
rect 38752 26936 38804 26988
rect 38844 26979 38896 26988
rect 38844 26945 38853 26979
rect 38853 26945 38887 26979
rect 38887 26945 38896 26979
rect 38844 26936 38896 26945
rect 39856 26979 39908 26988
rect 37280 26868 37332 26920
rect 38660 26800 38712 26852
rect 39856 26945 39865 26979
rect 39865 26945 39899 26979
rect 39899 26945 39908 26979
rect 39856 26936 39908 26945
rect 39948 26979 40000 26988
rect 39948 26945 39957 26979
rect 39957 26945 39991 26979
rect 39991 26945 40000 26979
rect 39948 26936 40000 26945
rect 40132 26936 40184 26988
rect 42432 26979 42484 26988
rect 40224 26911 40276 26920
rect 40224 26877 40233 26911
rect 40233 26877 40267 26911
rect 40267 26877 40276 26911
rect 40224 26868 40276 26877
rect 9956 26775 10008 26784
rect 9956 26741 9965 26775
rect 9965 26741 9999 26775
rect 9999 26741 10008 26775
rect 9956 26732 10008 26741
rect 10508 26732 10560 26784
rect 10600 26732 10652 26784
rect 11704 26775 11756 26784
rect 11704 26741 11713 26775
rect 11713 26741 11747 26775
rect 11747 26741 11756 26775
rect 11704 26732 11756 26741
rect 13360 26732 13412 26784
rect 36268 26775 36320 26784
rect 36268 26741 36277 26775
rect 36277 26741 36311 26775
rect 36311 26741 36320 26775
rect 36268 26732 36320 26741
rect 36728 26732 36780 26784
rect 37464 26775 37516 26784
rect 37464 26741 37473 26775
rect 37473 26741 37507 26775
rect 37507 26741 37516 26775
rect 37464 26732 37516 26741
rect 39120 26732 39172 26784
rect 40684 26732 40736 26784
rect 42432 26945 42441 26979
rect 42441 26945 42475 26979
rect 42475 26945 42484 26979
rect 42432 26936 42484 26945
rect 42616 26979 42668 26988
rect 42616 26945 42625 26979
rect 42625 26945 42659 26979
rect 42659 26945 42668 26979
rect 42616 26936 42668 26945
rect 43352 27013 43361 27047
rect 43361 27013 43395 27047
rect 43395 27013 43404 27047
rect 43352 27004 43404 27013
rect 46112 27072 46164 27124
rect 46480 27072 46532 27124
rect 43536 27047 43588 27056
rect 43536 27013 43571 27047
rect 43571 27013 43588 27047
rect 43536 27004 43588 27013
rect 43720 27004 43772 27056
rect 43996 27004 44048 27056
rect 44916 27047 44968 27056
rect 44916 27013 44925 27047
rect 44925 27013 44959 27047
rect 44959 27013 44968 27047
rect 44916 27004 44968 27013
rect 45928 27004 45980 27056
rect 43260 26979 43312 26988
rect 43260 26945 43269 26979
rect 43269 26945 43303 26979
rect 43303 26945 43312 26979
rect 43260 26936 43312 26945
rect 43904 26936 43956 26988
rect 45744 26979 45796 26988
rect 45744 26945 45753 26979
rect 45753 26945 45787 26979
rect 45787 26945 45796 26979
rect 45744 26936 45796 26945
rect 46020 26936 46072 26988
rect 47216 27004 47268 27056
rect 51448 27115 51500 27124
rect 51448 27081 51457 27115
rect 51457 27081 51491 27115
rect 51491 27081 51500 27115
rect 51448 27072 51500 27081
rect 51540 27072 51592 27124
rect 49976 27004 50028 27056
rect 46572 26979 46624 26988
rect 46572 26945 46581 26979
rect 46581 26945 46615 26979
rect 46615 26945 46624 26979
rect 46572 26936 46624 26945
rect 47676 26936 47728 26988
rect 48228 26979 48280 26988
rect 48228 26945 48237 26979
rect 48237 26945 48271 26979
rect 48271 26945 48280 26979
rect 48228 26936 48280 26945
rect 48780 26936 48832 26988
rect 49700 26936 49752 26988
rect 50896 26979 50948 26988
rect 50896 26945 50905 26979
rect 50905 26945 50939 26979
rect 50939 26945 50948 26979
rect 50896 26936 50948 26945
rect 54116 27072 54168 27124
rect 54576 27115 54628 27124
rect 54576 27081 54585 27115
rect 54585 27081 54619 27115
rect 54619 27081 54628 27115
rect 54576 27072 54628 27081
rect 58164 27072 58216 27124
rect 52184 27004 52236 27056
rect 42340 26732 42392 26784
rect 45836 26800 45888 26852
rect 46020 26800 46072 26852
rect 47308 26800 47360 26852
rect 50160 26911 50212 26920
rect 50160 26877 50169 26911
rect 50169 26877 50203 26911
rect 50203 26877 50212 26911
rect 50160 26868 50212 26877
rect 51632 26868 51684 26920
rect 53932 26936 53984 26988
rect 54852 26936 54904 26988
rect 57152 26936 57204 26988
rect 54484 26868 54536 26920
rect 56048 26911 56100 26920
rect 56048 26877 56057 26911
rect 56057 26877 56091 26911
rect 56091 26877 56100 26911
rect 56048 26868 56100 26877
rect 56324 26868 56376 26920
rect 47584 26732 47636 26784
rect 51724 26800 51776 26852
rect 48504 26732 48556 26784
rect 48780 26775 48832 26784
rect 48780 26741 48789 26775
rect 48789 26741 48823 26775
rect 48823 26741 48832 26775
rect 48780 26732 48832 26741
rect 50804 26775 50856 26784
rect 50804 26741 50813 26775
rect 50813 26741 50847 26775
rect 50847 26741 50856 26775
rect 50804 26732 50856 26741
rect 51632 26775 51684 26784
rect 51632 26741 51641 26775
rect 51641 26741 51675 26775
rect 51675 26741 51684 26775
rect 53656 26800 53708 26852
rect 51632 26732 51684 26741
rect 53380 26732 53432 26784
rect 55404 26775 55456 26784
rect 55404 26741 55413 26775
rect 55413 26741 55447 26775
rect 55447 26741 55456 26775
rect 55404 26732 55456 26741
rect 56968 26775 57020 26784
rect 56968 26741 56977 26775
rect 56977 26741 57011 26775
rect 57011 26741 57020 26775
rect 56968 26732 57020 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 5724 26528 5776 26580
rect 6552 26528 6604 26580
rect 7840 26528 7892 26580
rect 9680 26528 9732 26580
rect 10140 26528 10192 26580
rect 6092 26460 6144 26512
rect 9220 26460 9272 26512
rect 10600 26460 10652 26512
rect 3240 26392 3292 26444
rect 7104 26392 7156 26444
rect 7472 26392 7524 26444
rect 8392 26392 8444 26444
rect 1400 26324 1452 26376
rect 3976 26367 4028 26376
rect 3976 26333 3985 26367
rect 3985 26333 4019 26367
rect 4019 26333 4028 26367
rect 3976 26324 4028 26333
rect 4620 26367 4672 26376
rect 4620 26333 4629 26367
rect 4629 26333 4663 26367
rect 4663 26333 4672 26367
rect 4620 26324 4672 26333
rect 5172 26324 5224 26376
rect 1584 26299 1636 26308
rect 1584 26265 1593 26299
rect 1593 26265 1627 26299
rect 1627 26265 1636 26299
rect 1584 26256 1636 26265
rect 5448 26256 5500 26308
rect 7564 26256 7616 26308
rect 10968 26324 11020 26376
rect 11336 26324 11388 26376
rect 40224 26528 40276 26580
rect 40592 26528 40644 26580
rect 42432 26528 42484 26580
rect 42800 26528 42852 26580
rect 46388 26528 46440 26580
rect 47860 26571 47912 26580
rect 47860 26537 47869 26571
rect 47869 26537 47903 26571
rect 47903 26537 47912 26571
rect 47860 26528 47912 26537
rect 48504 26571 48556 26580
rect 48504 26537 48534 26571
rect 48534 26537 48556 26571
rect 48504 26528 48556 26537
rect 50160 26528 50212 26580
rect 39120 26503 39172 26512
rect 39120 26469 39129 26503
rect 39129 26469 39163 26503
rect 39163 26469 39172 26503
rect 39120 26460 39172 26469
rect 39212 26460 39264 26512
rect 39948 26460 40000 26512
rect 35440 26435 35492 26444
rect 35440 26401 35449 26435
rect 35449 26401 35483 26435
rect 35483 26401 35492 26435
rect 35440 26392 35492 26401
rect 10876 26256 10928 26308
rect 11612 26256 11664 26308
rect 12624 26256 12676 26308
rect 37832 26324 37884 26376
rect 38108 26324 38160 26376
rect 40316 26392 40368 26444
rect 41696 26460 41748 26512
rect 42340 26392 42392 26444
rect 39212 26324 39264 26376
rect 40408 26367 40460 26376
rect 40408 26333 40417 26367
rect 40417 26333 40451 26367
rect 40451 26333 40460 26367
rect 40408 26324 40460 26333
rect 51908 26528 51960 26580
rect 53748 26571 53800 26580
rect 53748 26537 53757 26571
rect 53757 26537 53791 26571
rect 53791 26537 53800 26571
rect 53748 26528 53800 26537
rect 53840 26528 53892 26580
rect 54484 26528 54536 26580
rect 54760 26528 54812 26580
rect 54944 26571 54996 26580
rect 54944 26537 54953 26571
rect 54953 26537 54987 26571
rect 54987 26537 54996 26571
rect 54944 26528 54996 26537
rect 56048 26528 56100 26580
rect 44824 26503 44876 26512
rect 44824 26469 44833 26503
rect 44833 26469 44867 26503
rect 44867 26469 44876 26503
rect 44824 26460 44876 26469
rect 43904 26324 43956 26376
rect 43996 26324 44048 26376
rect 44456 26324 44508 26376
rect 45192 26367 45244 26376
rect 45192 26333 45201 26367
rect 45201 26333 45235 26367
rect 45235 26333 45244 26367
rect 45192 26324 45244 26333
rect 45376 26314 45428 26366
rect 45652 26392 45704 26444
rect 51080 26460 51132 26512
rect 47124 26392 47176 26444
rect 48504 26392 48556 26444
rect 53472 26392 53524 26444
rect 35716 26299 35768 26308
rect 35716 26265 35725 26299
rect 35725 26265 35759 26299
rect 35759 26265 35768 26299
rect 35716 26256 35768 26265
rect 36728 26256 36780 26308
rect 3884 26231 3936 26240
rect 3884 26197 3893 26231
rect 3893 26197 3927 26231
rect 3927 26197 3936 26231
rect 3884 26188 3936 26197
rect 4804 26231 4856 26240
rect 4804 26197 4813 26231
rect 4813 26197 4847 26231
rect 4847 26197 4856 26231
rect 4804 26188 4856 26197
rect 7748 26231 7800 26240
rect 7748 26197 7757 26231
rect 7757 26197 7791 26231
rect 7791 26197 7800 26231
rect 7748 26188 7800 26197
rect 10140 26188 10192 26240
rect 10324 26188 10376 26240
rect 12348 26188 12400 26240
rect 13360 26188 13412 26240
rect 37096 26188 37148 26240
rect 38752 26256 38804 26308
rect 39120 26299 39172 26308
rect 39120 26265 39129 26299
rect 39129 26265 39163 26299
rect 39163 26265 39172 26299
rect 39120 26256 39172 26265
rect 37924 26231 37976 26240
rect 37924 26197 37933 26231
rect 37933 26197 37967 26231
rect 37967 26197 37976 26231
rect 37924 26188 37976 26197
rect 38844 26188 38896 26240
rect 40776 26188 40828 26240
rect 42156 26188 42208 26240
rect 43352 26188 43404 26240
rect 45744 26188 45796 26240
rect 46388 26367 46440 26376
rect 46388 26333 46397 26367
rect 46397 26333 46431 26367
rect 46431 26333 46440 26367
rect 46388 26324 46440 26333
rect 46940 26324 46992 26376
rect 47308 26324 47360 26376
rect 48044 26324 48096 26376
rect 51816 26324 51868 26376
rect 52736 26367 52788 26376
rect 52736 26333 52745 26367
rect 52745 26333 52779 26367
rect 52779 26333 52788 26367
rect 52736 26324 52788 26333
rect 46480 26299 46532 26308
rect 46480 26265 46489 26299
rect 46489 26265 46523 26299
rect 46523 26265 46532 26299
rect 46480 26256 46532 26265
rect 46848 26188 46900 26240
rect 48412 26256 48464 26308
rect 49792 26256 49844 26308
rect 52828 26256 52880 26308
rect 53656 26460 53708 26512
rect 55312 26460 55364 26512
rect 56508 26392 56560 26444
rect 53748 26367 53800 26376
rect 53748 26333 53757 26367
rect 53757 26333 53791 26367
rect 53791 26333 53800 26367
rect 53748 26324 53800 26333
rect 53840 26367 53892 26376
rect 53840 26333 53849 26367
rect 53849 26333 53883 26367
rect 53883 26333 53892 26367
rect 53840 26324 53892 26333
rect 54484 26367 54536 26376
rect 54484 26333 54493 26367
rect 54493 26333 54527 26367
rect 54527 26333 54536 26367
rect 54484 26324 54536 26333
rect 54576 26324 54628 26376
rect 54208 26299 54260 26308
rect 54208 26265 54217 26299
rect 54217 26265 54251 26299
rect 54251 26265 54260 26299
rect 54208 26256 54260 26265
rect 47676 26231 47728 26240
rect 47676 26197 47685 26231
rect 47685 26197 47719 26231
rect 47719 26197 47728 26231
rect 47676 26188 47728 26197
rect 53748 26188 53800 26240
rect 54116 26188 54168 26240
rect 54300 26231 54352 26240
rect 54300 26197 54309 26231
rect 54309 26197 54343 26231
rect 54343 26197 54352 26231
rect 54300 26188 54352 26197
rect 55220 26324 55272 26376
rect 58900 26324 58952 26376
rect 57060 26299 57112 26308
rect 57060 26265 57094 26299
rect 57094 26265 57112 26299
rect 57060 26256 57112 26265
rect 54852 26188 54904 26240
rect 55036 26188 55088 26240
rect 58256 26231 58308 26240
rect 58256 26197 58265 26231
rect 58265 26197 58299 26231
rect 58299 26197 58308 26231
rect 58256 26188 58308 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 1400 26027 1452 26036
rect 1400 25993 1409 26027
rect 1409 25993 1443 26027
rect 1443 25993 1452 26027
rect 1400 25984 1452 25993
rect 5448 26027 5500 26036
rect 5448 25993 5457 26027
rect 5457 25993 5491 26027
rect 5491 25993 5500 26027
rect 5448 25984 5500 25993
rect 7748 25984 7800 26036
rect 2412 25916 2464 25968
rect 9680 25984 9732 26036
rect 3884 25891 3936 25900
rect 3884 25857 3893 25891
rect 3893 25857 3927 25891
rect 3927 25857 3936 25891
rect 3884 25848 3936 25857
rect 4620 25848 4672 25900
rect 3148 25823 3200 25832
rect 3148 25789 3157 25823
rect 3157 25789 3191 25823
rect 3191 25789 3200 25823
rect 3148 25780 3200 25789
rect 4068 25823 4120 25832
rect 4068 25789 4077 25823
rect 4077 25789 4111 25823
rect 4111 25789 4120 25823
rect 4068 25780 4120 25789
rect 3424 25712 3476 25764
rect 7840 25848 7892 25900
rect 8484 25891 8536 25900
rect 8484 25857 8493 25891
rect 8493 25857 8527 25891
rect 8527 25857 8536 25891
rect 8484 25848 8536 25857
rect 8576 25891 8628 25900
rect 8576 25857 8585 25891
rect 8585 25857 8619 25891
rect 8619 25857 8628 25891
rect 8576 25848 8628 25857
rect 8668 25848 8720 25900
rect 9036 25848 9088 25900
rect 3240 25687 3292 25696
rect 3240 25653 3249 25687
rect 3249 25653 3283 25687
rect 3283 25653 3292 25687
rect 3240 25644 3292 25653
rect 7196 25687 7248 25696
rect 7196 25653 7205 25687
rect 7205 25653 7239 25687
rect 7239 25653 7248 25687
rect 7196 25644 7248 25653
rect 7472 25644 7524 25696
rect 8760 25687 8812 25696
rect 8760 25653 8769 25687
rect 8769 25653 8803 25687
rect 8803 25653 8812 25687
rect 8760 25644 8812 25653
rect 9128 25687 9180 25696
rect 9128 25653 9137 25687
rect 9137 25653 9171 25687
rect 9171 25653 9180 25687
rect 9128 25644 9180 25653
rect 9772 25916 9824 25968
rect 10416 25984 10468 26036
rect 10876 25984 10928 26036
rect 10968 25984 11020 26036
rect 11520 26027 11572 26036
rect 11520 25993 11529 26027
rect 11529 25993 11563 26027
rect 11563 25993 11572 26027
rect 11520 25984 11572 25993
rect 11888 25984 11940 26036
rect 10416 25848 10468 25900
rect 11612 25916 11664 25968
rect 12624 25984 12676 26036
rect 35716 26027 35768 26036
rect 35716 25993 35725 26027
rect 35725 25993 35759 26027
rect 35759 25993 35768 26027
rect 35716 25984 35768 25993
rect 36268 25984 36320 26036
rect 11152 25891 11204 25900
rect 11152 25857 11161 25891
rect 11161 25857 11195 25891
rect 11195 25857 11204 25891
rect 11152 25848 11204 25857
rect 11336 25891 11388 25900
rect 11336 25857 11345 25891
rect 11345 25857 11379 25891
rect 11379 25857 11388 25891
rect 11336 25848 11388 25857
rect 12072 25848 12124 25900
rect 14924 25848 14976 25900
rect 37096 25984 37148 26036
rect 37280 26027 37332 26036
rect 37280 25993 37289 26027
rect 37289 25993 37323 26027
rect 37323 25993 37332 26027
rect 37280 25984 37332 25993
rect 37832 26027 37884 26036
rect 37832 25993 37841 26027
rect 37841 25993 37875 26027
rect 37875 25993 37884 26027
rect 37832 25984 37884 25993
rect 37924 25984 37976 26036
rect 39120 26027 39172 26036
rect 39120 25993 39129 26027
rect 39129 25993 39163 26027
rect 39163 25993 39172 26027
rect 39120 25984 39172 25993
rect 45284 25984 45336 26036
rect 46020 25984 46072 26036
rect 46940 26027 46992 26036
rect 46940 25993 46949 26027
rect 46949 25993 46983 26027
rect 46983 25993 46992 26027
rect 46940 25984 46992 25993
rect 48780 25984 48832 26036
rect 37372 25916 37424 25968
rect 36912 25891 36964 25900
rect 36912 25857 36921 25891
rect 36921 25857 36955 25891
rect 36955 25857 36964 25891
rect 36912 25848 36964 25857
rect 37096 25848 37148 25900
rect 37648 25916 37700 25968
rect 37740 25891 37792 25900
rect 37740 25857 37749 25891
rect 37749 25857 37783 25891
rect 37783 25857 37792 25891
rect 37740 25848 37792 25857
rect 38844 25916 38896 25968
rect 39212 25897 39264 25900
rect 39212 25863 39221 25897
rect 39221 25863 39255 25897
rect 39255 25863 39264 25897
rect 40408 25916 40460 25968
rect 39212 25848 39264 25863
rect 42892 25848 42944 25900
rect 44456 25848 44508 25900
rect 45928 25916 45980 25968
rect 36544 25780 36596 25832
rect 10324 25712 10376 25764
rect 12164 25712 12216 25764
rect 12624 25712 12676 25764
rect 13176 25712 13228 25764
rect 13452 25712 13504 25764
rect 10140 25644 10192 25696
rect 11152 25644 11204 25696
rect 12348 25687 12400 25696
rect 12348 25653 12357 25687
rect 12357 25653 12391 25687
rect 12391 25653 12400 25687
rect 12348 25644 12400 25653
rect 31116 25712 31168 25764
rect 44088 25712 44140 25764
rect 45192 25780 45244 25832
rect 45560 25848 45612 25900
rect 46480 25780 46532 25832
rect 46296 25755 46348 25764
rect 46296 25721 46305 25755
rect 46305 25721 46339 25755
rect 46339 25721 46348 25755
rect 46296 25712 46348 25721
rect 47952 25848 48004 25900
rect 48044 25891 48096 25900
rect 48044 25857 48053 25891
rect 48053 25857 48087 25891
rect 48087 25857 48096 25891
rect 48044 25848 48096 25857
rect 48228 25959 48280 25968
rect 48228 25925 48237 25959
rect 48237 25925 48271 25959
rect 48271 25925 48280 25959
rect 48228 25916 48280 25925
rect 48412 25848 48464 25900
rect 47676 25780 47728 25832
rect 47860 25712 47912 25764
rect 51264 25984 51316 26036
rect 52736 25984 52788 26036
rect 53472 25984 53524 26036
rect 54208 25984 54260 26036
rect 55312 26027 55364 26036
rect 55312 25993 55321 26027
rect 55321 25993 55355 26027
rect 55355 25993 55364 26027
rect 55312 25984 55364 25993
rect 57060 25984 57112 26036
rect 58256 25984 58308 26036
rect 50804 25916 50856 25968
rect 51080 25891 51132 25900
rect 51080 25857 51089 25891
rect 51089 25857 51123 25891
rect 51123 25857 51132 25891
rect 51080 25848 51132 25857
rect 50160 25823 50212 25832
rect 50160 25789 50169 25823
rect 50169 25789 50203 25823
rect 50203 25789 50212 25823
rect 51356 25891 51408 25900
rect 51356 25857 51390 25891
rect 51390 25857 51408 25891
rect 51356 25848 51408 25857
rect 52460 25848 52512 25900
rect 53840 25916 53892 25968
rect 55404 25848 55456 25900
rect 50160 25780 50212 25789
rect 53196 25780 53248 25832
rect 56784 25848 56836 25900
rect 57980 25916 58032 25968
rect 56324 25780 56376 25832
rect 56508 25780 56560 25832
rect 56968 25823 57020 25832
rect 56968 25789 56977 25823
rect 56977 25789 57011 25823
rect 57011 25789 57020 25823
rect 56968 25780 57020 25789
rect 58624 25848 58676 25900
rect 49148 25712 49200 25764
rect 56876 25712 56928 25764
rect 37740 25644 37792 25696
rect 39396 25644 39448 25696
rect 41420 25644 41472 25696
rect 41604 25644 41656 25696
rect 42708 25644 42760 25696
rect 49424 25644 49476 25696
rect 49792 25687 49844 25696
rect 49792 25653 49801 25687
rect 49801 25653 49835 25687
rect 49835 25653 49844 25687
rect 49792 25644 49844 25653
rect 52736 25687 52788 25696
rect 52736 25653 52745 25687
rect 52745 25653 52779 25687
rect 52779 25653 52788 25687
rect 52736 25644 52788 25653
rect 58072 25687 58124 25696
rect 58072 25653 58081 25687
rect 58081 25653 58115 25687
rect 58115 25653 58124 25687
rect 58072 25644 58124 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3424 25483 3476 25492
rect 3424 25449 3433 25483
rect 3433 25449 3467 25483
rect 3467 25449 3476 25483
rect 3424 25440 3476 25449
rect 3792 25440 3844 25492
rect 4068 25440 4120 25492
rect 4620 25440 4672 25492
rect 5724 25483 5776 25492
rect 5724 25449 5733 25483
rect 5733 25449 5767 25483
rect 5767 25449 5776 25483
rect 5724 25440 5776 25449
rect 5816 25440 5868 25492
rect 7472 25483 7524 25492
rect 7472 25449 7481 25483
rect 7481 25449 7515 25483
rect 7515 25449 7524 25483
rect 7472 25440 7524 25449
rect 8760 25483 8812 25492
rect 8760 25449 8769 25483
rect 8769 25449 8803 25483
rect 8803 25449 8812 25483
rect 8760 25440 8812 25449
rect 9772 25440 9824 25492
rect 10416 25440 10468 25492
rect 11888 25440 11940 25492
rect 3332 25372 3384 25424
rect 3240 25304 3292 25356
rect 3700 25304 3752 25356
rect 4068 25279 4120 25288
rect 4068 25245 4077 25279
rect 4077 25245 4111 25279
rect 4111 25245 4120 25279
rect 4068 25236 4120 25245
rect 4712 25236 4764 25288
rect 4804 25279 4856 25288
rect 4804 25245 4813 25279
rect 4813 25245 4847 25279
rect 4847 25245 4856 25279
rect 4804 25236 4856 25245
rect 5172 25236 5224 25288
rect 5632 25236 5684 25288
rect 7288 25372 7340 25424
rect 9128 25372 9180 25424
rect 11152 25372 11204 25424
rect 12532 25483 12584 25492
rect 12532 25449 12541 25483
rect 12541 25449 12575 25483
rect 12575 25449 12584 25483
rect 13084 25483 13136 25492
rect 12532 25440 12584 25449
rect 13084 25449 13093 25483
rect 13093 25449 13127 25483
rect 13127 25449 13136 25483
rect 13084 25440 13136 25449
rect 13636 25440 13688 25492
rect 25320 25440 25372 25492
rect 36544 25440 36596 25492
rect 36912 25440 36964 25492
rect 37464 25440 37516 25492
rect 38568 25440 38620 25492
rect 40408 25440 40460 25492
rect 7196 25236 7248 25288
rect 7288 25279 7340 25288
rect 7288 25245 7297 25279
rect 7297 25245 7331 25279
rect 7331 25245 7340 25279
rect 7288 25236 7340 25245
rect 8576 25347 8628 25356
rect 8576 25313 8585 25347
rect 8585 25313 8619 25347
rect 8619 25313 8628 25347
rect 8576 25304 8628 25313
rect 7932 25236 7984 25288
rect 8484 25279 8536 25288
rect 8484 25245 8493 25279
rect 8493 25245 8527 25279
rect 8527 25245 8536 25279
rect 9680 25304 9732 25356
rect 12072 25304 12124 25356
rect 8484 25236 8536 25245
rect 4712 25143 4764 25152
rect 4712 25109 4721 25143
rect 4721 25109 4755 25143
rect 4755 25109 4764 25143
rect 4712 25100 4764 25109
rect 5448 25100 5500 25152
rect 5540 25143 5592 25152
rect 5540 25109 5549 25143
rect 5549 25109 5583 25143
rect 5583 25109 5592 25143
rect 5540 25100 5592 25109
rect 8024 25168 8076 25220
rect 8300 25143 8352 25152
rect 8300 25109 8309 25143
rect 8309 25109 8343 25143
rect 8343 25109 8352 25143
rect 8300 25100 8352 25109
rect 8852 25168 8904 25220
rect 9864 25211 9916 25220
rect 9864 25177 9873 25211
rect 9873 25177 9907 25211
rect 9907 25177 9916 25211
rect 9864 25168 9916 25177
rect 10232 25168 10284 25220
rect 10324 25143 10376 25152
rect 10324 25109 10333 25143
rect 10333 25109 10367 25143
rect 10367 25109 10376 25143
rect 10324 25100 10376 25109
rect 12716 25168 12768 25220
rect 13084 25279 13136 25288
rect 13084 25245 13093 25279
rect 13093 25245 13127 25279
rect 13127 25245 13136 25279
rect 13084 25236 13136 25245
rect 12532 25100 12584 25152
rect 36820 25279 36872 25288
rect 36820 25245 36829 25279
rect 36829 25245 36863 25279
rect 36863 25245 36872 25279
rect 36820 25236 36872 25245
rect 37648 25372 37700 25424
rect 41420 25483 41472 25492
rect 41420 25449 41429 25483
rect 41429 25449 41463 25483
rect 41463 25449 41472 25483
rect 41420 25440 41472 25449
rect 42248 25440 42300 25492
rect 42616 25440 42668 25492
rect 40776 25415 40828 25424
rect 40776 25381 40785 25415
rect 40785 25381 40819 25415
rect 40819 25381 40828 25415
rect 40776 25372 40828 25381
rect 41512 25372 41564 25424
rect 44088 25440 44140 25492
rect 47308 25440 47360 25492
rect 47952 25440 48004 25492
rect 48136 25440 48188 25492
rect 48412 25440 48464 25492
rect 51356 25483 51408 25492
rect 51356 25449 51365 25483
rect 51365 25449 51399 25483
rect 51399 25449 51408 25483
rect 51356 25440 51408 25449
rect 51632 25440 51684 25492
rect 52736 25440 52788 25492
rect 53104 25440 53156 25492
rect 53748 25440 53800 25492
rect 13452 25143 13504 25152
rect 13452 25109 13461 25143
rect 13461 25109 13495 25143
rect 13495 25109 13504 25143
rect 13452 25100 13504 25109
rect 37464 25279 37516 25288
rect 37464 25245 37473 25279
rect 37473 25245 37507 25279
rect 37507 25245 37516 25279
rect 37464 25236 37516 25245
rect 37648 25279 37700 25288
rect 37648 25245 37657 25279
rect 37657 25245 37691 25279
rect 37691 25245 37700 25279
rect 37648 25236 37700 25245
rect 37832 25279 37884 25288
rect 37832 25245 37841 25279
rect 37841 25245 37875 25279
rect 37875 25245 37884 25279
rect 37832 25236 37884 25245
rect 38936 25279 38988 25288
rect 38936 25245 38945 25279
rect 38945 25245 38979 25279
rect 38979 25245 38988 25279
rect 38936 25236 38988 25245
rect 40592 25304 40644 25356
rect 40040 25279 40092 25288
rect 40040 25245 40049 25279
rect 40049 25245 40083 25279
rect 40083 25245 40092 25279
rect 40040 25236 40092 25245
rect 39212 25100 39264 25152
rect 41604 25236 41656 25288
rect 41696 25279 41748 25288
rect 41696 25245 41705 25279
rect 41705 25245 41739 25279
rect 41739 25245 41748 25279
rect 41696 25236 41748 25245
rect 41880 25279 41932 25288
rect 41880 25245 41889 25279
rect 41889 25245 41923 25279
rect 41923 25245 41932 25279
rect 41880 25236 41932 25245
rect 42524 25347 42576 25356
rect 42524 25313 42533 25347
rect 42533 25313 42567 25347
rect 42567 25313 42576 25347
rect 42524 25304 42576 25313
rect 44088 25236 44140 25288
rect 41052 25168 41104 25220
rect 41788 25211 41840 25220
rect 41788 25177 41797 25211
rect 41797 25177 41831 25211
rect 41831 25177 41840 25211
rect 41788 25168 41840 25177
rect 42800 25211 42852 25220
rect 42800 25177 42809 25211
rect 42809 25177 42843 25211
rect 42843 25177 42852 25211
rect 42800 25168 42852 25177
rect 44824 25236 44876 25288
rect 45284 25236 45336 25288
rect 45928 25279 45980 25288
rect 45928 25245 45937 25279
rect 45937 25245 45971 25279
rect 45971 25245 45980 25279
rect 45928 25236 45980 25245
rect 46020 25279 46072 25288
rect 46020 25245 46029 25279
rect 46029 25245 46063 25279
rect 46063 25245 46072 25279
rect 46020 25236 46072 25245
rect 40960 25143 41012 25152
rect 40960 25109 40987 25143
rect 40987 25109 41012 25143
rect 40960 25100 41012 25109
rect 42892 25100 42944 25152
rect 45008 25143 45060 25152
rect 45008 25109 45017 25143
rect 45017 25109 45051 25143
rect 45051 25109 45060 25143
rect 45008 25100 45060 25109
rect 45560 25168 45612 25220
rect 46296 25236 46348 25288
rect 49424 25372 49476 25424
rect 46848 25347 46900 25356
rect 46848 25313 46857 25347
rect 46857 25313 46891 25347
rect 46891 25313 46900 25347
rect 46848 25304 46900 25313
rect 46949 25347 47001 25356
rect 46949 25313 46983 25347
rect 46983 25313 47001 25347
rect 46949 25304 47001 25313
rect 46204 25100 46256 25152
rect 46388 25143 46440 25152
rect 46388 25109 46397 25143
rect 46397 25109 46431 25143
rect 46431 25109 46440 25143
rect 46388 25100 46440 25109
rect 47032 25168 47084 25220
rect 48872 25236 48924 25288
rect 54852 25372 54904 25424
rect 53380 25279 53432 25288
rect 53380 25245 53389 25279
rect 53389 25245 53423 25279
rect 53423 25245 53432 25279
rect 53380 25236 53432 25245
rect 54484 25304 54536 25356
rect 53748 25279 53800 25288
rect 53748 25245 53757 25279
rect 53757 25245 53791 25279
rect 53791 25245 53800 25279
rect 53748 25236 53800 25245
rect 47400 25100 47452 25152
rect 48596 25100 48648 25152
rect 49148 25100 49200 25152
rect 53840 25168 53892 25220
rect 54300 25236 54352 25288
rect 54944 25304 54996 25356
rect 53472 25143 53524 25152
rect 53472 25109 53481 25143
rect 53481 25109 53515 25143
rect 53515 25109 53524 25143
rect 53472 25100 53524 25109
rect 56232 25236 56284 25288
rect 57152 25279 57204 25288
rect 57152 25245 57161 25279
rect 57161 25245 57195 25279
rect 57195 25245 57204 25279
rect 57152 25236 57204 25245
rect 57980 25304 58032 25356
rect 58072 25304 58124 25356
rect 55036 25168 55088 25220
rect 56600 25168 56652 25220
rect 58624 25168 58676 25220
rect 55312 25143 55364 25152
rect 55312 25109 55321 25143
rect 55321 25109 55355 25143
rect 55355 25109 55364 25143
rect 55312 25100 55364 25109
rect 57428 25143 57480 25152
rect 57428 25109 57437 25143
rect 57437 25109 57471 25143
rect 57471 25109 57480 25143
rect 57428 25100 57480 25109
rect 57612 25100 57664 25152
rect 57796 25100 57848 25152
rect 58072 25143 58124 25152
rect 58072 25109 58081 25143
rect 58081 25109 58115 25143
rect 58115 25109 58124 25143
rect 58072 25100 58124 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 3700 24896 3752 24948
rect 5724 24896 5776 24948
rect 12532 24896 12584 24948
rect 12624 24939 12676 24948
rect 12624 24905 12633 24939
rect 12633 24905 12667 24939
rect 12667 24905 12676 24939
rect 12624 24896 12676 24905
rect 13084 24896 13136 24948
rect 38936 24939 38988 24948
rect 38936 24905 38945 24939
rect 38945 24905 38979 24939
rect 38979 24905 38988 24939
rect 38936 24896 38988 24905
rect 40040 24896 40092 24948
rect 41052 24896 41104 24948
rect 41880 24896 41932 24948
rect 42708 24939 42760 24948
rect 42708 24905 42717 24939
rect 42717 24905 42751 24939
rect 42751 24905 42760 24939
rect 42708 24896 42760 24905
rect 42800 24939 42852 24948
rect 42800 24905 42809 24939
rect 42809 24905 42843 24939
rect 42843 24905 42852 24939
rect 42800 24896 42852 24905
rect 45008 24896 45060 24948
rect 45744 24896 45796 24948
rect 5448 24828 5500 24880
rect 10048 24828 10100 24880
rect 13452 24871 13504 24880
rect 13452 24837 13486 24871
rect 13486 24837 13504 24871
rect 13452 24828 13504 24837
rect 2688 24803 2740 24812
rect 2688 24769 2697 24803
rect 2697 24769 2731 24803
rect 2731 24769 2740 24803
rect 2688 24760 2740 24769
rect 940 24692 992 24744
rect 3700 24735 3752 24744
rect 3700 24701 3709 24735
rect 3709 24701 3743 24735
rect 3743 24701 3752 24735
rect 3700 24692 3752 24701
rect 7288 24692 7340 24744
rect 11336 24692 11388 24744
rect 7840 24624 7892 24676
rect 11888 24624 11940 24676
rect 12992 24760 13044 24812
rect 36820 24760 36872 24812
rect 37372 24760 37424 24812
rect 12716 24692 12768 24744
rect 37188 24692 37240 24744
rect 38476 24803 38528 24812
rect 38476 24769 38485 24803
rect 38485 24769 38519 24803
rect 38519 24769 38528 24803
rect 38476 24760 38528 24769
rect 39028 24803 39080 24812
rect 39028 24769 39037 24803
rect 39037 24769 39071 24803
rect 39071 24769 39080 24803
rect 39028 24760 39080 24769
rect 39764 24803 39816 24812
rect 39764 24769 39773 24803
rect 39773 24769 39807 24803
rect 39807 24769 39816 24803
rect 39764 24760 39816 24769
rect 3056 24556 3108 24608
rect 9680 24556 9732 24608
rect 10600 24556 10652 24608
rect 12532 24624 12584 24676
rect 37372 24624 37424 24676
rect 40684 24803 40736 24812
rect 40684 24769 40693 24803
rect 40693 24769 40727 24803
rect 40727 24769 40736 24803
rect 40684 24760 40736 24769
rect 40960 24760 41012 24812
rect 42892 24828 42944 24880
rect 41512 24803 41564 24812
rect 41512 24769 41521 24803
rect 41521 24769 41555 24803
rect 41555 24769 41564 24803
rect 41512 24760 41564 24769
rect 41604 24760 41656 24812
rect 43812 24803 43864 24812
rect 43812 24769 43821 24803
rect 43821 24769 43855 24803
rect 43855 24769 43864 24803
rect 43812 24760 43864 24769
rect 44180 24803 44232 24812
rect 44180 24769 44189 24803
rect 44189 24769 44223 24803
rect 44223 24769 44232 24803
rect 44180 24760 44232 24769
rect 44364 24760 44416 24812
rect 44456 24803 44508 24812
rect 44456 24769 44465 24803
rect 44465 24769 44499 24803
rect 44499 24769 44508 24803
rect 44456 24760 44508 24769
rect 44548 24803 44600 24812
rect 44548 24769 44557 24803
rect 44557 24769 44591 24803
rect 44591 24769 44600 24803
rect 44548 24760 44600 24769
rect 45192 24760 45244 24812
rect 45376 24760 45428 24812
rect 46204 24828 46256 24880
rect 46388 24803 46440 24812
rect 46388 24769 46397 24803
rect 46397 24769 46431 24803
rect 46431 24769 46440 24803
rect 46388 24760 46440 24769
rect 45008 24692 45060 24744
rect 46664 24803 46716 24812
rect 46664 24769 46673 24803
rect 46673 24769 46707 24803
rect 46707 24769 46716 24803
rect 46664 24760 46716 24769
rect 47032 24828 47084 24880
rect 47676 24828 47728 24880
rect 47216 24803 47268 24812
rect 47216 24769 47225 24803
rect 47225 24769 47259 24803
rect 47259 24769 47268 24803
rect 47216 24760 47268 24769
rect 47400 24803 47452 24812
rect 47400 24769 47409 24803
rect 47409 24769 47443 24803
rect 47443 24769 47452 24803
rect 48780 24896 48832 24948
rect 48412 24828 48464 24880
rect 49240 24828 49292 24880
rect 53104 24896 53156 24948
rect 53472 24896 53524 24948
rect 53748 24939 53800 24948
rect 53748 24905 53757 24939
rect 53757 24905 53791 24939
rect 53791 24905 53800 24939
rect 53748 24896 53800 24905
rect 57428 24896 57480 24948
rect 58072 24896 58124 24948
rect 47400 24760 47452 24769
rect 13176 24556 13228 24608
rect 35900 24556 35952 24608
rect 36728 24556 36780 24608
rect 37280 24599 37332 24608
rect 37280 24565 37289 24599
rect 37289 24565 37323 24599
rect 37323 24565 37332 24599
rect 37280 24556 37332 24565
rect 38016 24599 38068 24608
rect 38016 24565 38025 24599
rect 38025 24565 38059 24599
rect 38059 24565 38068 24599
rect 38016 24556 38068 24565
rect 42248 24556 42300 24608
rect 43996 24624 44048 24676
rect 45652 24624 45704 24676
rect 45836 24667 45888 24676
rect 45836 24633 45845 24667
rect 45845 24633 45879 24667
rect 45879 24633 45888 24667
rect 47492 24692 47544 24744
rect 48228 24803 48280 24812
rect 48228 24769 48237 24803
rect 48237 24769 48271 24803
rect 48271 24769 48280 24803
rect 48228 24760 48280 24769
rect 48504 24760 48556 24812
rect 48596 24735 48648 24744
rect 48596 24701 48605 24735
rect 48605 24701 48639 24735
rect 48639 24701 48648 24735
rect 48596 24692 48648 24701
rect 48964 24735 49016 24744
rect 48964 24701 48973 24735
rect 48973 24701 49007 24735
rect 49007 24701 49016 24735
rect 48964 24692 49016 24701
rect 45836 24624 45888 24633
rect 51632 24803 51684 24812
rect 51632 24769 51641 24803
rect 51641 24769 51675 24803
rect 51675 24769 51684 24803
rect 52460 24828 52512 24880
rect 51632 24760 51684 24769
rect 51816 24803 51868 24812
rect 51816 24769 51825 24803
rect 51825 24769 51859 24803
rect 51859 24769 51868 24803
rect 51816 24760 51868 24769
rect 52092 24803 52144 24812
rect 52092 24769 52101 24803
rect 52101 24769 52135 24803
rect 52135 24769 52144 24803
rect 52092 24760 52144 24769
rect 45376 24556 45428 24608
rect 45468 24599 45520 24608
rect 45468 24565 45477 24599
rect 45477 24565 45511 24599
rect 45511 24565 45520 24599
rect 45468 24556 45520 24565
rect 46204 24556 46256 24608
rect 47124 24556 47176 24608
rect 48412 24599 48464 24608
rect 48412 24565 48421 24599
rect 48421 24565 48455 24599
rect 48455 24565 48464 24599
rect 48412 24556 48464 24565
rect 53380 24760 53432 24812
rect 53564 24760 53616 24812
rect 51080 24556 51132 24608
rect 51448 24556 51500 24608
rect 51724 24599 51776 24608
rect 51724 24565 51733 24599
rect 51733 24565 51767 24599
rect 51767 24565 51776 24599
rect 51724 24556 51776 24565
rect 52368 24556 52420 24608
rect 54760 24735 54812 24744
rect 54760 24701 54769 24735
rect 54769 24701 54803 24735
rect 54803 24701 54812 24735
rect 54760 24692 54812 24701
rect 55128 24760 55180 24812
rect 54852 24556 54904 24608
rect 56048 24624 56100 24676
rect 57980 24692 58032 24744
rect 55312 24556 55364 24608
rect 55956 24556 56008 24608
rect 57060 24599 57112 24608
rect 57060 24565 57069 24599
rect 57069 24565 57103 24599
rect 57103 24565 57112 24599
rect 57060 24556 57112 24565
rect 57888 24599 57940 24608
rect 57888 24565 57897 24599
rect 57897 24565 57931 24599
rect 57931 24565 57940 24599
rect 57888 24556 57940 24565
rect 58716 24556 58768 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3056 24352 3108 24404
rect 3332 24395 3384 24404
rect 3332 24361 3341 24395
rect 3341 24361 3375 24395
rect 3375 24361 3384 24395
rect 3332 24352 3384 24361
rect 3700 24352 3752 24404
rect 6736 24352 6788 24404
rect 4896 24327 4948 24336
rect 4896 24293 4905 24327
rect 4905 24293 4939 24327
rect 4939 24293 4948 24327
rect 4896 24284 4948 24293
rect 3148 24259 3200 24268
rect 3148 24225 3157 24259
rect 3157 24225 3191 24259
rect 3191 24225 3200 24259
rect 3148 24216 3200 24225
rect 3240 24191 3292 24200
rect 3240 24157 3249 24191
rect 3249 24157 3283 24191
rect 3283 24157 3292 24191
rect 3240 24148 3292 24157
rect 4344 24191 4396 24200
rect 4344 24157 4353 24191
rect 4353 24157 4387 24191
rect 4387 24157 4396 24191
rect 4344 24148 4396 24157
rect 2412 24080 2464 24132
rect 2872 24080 2924 24132
rect 3332 24080 3384 24132
rect 4712 24191 4764 24200
rect 4712 24157 4721 24191
rect 4721 24157 4755 24191
rect 4755 24157 4764 24191
rect 4712 24148 4764 24157
rect 5724 24148 5776 24200
rect 6552 24148 6604 24200
rect 9680 24352 9732 24404
rect 9956 24352 10008 24404
rect 7656 24327 7708 24336
rect 7656 24293 7665 24327
rect 7665 24293 7699 24327
rect 7699 24293 7708 24327
rect 7656 24284 7708 24293
rect 8484 24327 8536 24336
rect 8484 24293 8493 24327
rect 8493 24293 8527 24327
rect 8527 24293 8536 24327
rect 8484 24284 8536 24293
rect 7012 24191 7064 24200
rect 7012 24157 7021 24191
rect 7021 24157 7055 24191
rect 7055 24157 7064 24191
rect 7012 24148 7064 24157
rect 7380 24191 7432 24200
rect 7380 24157 7389 24191
rect 7389 24157 7423 24191
rect 7423 24157 7432 24191
rect 7380 24148 7432 24157
rect 5264 24080 5316 24132
rect 2688 24012 2740 24064
rect 4620 24012 4672 24064
rect 6368 24012 6420 24064
rect 7564 24080 7616 24132
rect 7840 24080 7892 24132
rect 8208 24191 8260 24200
rect 8208 24157 8217 24191
rect 8217 24157 8251 24191
rect 8251 24157 8260 24191
rect 8208 24148 8260 24157
rect 8300 24191 8352 24200
rect 8300 24157 8309 24191
rect 8309 24157 8343 24191
rect 8343 24157 8352 24191
rect 8300 24148 8352 24157
rect 10048 24191 10100 24200
rect 10048 24157 10057 24191
rect 10057 24157 10091 24191
rect 10091 24157 10100 24191
rect 10048 24148 10100 24157
rect 10140 24191 10192 24200
rect 10140 24157 10149 24191
rect 10149 24157 10183 24191
rect 10183 24157 10192 24191
rect 10140 24148 10192 24157
rect 10508 24191 10560 24200
rect 10508 24157 10517 24191
rect 10517 24157 10551 24191
rect 10551 24157 10560 24191
rect 10508 24148 10560 24157
rect 12440 24352 12492 24404
rect 12900 24352 12952 24404
rect 13636 24352 13688 24404
rect 37188 24352 37240 24404
rect 39028 24352 39080 24404
rect 40040 24352 40092 24404
rect 43812 24352 43864 24404
rect 45008 24352 45060 24404
rect 45468 24352 45520 24404
rect 47124 24395 47176 24404
rect 47124 24361 47133 24395
rect 47133 24361 47167 24395
rect 47167 24361 47176 24395
rect 47124 24352 47176 24361
rect 47584 24352 47636 24404
rect 48228 24352 48280 24404
rect 48872 24352 48924 24404
rect 48964 24352 49016 24404
rect 51724 24352 51776 24404
rect 51816 24352 51868 24404
rect 52092 24352 52144 24404
rect 56692 24352 56744 24404
rect 57060 24352 57112 24404
rect 57888 24352 57940 24404
rect 13820 24327 13872 24336
rect 13820 24293 13829 24327
rect 13829 24293 13863 24327
rect 13863 24293 13872 24327
rect 13820 24284 13872 24293
rect 9772 24055 9824 24064
rect 9772 24021 9781 24055
rect 9781 24021 9815 24055
rect 9815 24021 9824 24055
rect 9772 24012 9824 24021
rect 10324 24012 10376 24064
rect 10600 24012 10652 24064
rect 11428 24012 11480 24064
rect 12716 24191 12768 24200
rect 12716 24157 12725 24191
rect 12725 24157 12759 24191
rect 12759 24157 12768 24191
rect 12716 24148 12768 24157
rect 12900 24148 12952 24200
rect 13360 24148 13412 24200
rect 34520 24216 34572 24268
rect 35440 24216 35492 24268
rect 37832 24216 37884 24268
rect 12624 24080 12676 24132
rect 12992 24080 13044 24132
rect 12532 24012 12584 24064
rect 12716 24055 12768 24064
rect 12716 24021 12725 24055
rect 12725 24021 12759 24055
rect 12759 24021 12768 24055
rect 37556 24191 37608 24200
rect 37556 24157 37565 24191
rect 37565 24157 37599 24191
rect 37599 24157 37608 24191
rect 37556 24148 37608 24157
rect 38568 24148 38620 24200
rect 39120 24191 39172 24200
rect 39120 24157 39129 24191
rect 39129 24157 39163 24191
rect 39163 24157 39172 24191
rect 39120 24148 39172 24157
rect 35440 24123 35492 24132
rect 35440 24089 35449 24123
rect 35449 24089 35483 24123
rect 35483 24089 35492 24123
rect 35440 24080 35492 24089
rect 35900 24080 35952 24132
rect 39396 24191 39448 24200
rect 39396 24157 39405 24191
rect 39405 24157 39439 24191
rect 39439 24157 39448 24191
rect 39396 24148 39448 24157
rect 42156 24216 42208 24268
rect 44088 24284 44140 24336
rect 39764 24148 39816 24200
rect 12716 24012 12768 24021
rect 13636 24055 13688 24064
rect 13636 24021 13645 24055
rect 13645 24021 13679 24055
rect 13679 24021 13688 24055
rect 13636 24012 13688 24021
rect 37004 24055 37056 24064
rect 37004 24021 37013 24055
rect 37013 24021 37047 24055
rect 37047 24021 37056 24055
rect 37004 24012 37056 24021
rect 38384 24012 38436 24064
rect 41328 24191 41380 24200
rect 41328 24157 41337 24191
rect 41337 24157 41371 24191
rect 41371 24157 41380 24191
rect 41328 24148 41380 24157
rect 42708 24148 42760 24200
rect 43904 24216 43956 24268
rect 41604 24123 41656 24132
rect 41604 24089 41613 24123
rect 41613 24089 41647 24123
rect 41647 24089 41656 24123
rect 41604 24080 41656 24089
rect 43904 24080 43956 24132
rect 44088 24080 44140 24132
rect 43444 24055 43496 24064
rect 43444 24021 43453 24055
rect 43453 24021 43487 24055
rect 43487 24021 43496 24055
rect 43444 24012 43496 24021
rect 44272 24012 44324 24064
rect 45284 24191 45336 24200
rect 45284 24157 45293 24191
rect 45293 24157 45327 24191
rect 45327 24157 45336 24191
rect 45284 24148 45336 24157
rect 51632 24284 51684 24336
rect 45652 24148 45704 24200
rect 48136 24216 48188 24268
rect 48780 24259 48832 24268
rect 48780 24225 48789 24259
rect 48789 24225 48823 24259
rect 48823 24225 48832 24259
rect 48780 24216 48832 24225
rect 55036 24284 55088 24336
rect 45100 24123 45152 24132
rect 45100 24089 45109 24123
rect 45109 24089 45143 24123
rect 45143 24089 45152 24123
rect 45100 24080 45152 24089
rect 47676 24148 47728 24200
rect 47492 24080 47544 24132
rect 48596 24148 48648 24200
rect 48964 24148 49016 24200
rect 50620 24148 50672 24200
rect 51448 24191 51500 24200
rect 51448 24157 51457 24191
rect 51457 24157 51491 24191
rect 51491 24157 51500 24191
rect 51448 24148 51500 24157
rect 47216 24012 47268 24064
rect 47676 24012 47728 24064
rect 48136 24055 48188 24064
rect 48136 24021 48145 24055
rect 48145 24021 48179 24055
rect 48179 24021 48188 24055
rect 48136 24012 48188 24021
rect 51080 24080 51132 24132
rect 52276 24148 52328 24200
rect 53288 24148 53340 24200
rect 53380 24148 53432 24200
rect 55956 24259 56008 24268
rect 55956 24225 55965 24259
rect 55965 24225 55999 24259
rect 55999 24225 56008 24259
rect 55956 24216 56008 24225
rect 56232 24284 56284 24336
rect 50620 24055 50672 24064
rect 50620 24021 50629 24055
rect 50629 24021 50663 24055
rect 50663 24021 50672 24055
rect 50620 24012 50672 24021
rect 50712 24012 50764 24064
rect 51356 24055 51408 24064
rect 51356 24021 51365 24055
rect 51365 24021 51399 24055
rect 51399 24021 51408 24055
rect 51356 24012 51408 24021
rect 51908 24012 51960 24064
rect 52920 24055 52972 24064
rect 52920 24021 52929 24055
rect 52929 24021 52963 24055
rect 52963 24021 52972 24055
rect 52920 24012 52972 24021
rect 54208 24012 54260 24064
rect 56508 24148 56560 24200
rect 57428 24148 57480 24200
rect 58164 24191 58216 24200
rect 58164 24157 58173 24191
rect 58173 24157 58207 24191
rect 58207 24157 58216 24191
rect 58164 24148 58216 24157
rect 57980 24055 58032 24064
rect 57980 24021 57989 24055
rect 57989 24021 58023 24055
rect 58023 24021 58032 24055
rect 57980 24012 58032 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 2688 23808 2740 23860
rect 3240 23808 3292 23860
rect 4344 23808 4396 23860
rect 4896 23808 4948 23860
rect 7288 23808 7340 23860
rect 7656 23808 7708 23860
rect 7932 23808 7984 23860
rect 8208 23808 8260 23860
rect 8484 23808 8536 23860
rect 10048 23808 10100 23860
rect 10140 23851 10192 23860
rect 10140 23817 10149 23851
rect 10149 23817 10183 23851
rect 10183 23817 10192 23851
rect 10140 23808 10192 23817
rect 10508 23851 10560 23860
rect 10508 23817 10517 23851
rect 10517 23817 10551 23851
rect 10551 23817 10560 23851
rect 10508 23808 10560 23817
rect 11336 23808 11388 23860
rect 12256 23808 12308 23860
rect 13636 23808 13688 23860
rect 13820 23808 13872 23860
rect 35440 23808 35492 23860
rect 3976 23715 4028 23724
rect 3976 23681 3985 23715
rect 3985 23681 4019 23715
rect 4019 23681 4028 23715
rect 3976 23672 4028 23681
rect 4068 23715 4120 23724
rect 4068 23681 4077 23715
rect 4077 23681 4111 23715
rect 4111 23681 4120 23715
rect 4068 23672 4120 23681
rect 3884 23604 3936 23656
rect 10140 23715 10192 23724
rect 10140 23681 10149 23715
rect 10149 23681 10183 23715
rect 10183 23681 10192 23715
rect 10140 23672 10192 23681
rect 10968 23672 11020 23724
rect 8116 23647 8168 23656
rect 8116 23613 8125 23647
rect 8125 23613 8159 23647
rect 8159 23613 8168 23647
rect 8116 23604 8168 23613
rect 12164 23740 12216 23792
rect 11980 23647 12032 23656
rect 11980 23613 11989 23647
rect 11989 23613 12023 23647
rect 12023 23613 12032 23647
rect 11980 23604 12032 23613
rect 12808 23672 12860 23724
rect 12992 23672 13044 23724
rect 12256 23536 12308 23588
rect 12624 23536 12676 23588
rect 37004 23808 37056 23860
rect 37280 23808 37332 23860
rect 36820 23715 36872 23724
rect 36820 23681 36829 23715
rect 36829 23681 36863 23715
rect 36863 23681 36872 23715
rect 36820 23672 36872 23681
rect 37096 23672 37148 23724
rect 38016 23808 38068 23860
rect 38384 23808 38436 23860
rect 38476 23851 38528 23860
rect 38476 23817 38485 23851
rect 38485 23817 38519 23851
rect 38519 23817 38528 23851
rect 38476 23808 38528 23817
rect 38568 23808 38620 23860
rect 39120 23808 39172 23860
rect 41604 23808 41656 23860
rect 43812 23808 43864 23860
rect 49792 23808 49844 23860
rect 50528 23808 50580 23860
rect 50620 23808 50672 23860
rect 53840 23851 53892 23860
rect 53840 23817 53849 23851
rect 53849 23817 53883 23851
rect 53883 23817 53892 23851
rect 53840 23808 53892 23817
rect 54852 23808 54904 23860
rect 39396 23740 39448 23792
rect 43444 23740 43496 23792
rect 39396 23647 39448 23656
rect 39396 23613 39405 23647
rect 39405 23613 39439 23647
rect 39439 23613 39448 23647
rect 39396 23604 39448 23613
rect 43996 23672 44048 23724
rect 42248 23604 42300 23656
rect 46572 23647 46624 23656
rect 46572 23613 46581 23647
rect 46581 23613 46615 23647
rect 46615 23613 46624 23647
rect 46572 23604 46624 23613
rect 48964 23672 49016 23724
rect 52828 23740 52880 23792
rect 44640 23536 44692 23588
rect 49792 23604 49844 23656
rect 50068 23647 50120 23656
rect 50068 23613 50077 23647
rect 50077 23613 50111 23647
rect 50111 23613 50120 23647
rect 50068 23604 50120 23613
rect 50528 23715 50580 23724
rect 50528 23681 50537 23715
rect 50537 23681 50571 23715
rect 50571 23681 50580 23715
rect 50528 23672 50580 23681
rect 52736 23715 52788 23724
rect 52736 23681 52745 23715
rect 52745 23681 52779 23715
rect 52779 23681 52788 23715
rect 52736 23672 52788 23681
rect 52920 23715 52972 23724
rect 52920 23681 52929 23715
rect 52929 23681 52963 23715
rect 52963 23681 52972 23715
rect 52920 23672 52972 23681
rect 53932 23672 53984 23724
rect 54208 23715 54260 23724
rect 54208 23681 54217 23715
rect 54217 23681 54251 23715
rect 54251 23681 54260 23715
rect 54208 23672 54260 23681
rect 54300 23715 54352 23724
rect 54300 23681 54309 23715
rect 54309 23681 54343 23715
rect 54343 23681 54352 23715
rect 54300 23672 54352 23681
rect 54392 23715 54444 23724
rect 54392 23681 54401 23715
rect 54401 23681 54435 23715
rect 54435 23681 54444 23715
rect 54392 23672 54444 23681
rect 57980 23808 58032 23860
rect 54944 23715 54996 23724
rect 54944 23681 54953 23715
rect 54953 23681 54987 23715
rect 54987 23681 54996 23715
rect 54944 23672 54996 23681
rect 56508 23715 56560 23724
rect 56508 23681 56542 23715
rect 56542 23681 56560 23715
rect 56508 23672 56560 23681
rect 50344 23536 50396 23588
rect 50712 23536 50764 23588
rect 56232 23647 56284 23656
rect 56232 23613 56241 23647
rect 56241 23613 56275 23647
rect 56275 23613 56284 23647
rect 56232 23604 56284 23613
rect 4712 23468 4764 23520
rect 4804 23468 4856 23520
rect 7012 23468 7064 23520
rect 7932 23468 7984 23520
rect 10968 23511 11020 23520
rect 10968 23477 10977 23511
rect 10977 23477 11011 23511
rect 11011 23477 11020 23511
rect 10968 23468 11020 23477
rect 11888 23468 11940 23520
rect 12072 23511 12124 23520
rect 12072 23477 12081 23511
rect 12081 23477 12115 23511
rect 12115 23477 12124 23511
rect 12072 23468 12124 23477
rect 12532 23511 12584 23520
rect 12532 23477 12541 23511
rect 12541 23477 12575 23511
rect 12575 23477 12584 23511
rect 12532 23468 12584 23477
rect 37556 23468 37608 23520
rect 37740 23511 37792 23520
rect 37740 23477 37749 23511
rect 37749 23477 37783 23511
rect 37783 23477 37792 23511
rect 37740 23468 37792 23477
rect 40868 23511 40920 23520
rect 40868 23477 40877 23511
rect 40877 23477 40911 23511
rect 40911 23477 40920 23511
rect 40868 23468 40920 23477
rect 44364 23468 44416 23520
rect 45100 23468 45152 23520
rect 45928 23511 45980 23520
rect 45928 23477 45937 23511
rect 45937 23477 45971 23511
rect 45971 23477 45980 23511
rect 45928 23468 45980 23477
rect 48044 23511 48096 23520
rect 48044 23477 48053 23511
rect 48053 23477 48087 23511
rect 48087 23477 48096 23511
rect 48044 23468 48096 23477
rect 48596 23468 48648 23520
rect 49332 23468 49384 23520
rect 50620 23511 50672 23520
rect 50620 23477 50629 23511
rect 50629 23477 50663 23511
rect 50663 23477 50672 23511
rect 50620 23468 50672 23477
rect 54484 23511 54536 23520
rect 54484 23477 54493 23511
rect 54493 23477 54527 23511
rect 54527 23477 54536 23511
rect 54484 23468 54536 23477
rect 56600 23468 56652 23520
rect 57888 23511 57940 23520
rect 57888 23477 57897 23511
rect 57897 23477 57931 23511
rect 57931 23477 57940 23511
rect 57888 23468 57940 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4620 23264 4672 23316
rect 6828 23264 6880 23316
rect 7380 23264 7432 23316
rect 7932 23264 7984 23316
rect 8116 23264 8168 23316
rect 11888 23264 11940 23316
rect 39396 23264 39448 23316
rect 3516 23196 3568 23248
rect 4712 23128 4764 23180
rect 940 22992 992 23044
rect 1400 22924 1452 22976
rect 3884 23060 3936 23112
rect 6552 23060 6604 23112
rect 40224 23264 40276 23316
rect 42708 23307 42760 23316
rect 42708 23273 42717 23307
rect 42717 23273 42751 23307
rect 42751 23273 42760 23307
rect 42708 23264 42760 23273
rect 47308 23307 47360 23316
rect 47308 23273 47317 23307
rect 47317 23273 47351 23307
rect 47351 23273 47360 23307
rect 47308 23264 47360 23273
rect 7012 23060 7064 23112
rect 7840 23060 7892 23112
rect 8392 23060 8444 23112
rect 9956 23103 10008 23112
rect 9956 23069 9965 23103
rect 9965 23069 9999 23103
rect 9999 23069 10008 23103
rect 9956 23060 10008 23069
rect 10140 23103 10192 23112
rect 10140 23069 10149 23103
rect 10149 23069 10183 23103
rect 10183 23069 10192 23103
rect 10140 23060 10192 23069
rect 39396 23060 39448 23112
rect 41236 23060 41288 23112
rect 44180 23060 44232 23112
rect 46664 23196 46716 23248
rect 48596 23307 48648 23316
rect 48596 23273 48605 23307
rect 48605 23273 48639 23307
rect 48639 23273 48648 23307
rect 48596 23264 48648 23273
rect 48044 23196 48096 23248
rect 48228 23196 48280 23248
rect 49976 23264 50028 23316
rect 52736 23264 52788 23316
rect 56508 23307 56560 23316
rect 56508 23273 56517 23307
rect 56517 23273 56551 23307
rect 56551 23273 56560 23307
rect 56508 23264 56560 23273
rect 56784 23264 56836 23316
rect 47860 23060 47912 23112
rect 48964 23239 49016 23248
rect 48964 23205 48973 23239
rect 48973 23205 49007 23239
rect 49007 23205 49016 23239
rect 48964 23196 49016 23205
rect 49608 23196 49660 23248
rect 51172 23239 51224 23248
rect 51172 23205 51181 23239
rect 51181 23205 51215 23239
rect 51215 23205 51224 23239
rect 51172 23196 51224 23205
rect 50068 23128 50120 23180
rect 37740 23035 37792 23044
rect 37740 23001 37749 23035
rect 37749 23001 37783 23035
rect 37783 23001 37792 23035
rect 37740 22992 37792 23001
rect 39764 22992 39816 23044
rect 40132 23035 40184 23044
rect 40132 23001 40141 23035
rect 40141 23001 40175 23035
rect 40175 23001 40184 23035
rect 40132 22992 40184 23001
rect 3516 22967 3568 22976
rect 3516 22933 3525 22967
rect 3525 22933 3559 22967
rect 3559 22933 3568 22967
rect 3516 22924 3568 22933
rect 4712 22924 4764 22976
rect 6644 22967 6696 22976
rect 6644 22933 6653 22967
rect 6653 22933 6687 22967
rect 6687 22933 6696 22967
rect 6644 22924 6696 22933
rect 10140 22967 10192 22976
rect 10140 22933 10149 22967
rect 10149 22933 10183 22967
rect 10183 22933 10192 22967
rect 10140 22924 10192 22933
rect 12900 22967 12952 22976
rect 12900 22933 12909 22967
rect 12909 22933 12943 22967
rect 12943 22933 12952 22967
rect 12900 22924 12952 22933
rect 45284 23035 45336 23044
rect 45284 23001 45293 23035
rect 45293 23001 45327 23035
rect 45327 23001 45336 23035
rect 45284 22992 45336 23001
rect 46940 22992 46992 23044
rect 50344 23060 50396 23112
rect 52460 23196 52512 23248
rect 51356 23103 51408 23112
rect 51356 23069 51365 23103
rect 51365 23069 51399 23103
rect 51399 23069 51408 23103
rect 51356 23060 51408 23069
rect 50528 22992 50580 23044
rect 42248 22967 42300 22976
rect 42248 22933 42257 22967
rect 42257 22933 42291 22967
rect 42291 22933 42300 22967
rect 42248 22924 42300 22933
rect 47032 22967 47084 22976
rect 47032 22933 47041 22967
rect 47041 22933 47075 22967
rect 47075 22933 47084 22967
rect 47032 22924 47084 22933
rect 47952 22967 48004 22976
rect 47952 22933 47961 22967
rect 47961 22933 47995 22967
rect 47995 22933 48004 22967
rect 47952 22924 48004 22933
rect 50804 22967 50856 22976
rect 50804 22933 50813 22967
rect 50813 22933 50847 22967
rect 50847 22933 50856 22967
rect 50804 22924 50856 22933
rect 51448 22967 51500 22976
rect 51448 22933 51457 22967
rect 51457 22933 51491 22967
rect 51491 22933 51500 22967
rect 51448 22924 51500 22933
rect 51724 23035 51776 23044
rect 51724 23001 51733 23035
rect 51733 23001 51767 23035
rect 51767 23001 51776 23035
rect 51724 22992 51776 23001
rect 51908 23103 51960 23112
rect 51908 23069 51917 23103
rect 51917 23069 51951 23103
rect 51951 23069 51960 23103
rect 51908 23060 51960 23069
rect 52368 23103 52420 23112
rect 52368 23069 52377 23103
rect 52377 23069 52411 23103
rect 52411 23069 52420 23103
rect 52368 23060 52420 23069
rect 52460 23103 52512 23112
rect 52460 23069 52469 23103
rect 52469 23069 52503 23103
rect 52503 23069 52512 23103
rect 52460 23060 52512 23069
rect 52276 22967 52328 22976
rect 52276 22933 52285 22967
rect 52285 22933 52319 22967
rect 52319 22933 52328 22967
rect 52276 22924 52328 22933
rect 53472 23103 53524 23112
rect 53472 23069 53481 23103
rect 53481 23069 53515 23103
rect 53515 23069 53524 23103
rect 53472 23060 53524 23069
rect 54484 23060 54536 23112
rect 55312 23103 55364 23112
rect 55312 23069 55321 23103
rect 55321 23069 55355 23103
rect 55355 23069 55364 23103
rect 55312 23060 55364 23069
rect 57888 23196 57940 23248
rect 54392 22924 54444 22976
rect 57336 23103 57388 23112
rect 57336 23069 57345 23103
rect 57345 23069 57379 23103
rect 57379 23069 57388 23103
rect 57336 23060 57388 23069
rect 57520 23103 57572 23112
rect 57520 23069 57529 23103
rect 57529 23069 57563 23103
rect 57563 23069 57572 23103
rect 57520 23060 57572 23069
rect 57612 23103 57664 23112
rect 57612 23069 57621 23103
rect 57621 23069 57655 23103
rect 57655 23069 57664 23103
rect 57612 23060 57664 23069
rect 57980 23103 58032 23112
rect 57980 23069 57989 23103
rect 57989 23069 58023 23103
rect 58023 23069 58032 23103
rect 57980 23060 58032 23069
rect 58256 23103 58308 23112
rect 58256 23069 58265 23103
rect 58265 23069 58299 23103
rect 58299 23069 58308 23103
rect 58256 23060 58308 23069
rect 56048 22967 56100 22976
rect 56048 22933 56057 22967
rect 56057 22933 56091 22967
rect 56091 22933 56100 22967
rect 56048 22924 56100 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 1400 22763 1452 22772
rect 1400 22729 1409 22763
rect 1409 22729 1443 22763
rect 1443 22729 1452 22763
rect 1400 22720 1452 22729
rect 3516 22720 3568 22772
rect 3976 22720 4028 22772
rect 4160 22720 4212 22772
rect 8024 22720 8076 22772
rect 8392 22720 8444 22772
rect 9956 22763 10008 22772
rect 9956 22729 9965 22763
rect 9965 22729 9999 22763
rect 9999 22729 10008 22763
rect 9956 22720 10008 22729
rect 11888 22720 11940 22772
rect 2412 22652 2464 22704
rect 3148 22627 3200 22636
rect 3148 22593 3157 22627
rect 3157 22593 3191 22627
rect 3191 22593 3200 22627
rect 3148 22584 3200 22593
rect 3332 22516 3384 22568
rect 4712 22627 4764 22636
rect 4712 22593 4721 22627
rect 4721 22593 4755 22627
rect 4755 22593 4764 22627
rect 4712 22584 4764 22593
rect 7380 22584 7432 22636
rect 9312 22695 9364 22704
rect 9312 22661 9321 22695
rect 9321 22661 9355 22695
rect 9355 22661 9364 22695
rect 9312 22652 9364 22661
rect 5356 22516 5408 22568
rect 7012 22516 7064 22568
rect 9220 22584 9272 22636
rect 9680 22584 9732 22636
rect 4804 22448 4856 22500
rect 10784 22584 10836 22636
rect 12440 22627 12492 22636
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 12716 22627 12768 22636
rect 12716 22593 12725 22627
rect 12725 22593 12759 22627
rect 12759 22593 12768 22627
rect 12716 22584 12768 22593
rect 12808 22627 12860 22636
rect 12808 22593 12817 22627
rect 12817 22593 12851 22627
rect 12851 22593 12860 22627
rect 12808 22584 12860 22593
rect 12992 22627 13044 22636
rect 12992 22593 13001 22627
rect 13001 22593 13035 22627
rect 13035 22593 13044 22627
rect 12992 22584 13044 22593
rect 9956 22516 10008 22568
rect 11336 22559 11388 22568
rect 11336 22525 11345 22559
rect 11345 22525 11379 22559
rect 11379 22525 11388 22559
rect 11336 22516 11388 22525
rect 39396 22763 39448 22772
rect 39396 22729 39405 22763
rect 39405 22729 39439 22763
rect 39439 22729 39448 22763
rect 39396 22720 39448 22729
rect 40132 22720 40184 22772
rect 40868 22720 40920 22772
rect 43260 22720 43312 22772
rect 43996 22720 44048 22772
rect 45284 22720 45336 22772
rect 46572 22720 46624 22772
rect 46940 22720 46992 22772
rect 47032 22720 47084 22772
rect 47860 22720 47912 22772
rect 47952 22763 48004 22772
rect 47952 22729 47961 22763
rect 47961 22729 47995 22763
rect 47995 22729 48004 22763
rect 47952 22720 48004 22729
rect 48044 22720 48096 22772
rect 49792 22720 49844 22772
rect 43168 22584 43220 22636
rect 44272 22584 44324 22636
rect 39764 22559 39816 22568
rect 39764 22525 39773 22559
rect 39773 22525 39807 22559
rect 39807 22525 39816 22559
rect 39764 22516 39816 22525
rect 41236 22516 41288 22568
rect 42984 22559 43036 22568
rect 42984 22525 42993 22559
rect 42993 22525 43027 22559
rect 43027 22525 43036 22559
rect 42984 22516 43036 22525
rect 43444 22516 43496 22568
rect 3240 22423 3292 22432
rect 3240 22389 3249 22423
rect 3249 22389 3283 22423
rect 3283 22389 3292 22423
rect 3240 22380 3292 22389
rect 4620 22423 4672 22432
rect 4620 22389 4629 22423
rect 4629 22389 4663 22423
rect 4663 22389 4672 22423
rect 4620 22380 4672 22389
rect 8024 22423 8076 22432
rect 8024 22389 8033 22423
rect 8033 22389 8067 22423
rect 8067 22389 8076 22423
rect 8024 22380 8076 22389
rect 8576 22380 8628 22432
rect 9680 22423 9732 22432
rect 9680 22389 9689 22423
rect 9689 22389 9723 22423
rect 9723 22389 9732 22423
rect 9680 22380 9732 22389
rect 44824 22448 44876 22500
rect 45928 22516 45980 22568
rect 46756 22584 46808 22636
rect 49240 22652 49292 22704
rect 50804 22720 50856 22772
rect 52828 22720 52880 22772
rect 53104 22720 53156 22772
rect 53472 22720 53524 22772
rect 55312 22763 55364 22772
rect 55312 22729 55321 22763
rect 55321 22729 55355 22763
rect 55355 22729 55364 22763
rect 55312 22720 55364 22729
rect 57336 22720 57388 22772
rect 57428 22763 57480 22772
rect 57428 22729 57437 22763
rect 57437 22729 57471 22763
rect 57471 22729 57480 22763
rect 57428 22720 57480 22729
rect 57520 22720 57572 22772
rect 58164 22720 58216 22772
rect 58256 22720 58308 22772
rect 58900 22720 58952 22772
rect 10968 22380 11020 22432
rect 11888 22423 11940 22432
rect 11888 22389 11897 22423
rect 11897 22389 11931 22423
rect 11931 22389 11940 22423
rect 11888 22380 11940 22389
rect 12440 22423 12492 22432
rect 12440 22389 12449 22423
rect 12449 22389 12483 22423
rect 12483 22389 12492 22423
rect 12440 22380 12492 22389
rect 42432 22423 42484 22432
rect 42432 22389 42441 22423
rect 42441 22389 42475 22423
rect 42475 22389 42484 22423
rect 42432 22380 42484 22389
rect 43444 22423 43496 22432
rect 43444 22389 43453 22423
rect 43453 22389 43487 22423
rect 43487 22389 43496 22423
rect 43444 22380 43496 22389
rect 43812 22380 43864 22432
rect 47216 22448 47268 22500
rect 48044 22627 48096 22636
rect 48044 22593 48053 22627
rect 48053 22593 48087 22627
rect 48087 22593 48096 22627
rect 48044 22584 48096 22593
rect 54760 22584 54812 22636
rect 55312 22627 55364 22636
rect 55312 22593 55321 22627
rect 55321 22593 55355 22627
rect 55355 22593 55364 22627
rect 55312 22584 55364 22593
rect 50804 22559 50856 22568
rect 50804 22525 50813 22559
rect 50813 22525 50847 22559
rect 50847 22525 50856 22559
rect 50804 22516 50856 22525
rect 57428 22627 57480 22636
rect 57428 22593 57437 22627
rect 57437 22593 57471 22627
rect 57471 22593 57480 22627
rect 57428 22584 57480 22593
rect 58808 22584 58860 22636
rect 48872 22380 48924 22432
rect 52460 22380 52512 22432
rect 53196 22380 53248 22432
rect 56692 22380 56744 22432
rect 56968 22380 57020 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3240 22176 3292 22228
rect 3332 22219 3384 22228
rect 3332 22185 3341 22219
rect 3341 22185 3375 22219
rect 3375 22185 3384 22219
rect 3332 22176 3384 22185
rect 4804 22176 4856 22228
rect 7380 22219 7432 22228
rect 7380 22185 7389 22219
rect 7389 22185 7423 22219
rect 7423 22185 7432 22219
rect 7380 22176 7432 22185
rect 8576 22176 8628 22228
rect 2872 22108 2924 22160
rect 4068 22108 4120 22160
rect 5724 22151 5776 22160
rect 5724 22117 5733 22151
rect 5733 22117 5767 22151
rect 5767 22117 5776 22151
rect 5724 22108 5776 22117
rect 3792 21972 3844 22024
rect 5356 21972 5408 22024
rect 5632 22015 5684 22024
rect 5632 21981 5641 22015
rect 5641 21981 5675 22015
rect 5675 21981 5684 22015
rect 5632 21972 5684 21981
rect 4436 21947 4488 21956
rect 4436 21913 4470 21947
rect 4470 21913 4488 21947
rect 4436 21904 4488 21913
rect 6000 21972 6052 22024
rect 6644 21904 6696 21956
rect 9220 22176 9272 22228
rect 9956 22219 10008 22228
rect 9956 22185 9965 22219
rect 9965 22185 9999 22219
rect 9999 22185 10008 22219
rect 9956 22176 10008 22185
rect 11888 22176 11940 22228
rect 42432 22176 42484 22228
rect 42708 22176 42760 22228
rect 54760 22219 54812 22228
rect 54760 22185 54769 22219
rect 54769 22185 54803 22219
rect 54803 22185 54812 22219
rect 54760 22176 54812 22185
rect 55312 22176 55364 22228
rect 57428 22176 57480 22228
rect 10784 22108 10836 22160
rect 10968 22108 11020 22160
rect 11520 22083 11572 22092
rect 11520 22049 11529 22083
rect 11529 22049 11563 22083
rect 11563 22049 11572 22083
rect 11520 22040 11572 22049
rect 10140 22015 10192 22024
rect 10140 21981 10149 22015
rect 10149 21981 10183 22015
rect 10183 21981 10192 22015
rect 10140 21972 10192 21981
rect 10324 21972 10376 22024
rect 41328 22040 41380 22092
rect 44180 22040 44232 22092
rect 47952 22040 48004 22092
rect 48136 22040 48188 22092
rect 8208 21904 8260 21956
rect 10600 21904 10652 21956
rect 9956 21836 10008 21888
rect 42616 21972 42668 22024
rect 12440 21904 12492 21956
rect 13084 21836 13136 21888
rect 42892 21972 42944 22024
rect 44272 22015 44324 22024
rect 44272 21981 44281 22015
rect 44281 21981 44315 22015
rect 44315 21981 44324 22015
rect 44272 21972 44324 21981
rect 43168 21904 43220 21956
rect 45652 22015 45704 22024
rect 45652 21981 45661 22015
rect 45661 21981 45695 22015
rect 45695 21981 45704 22015
rect 45652 21972 45704 21981
rect 44548 21904 44600 21956
rect 47124 22015 47176 22024
rect 47124 21981 47133 22015
rect 47133 21981 47167 22015
rect 47167 21981 47176 22015
rect 47124 21972 47176 21981
rect 50160 22040 50212 22092
rect 49332 22015 49384 22024
rect 49332 21981 49341 22015
rect 49341 21981 49375 22015
rect 49375 21981 49384 22015
rect 49332 21972 49384 21981
rect 48688 21904 48740 21956
rect 49148 21904 49200 21956
rect 43536 21879 43588 21888
rect 43536 21845 43545 21879
rect 43545 21845 43579 21879
rect 43579 21845 43588 21879
rect 43536 21836 43588 21845
rect 43996 21836 44048 21888
rect 44732 21836 44784 21888
rect 46204 21836 46256 21888
rect 49240 21879 49292 21888
rect 49240 21845 49249 21879
rect 49249 21845 49283 21879
rect 49283 21845 49292 21879
rect 49240 21836 49292 21845
rect 54300 22108 54352 22160
rect 51172 22015 51224 22024
rect 51172 21981 51181 22015
rect 51181 21981 51215 22015
rect 51215 21981 51224 22015
rect 51172 21972 51224 21981
rect 52460 22015 52512 22024
rect 52460 21981 52469 22015
rect 52469 21981 52503 22015
rect 52503 21981 52512 22015
rect 52460 21972 52512 21981
rect 53564 22015 53616 22024
rect 53564 21981 53573 22015
rect 53573 21981 53607 22015
rect 53607 21981 53616 22015
rect 53564 21972 53616 21981
rect 54024 21972 54076 22024
rect 54116 22015 54168 22024
rect 54116 21981 54125 22015
rect 54125 21981 54159 22015
rect 54159 21981 54168 22015
rect 54116 21972 54168 21981
rect 52184 21904 52236 21956
rect 54484 22040 54536 22092
rect 55128 22108 55180 22160
rect 57612 22151 57664 22160
rect 57612 22117 57621 22151
rect 57621 22117 57655 22151
rect 57655 22117 57664 22151
rect 57612 22108 57664 22117
rect 57428 22083 57480 22092
rect 57428 22049 57437 22083
rect 57437 22049 57471 22083
rect 57471 22049 57480 22083
rect 57428 22040 57480 22049
rect 52368 21836 52420 21888
rect 52736 21879 52788 21888
rect 52736 21845 52745 21879
rect 52745 21845 52779 21879
rect 52779 21845 52788 21879
rect 52736 21836 52788 21845
rect 53932 21836 53984 21888
rect 54208 21836 54260 21888
rect 54484 21947 54536 21956
rect 54484 21913 54493 21947
rect 54493 21913 54527 21947
rect 54527 21913 54536 21947
rect 54484 21904 54536 21913
rect 54944 22015 54996 22024
rect 54944 21981 54953 22015
rect 54953 21981 54987 22015
rect 54987 21981 54996 22015
rect 54944 21972 54996 21981
rect 55220 21904 55272 21956
rect 55956 22015 56008 22024
rect 55956 21981 55965 22015
rect 55965 21981 55999 22015
rect 55999 21981 56008 22015
rect 55956 21972 56008 21981
rect 56876 22015 56928 22024
rect 56876 21981 56885 22015
rect 56885 21981 56919 22015
rect 56919 21981 56928 22015
rect 56876 21972 56928 21981
rect 56784 21947 56836 21956
rect 56784 21913 56793 21947
rect 56793 21913 56827 21947
rect 56827 21913 56836 21947
rect 56784 21904 56836 21913
rect 57152 22015 57204 22024
rect 57152 21981 57161 22015
rect 57161 21981 57195 22015
rect 57195 21981 57204 22015
rect 57152 21972 57204 21981
rect 57060 21904 57112 21956
rect 57888 21947 57940 21956
rect 57888 21913 57897 21947
rect 57897 21913 57931 21947
rect 57931 21913 57940 21947
rect 57888 21904 57940 21913
rect 57980 21836 58032 21888
rect 58072 21836 58124 21888
rect 58256 21879 58308 21888
rect 58256 21845 58265 21879
rect 58265 21845 58299 21879
rect 58299 21845 58308 21879
rect 58256 21836 58308 21845
rect 58348 21879 58400 21888
rect 58348 21845 58357 21879
rect 58357 21845 58391 21879
rect 58391 21845 58400 21879
rect 58348 21836 58400 21845
rect 58900 21904 58952 21956
rect 58716 21836 58768 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 3792 21632 3844 21684
rect 5724 21564 5776 21616
rect 6644 21632 6696 21684
rect 7012 21675 7064 21684
rect 7012 21641 7021 21675
rect 7021 21641 7055 21675
rect 7055 21641 7064 21675
rect 7012 21632 7064 21641
rect 8208 21632 8260 21684
rect 42892 21632 42944 21684
rect 42984 21632 43036 21684
rect 43168 21632 43220 21684
rect 2688 21539 2740 21548
rect 2688 21505 2697 21539
rect 2697 21505 2731 21539
rect 2731 21505 2740 21539
rect 2688 21496 2740 21505
rect 4712 21539 4764 21548
rect 4712 21505 4721 21539
rect 4721 21505 4755 21539
rect 4755 21505 4764 21539
rect 4712 21496 4764 21505
rect 4804 21539 4856 21548
rect 4804 21505 4813 21539
rect 4813 21505 4847 21539
rect 4847 21505 4856 21539
rect 4804 21496 4856 21505
rect 940 21428 992 21480
rect 3700 21471 3752 21480
rect 3700 21437 3709 21471
rect 3709 21437 3743 21471
rect 3743 21437 3752 21471
rect 3700 21428 3752 21437
rect 4436 21428 4488 21480
rect 6000 21539 6052 21548
rect 6000 21505 6009 21539
rect 6009 21505 6043 21539
rect 6043 21505 6052 21539
rect 6000 21496 6052 21505
rect 6460 21539 6512 21548
rect 6460 21505 6469 21539
rect 6469 21505 6503 21539
rect 6503 21505 6512 21539
rect 6460 21496 6512 21505
rect 7564 21564 7616 21616
rect 7012 21496 7064 21548
rect 8208 21539 8260 21548
rect 8208 21505 8217 21539
rect 8217 21505 8251 21539
rect 8251 21505 8260 21539
rect 8208 21496 8260 21505
rect 43536 21632 43588 21684
rect 44180 21632 44232 21684
rect 45468 21632 45520 21684
rect 10692 21471 10744 21480
rect 10692 21437 10701 21471
rect 10701 21437 10735 21471
rect 10735 21437 10744 21471
rect 10692 21428 10744 21437
rect 8116 21360 8168 21412
rect 9864 21360 9916 21412
rect 11980 21360 12032 21412
rect 19984 21360 20036 21412
rect 34520 21360 34572 21412
rect 44548 21607 44600 21616
rect 44548 21573 44557 21607
rect 44557 21573 44591 21607
rect 44591 21573 44600 21607
rect 44548 21564 44600 21573
rect 44732 21564 44784 21616
rect 46204 21564 46256 21616
rect 43996 21496 44048 21548
rect 44088 21496 44140 21548
rect 44364 21539 44416 21548
rect 44364 21505 44373 21539
rect 44373 21505 44407 21539
rect 44407 21505 44416 21539
rect 44364 21496 44416 21505
rect 46664 21675 46716 21684
rect 46664 21641 46673 21675
rect 46673 21641 46707 21675
rect 46707 21641 46716 21675
rect 46664 21632 46716 21641
rect 49424 21632 49476 21684
rect 49424 21539 49476 21548
rect 49424 21505 49433 21539
rect 49433 21505 49467 21539
rect 49467 21505 49476 21539
rect 49424 21496 49476 21505
rect 49516 21539 49568 21548
rect 49516 21505 49525 21539
rect 49525 21505 49559 21539
rect 49559 21505 49568 21539
rect 49516 21496 49568 21505
rect 52184 21632 52236 21684
rect 49884 21539 49936 21548
rect 49884 21505 49893 21539
rect 49893 21505 49927 21539
rect 49927 21505 49936 21539
rect 49884 21496 49936 21505
rect 44732 21360 44784 21412
rect 48780 21428 48832 21480
rect 50160 21539 50212 21548
rect 50160 21505 50169 21539
rect 50169 21505 50203 21539
rect 50203 21505 50212 21539
rect 50160 21496 50212 21505
rect 49608 21360 49660 21412
rect 3056 21292 3108 21344
rect 10048 21335 10100 21344
rect 10048 21301 10057 21335
rect 10057 21301 10091 21335
rect 10091 21301 10100 21335
rect 10048 21292 10100 21301
rect 12164 21335 12216 21344
rect 12164 21301 12173 21335
rect 12173 21301 12207 21335
rect 12207 21301 12216 21335
rect 12164 21292 12216 21301
rect 42892 21335 42944 21344
rect 42892 21301 42901 21335
rect 42901 21301 42935 21335
rect 42935 21301 42944 21335
rect 42892 21292 42944 21301
rect 43812 21335 43864 21344
rect 43812 21301 43821 21335
rect 43821 21301 43855 21335
rect 43855 21301 43864 21335
rect 43812 21292 43864 21301
rect 44640 21335 44692 21344
rect 44640 21301 44649 21335
rect 44649 21301 44683 21335
rect 44683 21301 44692 21335
rect 44640 21292 44692 21301
rect 47768 21335 47820 21344
rect 47768 21301 47777 21335
rect 47777 21301 47811 21335
rect 47811 21301 47820 21335
rect 47768 21292 47820 21301
rect 49700 21335 49752 21344
rect 49700 21301 49709 21335
rect 49709 21301 49743 21335
rect 49743 21301 49752 21335
rect 49700 21292 49752 21301
rect 50528 21539 50580 21548
rect 50528 21505 50537 21539
rect 50537 21505 50571 21539
rect 50571 21505 50580 21539
rect 50528 21496 50580 21505
rect 51080 21564 51132 21616
rect 50988 21539 51040 21548
rect 50988 21505 50997 21539
rect 50997 21505 51031 21539
rect 51031 21505 51040 21539
rect 50988 21496 51040 21505
rect 52736 21632 52788 21684
rect 54116 21675 54168 21684
rect 54116 21641 54125 21675
rect 54125 21641 54159 21675
rect 54159 21641 54168 21675
rect 54116 21632 54168 21641
rect 54484 21632 54536 21684
rect 55956 21632 56008 21684
rect 56784 21632 56836 21684
rect 57888 21632 57940 21684
rect 58072 21632 58124 21684
rect 51448 21360 51500 21412
rect 53564 21496 53616 21548
rect 54760 21539 54812 21548
rect 54760 21505 54794 21539
rect 54794 21505 54812 21539
rect 54760 21496 54812 21505
rect 56416 21428 56468 21480
rect 57888 21471 57940 21480
rect 57888 21437 57897 21471
rect 57897 21437 57931 21471
rect 57931 21437 57940 21471
rect 57888 21428 57940 21437
rect 55220 21292 55272 21344
rect 55404 21292 55456 21344
rect 56600 21292 56652 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 3056 21088 3108 21140
rect 3700 21088 3752 21140
rect 4712 21088 4764 21140
rect 6460 21088 6512 21140
rect 8116 21088 8168 21140
rect 9864 21088 9916 21140
rect 9956 21088 10008 21140
rect 10048 21088 10100 21140
rect 10416 21088 10468 21140
rect 12164 21088 12216 21140
rect 42892 21088 42944 21140
rect 44364 21088 44416 21140
rect 44732 21131 44784 21140
rect 44732 21097 44741 21131
rect 44741 21097 44775 21131
rect 44775 21097 44784 21131
rect 44732 21088 44784 21097
rect 45652 21088 45704 21140
rect 47768 21088 47820 21140
rect 49424 21088 49476 21140
rect 49608 21088 49660 21140
rect 49700 21088 49752 21140
rect 50528 21088 50580 21140
rect 50988 21088 51040 21140
rect 54576 21088 54628 21140
rect 54760 21088 54812 21140
rect 3148 20927 3200 20936
rect 3148 20893 3157 20927
rect 3157 20893 3191 20927
rect 3191 20893 3200 20927
rect 3148 20884 3200 20893
rect 2412 20816 2464 20868
rect 2872 20816 2924 20868
rect 3516 20927 3568 20936
rect 3516 20893 3525 20927
rect 3525 20893 3559 20927
rect 3559 20893 3568 20927
rect 3516 20884 3568 20893
rect 4344 20927 4396 20936
rect 4344 20893 4353 20927
rect 4353 20893 4387 20927
rect 4387 20893 4396 20927
rect 4344 20884 4396 20893
rect 5356 20884 5408 20936
rect 4620 20816 4672 20868
rect 9956 20884 10008 20936
rect 11980 20952 12032 21004
rect 13728 20927 13780 20936
rect 13728 20893 13737 20927
rect 13737 20893 13771 20927
rect 13771 20893 13780 20927
rect 13728 20884 13780 20893
rect 18236 20884 18288 20936
rect 43444 20927 43496 20936
rect 43444 20893 43453 20927
rect 43453 20893 43487 20927
rect 43487 20893 43496 20927
rect 43444 20884 43496 20893
rect 43996 20952 44048 21004
rect 44640 20884 44692 20936
rect 45468 20952 45520 21004
rect 2688 20748 2740 20800
rect 6920 20816 6972 20868
rect 8024 20816 8076 20868
rect 8576 20816 8628 20868
rect 8852 20816 8904 20868
rect 9772 20816 9824 20868
rect 10048 20748 10100 20800
rect 10140 20791 10192 20800
rect 10140 20757 10149 20791
rect 10149 20757 10183 20791
rect 10183 20757 10192 20791
rect 10140 20748 10192 20757
rect 10968 20816 11020 20868
rect 44088 20816 44140 20868
rect 47032 20884 47084 20936
rect 49056 21020 49108 21072
rect 47952 20952 48004 21004
rect 47124 20748 47176 20800
rect 48320 20884 48372 20936
rect 48412 20816 48464 20868
rect 48504 20791 48556 20800
rect 48504 20757 48513 20791
rect 48513 20757 48547 20791
rect 48547 20757 48556 20791
rect 48504 20748 48556 20757
rect 50068 20952 50120 21004
rect 49976 20884 50028 20936
rect 55404 20952 55456 21004
rect 56600 21088 56652 21140
rect 57428 21088 57480 21140
rect 57888 21088 57940 21140
rect 50988 20884 51040 20936
rect 51448 20927 51500 20936
rect 51448 20893 51457 20927
rect 51457 20893 51491 20927
rect 51491 20893 51500 20927
rect 51448 20884 51500 20893
rect 52276 20884 52328 20936
rect 55864 20884 55916 20936
rect 55956 20927 56008 20936
rect 55956 20893 55965 20927
rect 55965 20893 55999 20927
rect 55999 20893 56008 20927
rect 55956 20884 56008 20893
rect 50712 20816 50764 20868
rect 55128 20748 55180 20800
rect 56416 20927 56468 20936
rect 56416 20893 56425 20927
rect 56425 20893 56459 20927
rect 56459 20893 56468 20927
rect 56416 20884 56468 20893
rect 57980 20927 58032 20936
rect 57980 20893 57989 20927
rect 57989 20893 58023 20927
rect 58023 20893 58032 20927
rect 57980 20884 58032 20893
rect 58348 20884 58400 20936
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 4344 20544 4396 20596
rect 6460 20544 6512 20596
rect 6920 20544 6972 20596
rect 8116 20587 8168 20596
rect 8116 20553 8125 20587
rect 8125 20553 8159 20587
rect 8159 20553 8168 20587
rect 8116 20544 8168 20553
rect 8208 20544 8260 20596
rect 10692 20544 10744 20596
rect 13176 20587 13228 20596
rect 13176 20553 13185 20587
rect 13185 20553 13219 20587
rect 13219 20553 13228 20587
rect 13176 20544 13228 20553
rect 19984 20544 20036 20596
rect 48228 20544 48280 20596
rect 48504 20544 48556 20596
rect 48780 20587 48832 20596
rect 48780 20553 48789 20587
rect 48789 20553 48823 20587
rect 48823 20553 48832 20587
rect 48780 20544 48832 20553
rect 49148 20544 49200 20596
rect 49332 20544 49384 20596
rect 49700 20544 49752 20596
rect 50620 20544 50672 20596
rect 51448 20544 51500 20596
rect 55864 20544 55916 20596
rect 55956 20544 56008 20596
rect 2688 20451 2740 20460
rect 2688 20417 2697 20451
rect 2697 20417 2731 20451
rect 2731 20417 2740 20451
rect 2688 20408 2740 20417
rect 3976 20451 4028 20460
rect 3976 20417 3985 20451
rect 3985 20417 4019 20451
rect 4019 20417 4028 20451
rect 3976 20408 4028 20417
rect 5080 20408 5132 20460
rect 5908 20408 5960 20460
rect 4620 20340 4672 20392
rect 3884 20272 3936 20324
rect 8300 20451 8352 20460
rect 8300 20417 8309 20451
rect 8309 20417 8343 20451
rect 8343 20417 8352 20451
rect 8300 20408 8352 20417
rect 8576 20476 8628 20528
rect 11244 20476 11296 20528
rect 18236 20451 18288 20460
rect 18236 20417 18245 20451
rect 18245 20417 18279 20451
rect 18279 20417 18288 20451
rect 48412 20476 48464 20528
rect 18236 20408 18288 20417
rect 10140 20383 10192 20392
rect 10140 20349 10149 20383
rect 10149 20349 10183 20383
rect 10183 20349 10192 20383
rect 10140 20340 10192 20349
rect 10324 20340 10376 20392
rect 10968 20340 11020 20392
rect 10600 20272 10652 20324
rect 4620 20204 4672 20256
rect 5816 20204 5868 20256
rect 6276 20204 6328 20256
rect 6736 20204 6788 20256
rect 7932 20247 7984 20256
rect 7932 20213 7941 20247
rect 7941 20213 7975 20247
rect 7975 20213 7984 20247
rect 7932 20204 7984 20213
rect 8024 20204 8076 20256
rect 9036 20204 9088 20256
rect 31116 20204 31168 20256
rect 45744 20204 45796 20256
rect 48504 20451 48556 20460
rect 48504 20417 48513 20451
rect 48513 20417 48547 20451
rect 48547 20417 48556 20451
rect 48504 20408 48556 20417
rect 48596 20451 48648 20460
rect 48596 20417 48605 20451
rect 48605 20417 48639 20451
rect 48639 20417 48648 20451
rect 48596 20408 48648 20417
rect 53012 20519 53064 20528
rect 53012 20485 53021 20519
rect 53021 20485 53055 20519
rect 53055 20485 53064 20519
rect 53012 20476 53064 20485
rect 57152 20476 57204 20528
rect 49056 20340 49108 20392
rect 49424 20340 49476 20392
rect 52828 20408 52880 20460
rect 48320 20247 48372 20256
rect 48320 20213 48329 20247
rect 48329 20213 48363 20247
rect 48363 20213 48372 20247
rect 48320 20204 48372 20213
rect 51816 20204 51868 20256
rect 52920 20204 52972 20256
rect 54300 20204 54352 20256
rect 56324 20408 56376 20460
rect 56692 20340 56744 20392
rect 57796 20204 57848 20256
rect 58532 20204 58584 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3884 20000 3936 20052
rect 4160 20000 4212 20052
rect 5080 20000 5132 20052
rect 5816 20000 5868 20052
rect 7104 20000 7156 20052
rect 5908 19975 5960 19984
rect 5908 19941 5917 19975
rect 5917 19941 5951 19975
rect 5951 19941 5960 19975
rect 5908 19932 5960 19941
rect 940 19728 992 19780
rect 1400 19660 1452 19712
rect 4068 19839 4120 19848
rect 4068 19805 4077 19839
rect 4077 19805 4111 19839
rect 4111 19805 4120 19839
rect 4068 19796 4120 19805
rect 4160 19796 4212 19848
rect 4620 19864 4672 19916
rect 4528 19839 4580 19848
rect 4528 19805 4537 19839
rect 4537 19805 4571 19839
rect 4571 19805 4580 19839
rect 4528 19796 4580 19805
rect 6276 19864 6328 19916
rect 10048 20000 10100 20052
rect 48320 20000 48372 20052
rect 48504 20000 48556 20052
rect 51080 20000 51132 20052
rect 51264 20000 51316 20052
rect 51816 20043 51868 20052
rect 51816 20009 51825 20043
rect 51825 20009 51859 20043
rect 51859 20009 51868 20043
rect 51816 20000 51868 20009
rect 52368 20000 52420 20052
rect 47032 19907 47084 19916
rect 47032 19873 47041 19907
rect 47041 19873 47075 19907
rect 47075 19873 47084 19907
rect 47032 19864 47084 19873
rect 6736 19796 6788 19848
rect 7932 19796 7984 19848
rect 9312 19796 9364 19848
rect 11428 19839 11480 19848
rect 11428 19805 11437 19839
rect 11437 19805 11471 19839
rect 11471 19805 11480 19839
rect 11428 19796 11480 19805
rect 3516 19703 3568 19712
rect 3516 19669 3525 19703
rect 3525 19669 3559 19703
rect 3559 19669 3568 19703
rect 3516 19660 3568 19669
rect 3792 19703 3844 19712
rect 3792 19669 3801 19703
rect 3801 19669 3835 19703
rect 3835 19669 3844 19703
rect 3792 19660 3844 19669
rect 4620 19660 4672 19712
rect 4712 19660 4764 19712
rect 8300 19728 8352 19780
rect 10968 19728 11020 19780
rect 41788 19796 41840 19848
rect 48596 19839 48648 19848
rect 48596 19805 48605 19839
rect 48605 19805 48639 19839
rect 48639 19805 48648 19839
rect 48596 19796 48648 19805
rect 49424 19864 49476 19916
rect 49608 19839 49660 19848
rect 49608 19805 49617 19839
rect 49617 19805 49651 19839
rect 49651 19805 49660 19839
rect 49608 19796 49660 19805
rect 49792 19839 49844 19848
rect 49792 19805 49801 19839
rect 49801 19805 49835 19839
rect 49835 19805 49844 19839
rect 49792 19796 49844 19805
rect 10876 19703 10928 19712
rect 10876 19669 10885 19703
rect 10885 19669 10919 19703
rect 10919 19669 10928 19703
rect 10876 19660 10928 19669
rect 11796 19660 11848 19712
rect 45744 19660 45796 19712
rect 47216 19660 47268 19712
rect 48412 19660 48464 19712
rect 49516 19660 49568 19712
rect 50344 19839 50396 19848
rect 50344 19805 50353 19839
rect 50353 19805 50387 19839
rect 50387 19805 50396 19839
rect 50344 19796 50396 19805
rect 50436 19839 50488 19848
rect 50436 19805 50445 19839
rect 50445 19805 50479 19839
rect 50479 19805 50488 19839
rect 50436 19796 50488 19805
rect 50896 19932 50948 19984
rect 51356 19796 51408 19848
rect 51816 19796 51868 19848
rect 51172 19660 51224 19712
rect 51632 19660 51684 19712
rect 53472 19660 53524 19712
rect 55220 20000 55272 20052
rect 56692 20043 56744 20052
rect 56692 20009 56701 20043
rect 56701 20009 56735 20043
rect 56735 20009 56744 20043
rect 56692 20000 56744 20009
rect 53656 19771 53708 19780
rect 53656 19737 53665 19771
rect 53665 19737 53699 19771
rect 53699 19737 53708 19771
rect 53656 19728 53708 19737
rect 54024 19839 54076 19848
rect 54024 19805 54033 19839
rect 54033 19805 54067 19839
rect 54067 19805 54076 19839
rect 54024 19796 54076 19805
rect 54208 19796 54260 19848
rect 54300 19839 54352 19848
rect 54300 19805 54309 19839
rect 54309 19805 54343 19839
rect 54343 19805 54352 19839
rect 54300 19796 54352 19805
rect 55036 19728 55088 19780
rect 55312 19839 55364 19848
rect 55312 19805 55321 19839
rect 55321 19805 55355 19839
rect 55355 19805 55364 19839
rect 55312 19796 55364 19805
rect 56416 19796 56468 19848
rect 58256 19839 58308 19848
rect 58256 19805 58265 19839
rect 58265 19805 58299 19839
rect 58299 19805 58308 19839
rect 58256 19796 58308 19805
rect 55220 19728 55272 19780
rect 57060 19771 57112 19780
rect 57060 19737 57094 19771
rect 57094 19737 57112 19771
rect 57060 19728 57112 19737
rect 55680 19660 55732 19712
rect 56324 19660 56376 19712
rect 57336 19660 57388 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 1400 19499 1452 19508
rect 1400 19465 1409 19499
rect 1409 19465 1443 19499
rect 1443 19465 1452 19499
rect 1400 19456 1452 19465
rect 8852 19499 8904 19508
rect 8852 19465 8861 19499
rect 8861 19465 8895 19499
rect 8895 19465 8904 19499
rect 8852 19456 8904 19465
rect 2412 19388 2464 19440
rect 5356 19388 5408 19440
rect 10324 19388 10376 19440
rect 10876 19456 10928 19508
rect 11980 19456 12032 19508
rect 47216 19456 47268 19508
rect 3148 19363 3200 19372
rect 3148 19329 3157 19363
rect 3157 19329 3191 19363
rect 3191 19329 3200 19363
rect 3148 19320 3200 19329
rect 3516 19320 3568 19372
rect 2872 19295 2924 19304
rect 2872 19261 2881 19295
rect 2881 19261 2915 19295
rect 2915 19261 2924 19295
rect 2872 19252 2924 19261
rect 6828 19252 6880 19304
rect 9312 19320 9364 19372
rect 10968 19363 11020 19372
rect 10968 19329 10977 19363
rect 10977 19329 11011 19363
rect 11011 19329 11020 19363
rect 10968 19320 11020 19329
rect 11244 19320 11296 19372
rect 47952 19456 48004 19508
rect 49148 19456 49200 19508
rect 49332 19499 49384 19508
rect 49332 19465 49341 19499
rect 49341 19465 49375 19499
rect 49375 19465 49384 19499
rect 49332 19456 49384 19465
rect 50620 19456 50672 19508
rect 51356 19456 51408 19508
rect 53656 19456 53708 19508
rect 55220 19456 55272 19508
rect 57060 19456 57112 19508
rect 42616 19252 42668 19304
rect 47216 19184 47268 19236
rect 49056 19252 49108 19304
rect 49700 19363 49752 19372
rect 49700 19329 49709 19363
rect 49709 19329 49743 19363
rect 49743 19329 49752 19363
rect 49700 19320 49752 19329
rect 49884 19363 49936 19372
rect 49884 19329 49893 19363
rect 49893 19329 49927 19363
rect 49927 19329 49936 19363
rect 49884 19320 49936 19329
rect 50160 19320 50212 19372
rect 56600 19388 56652 19440
rect 57612 19456 57664 19508
rect 58348 19456 58400 19508
rect 50988 19320 51040 19372
rect 49792 19252 49844 19304
rect 50896 19252 50948 19304
rect 51172 19252 51224 19304
rect 51632 19363 51684 19372
rect 51632 19329 51641 19363
rect 51641 19329 51675 19363
rect 51675 19329 51684 19363
rect 51632 19320 51684 19329
rect 51724 19363 51776 19372
rect 51724 19329 51733 19363
rect 51733 19329 51767 19363
rect 51767 19329 51776 19363
rect 51724 19320 51776 19329
rect 51908 19363 51960 19372
rect 51908 19329 51917 19363
rect 51917 19329 51951 19363
rect 51951 19329 51960 19363
rect 51908 19320 51960 19329
rect 53656 19320 53708 19372
rect 54208 19320 54260 19372
rect 55680 19320 55732 19372
rect 56140 19320 56192 19372
rect 53840 19252 53892 19304
rect 55128 19252 55180 19304
rect 57060 19252 57112 19304
rect 3240 19159 3292 19168
rect 3240 19125 3249 19159
rect 3249 19125 3283 19159
rect 3283 19125 3292 19159
rect 3240 19116 3292 19125
rect 4068 19116 4120 19168
rect 8392 19116 8444 19168
rect 11060 19159 11112 19168
rect 11060 19125 11069 19159
rect 11069 19125 11103 19159
rect 11103 19125 11112 19159
rect 11060 19116 11112 19125
rect 47400 19116 47452 19168
rect 48320 19159 48372 19168
rect 48320 19125 48329 19159
rect 48329 19125 48363 19159
rect 48363 19125 48372 19159
rect 48320 19116 48372 19125
rect 57336 19363 57388 19372
rect 57336 19329 57345 19363
rect 57345 19329 57379 19363
rect 57379 19329 57388 19363
rect 57336 19320 57388 19329
rect 57796 19320 57848 19372
rect 57428 19252 57480 19304
rect 57612 19184 57664 19236
rect 52276 19116 52328 19168
rect 54852 19159 54904 19168
rect 54852 19125 54861 19159
rect 54861 19125 54895 19159
rect 54895 19125 54904 19159
rect 54852 19116 54904 19125
rect 55036 19116 55088 19168
rect 57336 19116 57388 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 2872 18912 2924 18964
rect 3792 18912 3844 18964
rect 4804 18912 4856 18964
rect 4712 18844 4764 18896
rect 3240 18776 3292 18828
rect 2228 18751 2280 18760
rect 2228 18717 2237 18751
rect 2237 18717 2271 18751
rect 2271 18717 2280 18751
rect 2228 18708 2280 18717
rect 3608 18751 3660 18760
rect 3608 18717 3617 18751
rect 3617 18717 3651 18751
rect 3651 18717 3660 18751
rect 3608 18708 3660 18717
rect 4068 18708 4120 18760
rect 4896 18776 4948 18828
rect 6828 18912 6880 18964
rect 11428 18912 11480 18964
rect 49884 18912 49936 18964
rect 51724 18955 51776 18964
rect 51724 18921 51733 18955
rect 51733 18921 51767 18955
rect 51767 18921 51776 18955
rect 51724 18912 51776 18921
rect 51908 18912 51960 18964
rect 9956 18844 10008 18896
rect 6828 18819 6880 18828
rect 6828 18785 6837 18819
rect 6837 18785 6871 18819
rect 6871 18785 6880 18819
rect 6828 18776 6880 18785
rect 8392 18776 8444 18828
rect 9772 18776 9824 18828
rect 11060 18819 11112 18828
rect 11060 18785 11069 18819
rect 11069 18785 11103 18819
rect 11103 18785 11112 18819
rect 11060 18776 11112 18785
rect 47032 18819 47084 18828
rect 47032 18785 47041 18819
rect 47041 18785 47075 18819
rect 47075 18785 47084 18819
rect 47032 18776 47084 18785
rect 6368 18708 6420 18760
rect 6644 18751 6696 18760
rect 6644 18717 6653 18751
rect 6653 18717 6687 18751
rect 6687 18717 6696 18751
rect 6644 18708 6696 18717
rect 3792 18615 3844 18624
rect 3792 18581 3801 18615
rect 3801 18581 3835 18615
rect 3835 18581 3844 18615
rect 3792 18572 3844 18581
rect 4528 18572 4580 18624
rect 5908 18615 5960 18624
rect 5908 18581 5917 18615
rect 5917 18581 5951 18615
rect 5951 18581 5960 18615
rect 5908 18572 5960 18581
rect 7012 18615 7064 18624
rect 7012 18581 7021 18615
rect 7021 18581 7055 18615
rect 7055 18581 7064 18615
rect 7012 18572 7064 18581
rect 12072 18640 12124 18692
rect 46940 18640 46992 18692
rect 47400 18708 47452 18760
rect 48320 18708 48372 18760
rect 48412 18708 48464 18760
rect 49424 18776 49476 18828
rect 49516 18776 49568 18828
rect 50988 18844 51040 18896
rect 52276 18819 52328 18828
rect 49792 18751 49844 18760
rect 49792 18717 49801 18751
rect 49801 18717 49835 18751
rect 49835 18717 49844 18751
rect 49792 18708 49844 18717
rect 52276 18785 52285 18819
rect 52285 18785 52319 18819
rect 52319 18785 52328 18819
rect 52276 18776 52328 18785
rect 53840 18844 53892 18896
rect 49332 18640 49384 18692
rect 50620 18751 50672 18760
rect 50620 18717 50629 18751
rect 50629 18717 50663 18751
rect 50663 18717 50672 18751
rect 50620 18708 50672 18717
rect 51264 18708 51316 18760
rect 51632 18708 51684 18760
rect 51724 18751 51776 18760
rect 51724 18717 51733 18751
rect 51733 18717 51767 18751
rect 51767 18717 51776 18751
rect 51724 18708 51776 18717
rect 8300 18572 8352 18624
rect 10324 18572 10376 18624
rect 45652 18615 45704 18624
rect 45652 18581 45661 18615
rect 45661 18581 45695 18615
rect 45695 18581 45704 18615
rect 45652 18572 45704 18581
rect 47308 18615 47360 18624
rect 47308 18581 47317 18615
rect 47317 18581 47351 18615
rect 47351 18581 47360 18615
rect 47308 18572 47360 18581
rect 49148 18615 49200 18624
rect 49148 18581 49157 18615
rect 49157 18581 49191 18615
rect 49191 18581 49200 18615
rect 49148 18572 49200 18581
rect 49884 18572 49936 18624
rect 51540 18572 51592 18624
rect 52276 18572 52328 18624
rect 54760 18751 54812 18760
rect 54760 18717 54769 18751
rect 54769 18717 54803 18751
rect 54803 18717 54812 18751
rect 54760 18708 54812 18717
rect 56784 18844 56836 18896
rect 57612 18955 57664 18964
rect 57612 18921 57621 18955
rect 57621 18921 57655 18955
rect 57655 18921 57664 18955
rect 57612 18912 57664 18921
rect 58348 18955 58400 18964
rect 58348 18921 58357 18955
rect 58357 18921 58391 18955
rect 58391 18921 58400 18955
rect 58348 18912 58400 18921
rect 55404 18708 55456 18760
rect 56324 18708 56376 18760
rect 53932 18615 53984 18624
rect 53932 18581 53941 18615
rect 53941 18581 53975 18615
rect 53975 18581 53984 18615
rect 53932 18572 53984 18581
rect 58164 18844 58216 18896
rect 57336 18776 57388 18828
rect 57796 18708 57848 18760
rect 58072 18751 58124 18760
rect 58072 18717 58081 18751
rect 58081 18717 58115 18751
rect 58115 18717 58124 18751
rect 58072 18708 58124 18717
rect 58348 18708 58400 18760
rect 58900 18708 58952 18760
rect 57888 18572 57940 18624
rect 57980 18615 58032 18624
rect 57980 18581 57989 18615
rect 57989 18581 58023 18615
rect 58023 18581 58032 18615
rect 57980 18572 58032 18581
rect 58072 18572 58124 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 3608 18368 3660 18420
rect 6828 18368 6880 18420
rect 46940 18368 46992 18420
rect 47216 18411 47268 18420
rect 47216 18377 47225 18411
rect 47225 18377 47259 18411
rect 47259 18377 47268 18411
rect 47216 18368 47268 18377
rect 47676 18368 47728 18420
rect 48596 18368 48648 18420
rect 49148 18368 49200 18420
rect 49332 18411 49384 18420
rect 49332 18377 49341 18411
rect 49341 18377 49375 18411
rect 49375 18377 49384 18411
rect 49332 18368 49384 18377
rect 49884 18368 49936 18420
rect 51724 18368 51776 18420
rect 52276 18368 52328 18420
rect 53656 18368 53708 18420
rect 2504 18300 2556 18352
rect 4528 18300 4580 18352
rect 5448 18300 5500 18352
rect 2688 18275 2740 18284
rect 2688 18241 2697 18275
rect 2697 18241 2731 18275
rect 2731 18241 2740 18275
rect 2688 18232 2740 18241
rect 1584 18207 1636 18216
rect 1584 18173 1593 18207
rect 1593 18173 1627 18207
rect 1627 18173 1636 18207
rect 1584 18164 1636 18173
rect 3516 18207 3568 18216
rect 3516 18173 3525 18207
rect 3525 18173 3559 18207
rect 3559 18173 3568 18207
rect 3516 18164 3568 18173
rect 5908 18207 5960 18216
rect 5908 18173 5917 18207
rect 5917 18173 5951 18207
rect 5951 18173 5960 18207
rect 5908 18164 5960 18173
rect 6276 18164 6328 18216
rect 7012 18300 7064 18352
rect 6920 18275 6972 18284
rect 6920 18241 6929 18275
rect 6929 18241 6963 18275
rect 6963 18241 6972 18275
rect 6920 18232 6972 18241
rect 8300 18300 8352 18352
rect 9680 18232 9732 18284
rect 11060 18164 11112 18216
rect 9956 18096 10008 18148
rect 2872 18028 2924 18080
rect 4712 18028 4764 18080
rect 9220 18071 9272 18080
rect 9220 18037 9229 18071
rect 9229 18037 9263 18071
rect 9263 18037 9272 18071
rect 9220 18028 9272 18037
rect 12164 18071 12216 18080
rect 12164 18037 12173 18071
rect 12173 18037 12207 18071
rect 12207 18037 12216 18071
rect 12164 18028 12216 18037
rect 38660 18028 38712 18080
rect 45652 18028 45704 18080
rect 47308 18232 47360 18284
rect 49608 18300 49660 18352
rect 48872 18232 48924 18284
rect 53932 18368 53984 18420
rect 51540 18275 51592 18284
rect 51540 18241 51549 18275
rect 51549 18241 51583 18275
rect 51583 18241 51592 18275
rect 51540 18232 51592 18241
rect 51724 18275 51776 18284
rect 51724 18241 51733 18275
rect 51733 18241 51767 18275
rect 51767 18241 51776 18275
rect 51724 18232 51776 18241
rect 51816 18275 51868 18284
rect 51816 18241 51825 18275
rect 51825 18241 51859 18275
rect 51859 18241 51868 18275
rect 51816 18232 51868 18241
rect 53840 18300 53892 18352
rect 51540 18096 51592 18148
rect 53564 18232 53616 18284
rect 53656 18275 53708 18284
rect 53656 18241 53665 18275
rect 53665 18241 53699 18275
rect 53699 18241 53708 18275
rect 53656 18232 53708 18241
rect 53840 18164 53892 18216
rect 54760 18368 54812 18420
rect 56600 18368 56652 18420
rect 56968 18232 57020 18284
rect 57980 18368 58032 18420
rect 58072 18368 58124 18420
rect 58348 18411 58400 18420
rect 58348 18377 58357 18411
rect 58357 18377 58391 18411
rect 58391 18377 58400 18411
rect 58348 18368 58400 18377
rect 58900 18368 58952 18420
rect 57796 18164 57848 18216
rect 53564 18096 53616 18148
rect 57612 18096 57664 18148
rect 49792 18028 49844 18080
rect 50988 18028 51040 18080
rect 51356 18071 51408 18080
rect 51356 18037 51365 18071
rect 51365 18037 51399 18071
rect 51399 18037 51408 18071
rect 51356 18028 51408 18037
rect 53748 18028 53800 18080
rect 55220 18028 55272 18080
rect 58348 18028 58400 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 2688 17824 2740 17876
rect 3516 17824 3568 17876
rect 3792 17824 3844 17876
rect 4620 17824 4672 17876
rect 4896 17824 4948 17876
rect 2872 17731 2924 17740
rect 2872 17697 2881 17731
rect 2881 17697 2915 17731
rect 2915 17697 2924 17731
rect 2872 17688 2924 17697
rect 3148 17663 3200 17672
rect 3148 17629 3157 17663
rect 3157 17629 3191 17663
rect 3191 17629 3200 17663
rect 3148 17620 3200 17629
rect 4712 17756 4764 17808
rect 2412 17552 2464 17604
rect 2228 17484 2280 17536
rect 4068 17620 4120 17672
rect 6920 17620 6972 17672
rect 9864 17824 9916 17876
rect 11980 17824 12032 17876
rect 48320 17824 48372 17876
rect 49608 17824 49660 17876
rect 50068 17824 50120 17876
rect 53564 17824 53616 17876
rect 53840 17824 53892 17876
rect 54852 17824 54904 17876
rect 55220 17824 55272 17876
rect 57888 17824 57940 17876
rect 57980 17824 58032 17876
rect 58256 17867 58308 17876
rect 58256 17833 58265 17867
rect 58265 17833 58299 17867
rect 58299 17833 58308 17867
rect 58256 17824 58308 17833
rect 8668 17731 8720 17740
rect 8668 17697 8677 17731
rect 8677 17697 8711 17731
rect 8711 17697 8720 17731
rect 8668 17688 8720 17697
rect 6644 17552 6696 17604
rect 9036 17595 9088 17604
rect 9036 17561 9045 17595
rect 9045 17561 9079 17595
rect 9079 17561 9088 17595
rect 9036 17552 9088 17561
rect 9956 17620 10008 17672
rect 10324 17620 10376 17672
rect 47860 17663 47912 17672
rect 47860 17629 47869 17663
rect 47869 17629 47903 17663
rect 47903 17629 47912 17663
rect 47860 17620 47912 17629
rect 12164 17552 12216 17604
rect 49240 17620 49292 17672
rect 51356 17620 51408 17672
rect 49608 17552 49660 17604
rect 53380 17552 53432 17604
rect 53748 17620 53800 17672
rect 53932 17663 53984 17672
rect 53932 17629 53941 17663
rect 53941 17629 53975 17663
rect 53975 17629 53984 17663
rect 53932 17620 53984 17629
rect 55128 17731 55180 17740
rect 55128 17697 55137 17731
rect 55137 17697 55171 17731
rect 55171 17697 55180 17731
rect 55128 17688 55180 17697
rect 55312 17663 55364 17672
rect 55312 17629 55321 17663
rect 55321 17629 55355 17663
rect 55355 17629 55364 17663
rect 55312 17620 55364 17629
rect 9220 17484 9272 17536
rect 10048 17527 10100 17536
rect 10048 17493 10057 17527
rect 10057 17493 10091 17527
rect 10091 17493 10100 17527
rect 10048 17484 10100 17493
rect 10232 17527 10284 17536
rect 10232 17493 10241 17527
rect 10241 17493 10275 17527
rect 10275 17493 10284 17527
rect 10232 17484 10284 17493
rect 47308 17527 47360 17536
rect 47308 17493 47317 17527
rect 47317 17493 47351 17527
rect 47351 17493 47360 17527
rect 47308 17484 47360 17493
rect 49148 17484 49200 17536
rect 49240 17527 49292 17536
rect 49240 17493 49249 17527
rect 49249 17493 49283 17527
rect 49283 17493 49292 17527
rect 49240 17484 49292 17493
rect 52736 17484 52788 17536
rect 56508 17484 56560 17536
rect 57612 17620 57664 17672
rect 58072 17665 58124 17672
rect 58072 17631 58090 17665
rect 58090 17631 58124 17665
rect 57704 17595 57756 17604
rect 57704 17561 57713 17595
rect 57713 17561 57747 17595
rect 57747 17561 57756 17595
rect 57704 17552 57756 17561
rect 58072 17620 58124 17631
rect 58256 17620 58308 17672
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 2228 17144 2280 17196
rect 4160 17119 4212 17128
rect 4160 17085 4169 17119
rect 4169 17085 4203 17119
rect 4203 17085 4212 17119
rect 4160 17076 4212 17085
rect 5540 17280 5592 17332
rect 6184 17280 6236 17332
rect 8668 17280 8720 17332
rect 11060 17323 11112 17332
rect 11060 17289 11069 17323
rect 11069 17289 11103 17323
rect 11103 17289 11112 17323
rect 11060 17280 11112 17289
rect 11244 17280 11296 17332
rect 47308 17280 47360 17332
rect 47860 17280 47912 17332
rect 48688 17280 48740 17332
rect 6460 17187 6512 17196
rect 6460 17153 6469 17187
rect 6469 17153 6503 17187
rect 6503 17153 6512 17187
rect 6460 17144 6512 17153
rect 6644 17144 6696 17196
rect 6920 17212 6972 17264
rect 6184 17119 6236 17128
rect 6184 17085 6193 17119
rect 6193 17085 6227 17119
rect 6227 17085 6236 17119
rect 6184 17076 6236 17085
rect 8116 17119 8168 17128
rect 8116 17085 8125 17119
rect 8125 17085 8159 17119
rect 8159 17085 8168 17119
rect 8116 17076 8168 17085
rect 9036 17076 9088 17128
rect 10232 17119 10284 17128
rect 10232 17085 10241 17119
rect 10241 17085 10275 17119
rect 10275 17085 10284 17119
rect 10232 17076 10284 17085
rect 48044 17212 48096 17264
rect 49240 17280 49292 17332
rect 55128 17280 55180 17332
rect 56968 17280 57020 17332
rect 57704 17280 57756 17332
rect 57980 17280 58032 17332
rect 58256 17280 58308 17332
rect 48780 17187 48832 17196
rect 48780 17153 48789 17187
rect 48789 17153 48823 17187
rect 48823 17153 48832 17187
rect 48780 17144 48832 17153
rect 55404 17212 55456 17264
rect 49332 17187 49384 17196
rect 49332 17153 49341 17187
rect 49341 17153 49375 17187
rect 49375 17153 49384 17187
rect 49332 17144 49384 17153
rect 47676 17076 47728 17128
rect 48044 17119 48096 17128
rect 48044 17085 48053 17119
rect 48053 17085 48087 17119
rect 48087 17085 48096 17119
rect 48044 17076 48096 17085
rect 3424 16983 3476 16992
rect 3424 16949 3433 16983
rect 3433 16949 3467 16983
rect 3467 16949 3476 16983
rect 3424 16940 3476 16949
rect 48780 17008 48832 17060
rect 56508 17187 56560 17196
rect 56508 17153 56517 17187
rect 56517 17153 56551 17187
rect 56551 17153 56560 17187
rect 56508 17144 56560 17153
rect 57336 17144 57388 17196
rect 57612 17187 57664 17196
rect 57612 17153 57621 17187
rect 57621 17153 57655 17187
rect 57655 17153 57664 17187
rect 57612 17144 57664 17153
rect 4804 16940 4856 16992
rect 5448 16983 5500 16992
rect 5448 16949 5457 16983
rect 5457 16949 5491 16983
rect 5491 16949 5500 16983
rect 5448 16940 5500 16949
rect 7472 16983 7524 16992
rect 7472 16949 7481 16983
rect 7481 16949 7515 16983
rect 7515 16949 7524 16983
rect 7472 16940 7524 16949
rect 46940 16940 46992 16992
rect 47124 16983 47176 16992
rect 47124 16949 47133 16983
rect 47133 16949 47167 16983
rect 47167 16949 47176 16983
rect 47124 16940 47176 16949
rect 58348 17144 58400 17196
rect 58164 17008 58216 17060
rect 58900 17008 58952 17060
rect 49240 16940 49292 16992
rect 49332 16940 49384 16992
rect 52736 16940 52788 16992
rect 57980 16940 58032 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3424 16736 3476 16788
rect 5448 16736 5500 16788
rect 6184 16736 6236 16788
rect 7472 16736 7524 16788
rect 10048 16736 10100 16788
rect 3148 16600 3200 16652
rect 6276 16600 6328 16652
rect 9772 16600 9824 16652
rect 45928 16600 45980 16652
rect 47032 16736 47084 16788
rect 48044 16779 48096 16788
rect 48044 16745 48053 16779
rect 48053 16745 48087 16779
rect 48087 16745 48096 16779
rect 48044 16736 48096 16745
rect 48688 16736 48740 16788
rect 49240 16736 49292 16788
rect 49424 16736 49476 16788
rect 3792 16575 3844 16584
rect 3792 16541 3801 16575
rect 3801 16541 3835 16575
rect 3835 16541 3844 16575
rect 3792 16532 3844 16541
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 4068 16532 4120 16584
rect 1676 16439 1728 16448
rect 1676 16405 1685 16439
rect 1685 16405 1719 16439
rect 1719 16405 1728 16439
rect 1676 16396 1728 16405
rect 2412 16396 2464 16448
rect 4528 16396 4580 16448
rect 5356 16464 5408 16516
rect 6368 16575 6420 16584
rect 6368 16541 6377 16575
rect 6377 16541 6411 16575
rect 6411 16541 6420 16575
rect 6368 16532 6420 16541
rect 6920 16532 6972 16584
rect 46940 16575 46992 16584
rect 46940 16541 46974 16575
rect 46974 16541 46992 16575
rect 46940 16532 46992 16541
rect 47676 16532 47728 16584
rect 49976 16643 50028 16652
rect 49976 16609 49985 16643
rect 49985 16609 50019 16643
rect 50019 16609 50028 16643
rect 49976 16600 50028 16609
rect 50896 16736 50948 16788
rect 52828 16736 52880 16788
rect 52920 16779 52972 16788
rect 52920 16745 52929 16779
rect 52929 16745 52963 16779
rect 52963 16745 52972 16779
rect 52920 16736 52972 16745
rect 53472 16736 53524 16788
rect 57796 16779 57848 16788
rect 57796 16745 57805 16779
rect 57805 16745 57839 16779
rect 57839 16745 57848 16779
rect 57796 16736 57848 16745
rect 57980 16779 58032 16788
rect 57980 16745 57989 16779
rect 57989 16745 58023 16779
rect 58023 16745 58032 16779
rect 57980 16736 58032 16745
rect 53564 16668 53616 16720
rect 52736 16600 52788 16652
rect 6736 16439 6788 16448
rect 6736 16405 6745 16439
rect 6745 16405 6779 16439
rect 6779 16405 6788 16439
rect 6736 16396 6788 16405
rect 9036 16439 9088 16448
rect 9036 16405 9045 16439
rect 9045 16405 9079 16439
rect 9079 16405 9088 16439
rect 9036 16396 9088 16405
rect 10324 16396 10376 16448
rect 51172 16532 51224 16584
rect 51816 16464 51868 16516
rect 51264 16396 51316 16448
rect 52920 16507 52972 16516
rect 52920 16473 52929 16507
rect 52929 16473 52963 16507
rect 52963 16473 52972 16507
rect 52920 16464 52972 16473
rect 53196 16575 53248 16584
rect 53196 16541 53205 16575
rect 53205 16541 53239 16575
rect 53239 16541 53248 16575
rect 53196 16532 53248 16541
rect 53288 16575 53340 16584
rect 53288 16541 53297 16575
rect 53297 16541 53331 16575
rect 53331 16541 53340 16575
rect 53288 16532 53340 16541
rect 53564 16532 53616 16584
rect 56876 16668 56928 16720
rect 55588 16575 55640 16584
rect 55588 16541 55597 16575
rect 55597 16541 55631 16575
rect 55631 16541 55640 16575
rect 55588 16532 55640 16541
rect 56600 16575 56652 16584
rect 56600 16541 56609 16575
rect 56609 16541 56643 16575
rect 56643 16541 56652 16575
rect 56600 16532 56652 16541
rect 58164 16575 58216 16584
rect 58164 16541 58173 16575
rect 58173 16541 58207 16575
rect 58207 16541 58216 16575
rect 58164 16532 58216 16541
rect 52552 16396 52604 16448
rect 52828 16439 52880 16448
rect 52828 16405 52837 16439
rect 52837 16405 52871 16439
rect 52871 16405 52880 16439
rect 52828 16396 52880 16405
rect 53656 16396 53708 16448
rect 56876 16464 56928 16516
rect 54116 16396 54168 16448
rect 55496 16439 55548 16448
rect 55496 16405 55505 16439
rect 55505 16405 55539 16439
rect 55539 16405 55548 16439
rect 55496 16396 55548 16405
rect 56784 16396 56836 16448
rect 57980 16396 58032 16448
rect 58900 16396 58952 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 3792 16192 3844 16244
rect 6368 16235 6420 16244
rect 6368 16201 6377 16235
rect 6377 16201 6411 16235
rect 6411 16201 6420 16235
rect 6368 16192 6420 16201
rect 6920 16192 6972 16244
rect 8116 16192 8168 16244
rect 940 16056 992 16108
rect 4712 16056 4764 16108
rect 6736 16056 6788 16108
rect 48320 16124 48372 16176
rect 1676 15988 1728 16040
rect 4620 15988 4672 16040
rect 45928 16099 45980 16108
rect 45928 16065 45937 16099
rect 45937 16065 45971 16099
rect 45971 16065 45980 16099
rect 45928 16056 45980 16065
rect 47676 16056 47728 16108
rect 48044 16099 48096 16108
rect 48044 16065 48053 16099
rect 48053 16065 48087 16099
rect 48087 16065 48096 16099
rect 48044 16056 48096 16065
rect 48412 16099 48464 16108
rect 48412 16065 48421 16099
rect 48421 16065 48455 16099
rect 48455 16065 48464 16099
rect 48412 16056 48464 16065
rect 48688 16056 48740 16108
rect 44824 15988 44876 16040
rect 48504 15988 48556 16040
rect 49240 16192 49292 16244
rect 49976 16192 50028 16244
rect 52828 16192 52880 16244
rect 53288 16192 53340 16244
rect 53564 16235 53616 16244
rect 53564 16201 53573 16235
rect 53573 16201 53607 16235
rect 53607 16201 53616 16235
rect 53564 16192 53616 16201
rect 54116 16235 54168 16244
rect 54116 16201 54125 16235
rect 54125 16201 54159 16235
rect 54159 16201 54168 16235
rect 54116 16192 54168 16201
rect 49608 16124 49660 16176
rect 48320 15920 48372 15972
rect 51080 16099 51132 16108
rect 51080 16065 51089 16099
rect 51089 16065 51123 16099
rect 51123 16065 51132 16099
rect 51080 16056 51132 16065
rect 51264 16099 51316 16108
rect 51264 16065 51273 16099
rect 51273 16065 51307 16099
rect 51307 16065 51316 16099
rect 51264 16056 51316 16065
rect 53380 16124 53432 16176
rect 53656 16124 53708 16176
rect 55588 16192 55640 16244
rect 56600 16192 56652 16244
rect 57336 16192 57388 16244
rect 49424 15920 49476 15972
rect 2688 15852 2740 15904
rect 47952 15895 48004 15904
rect 47952 15861 47961 15895
rect 47961 15861 47995 15895
rect 47995 15861 48004 15895
rect 47952 15852 48004 15861
rect 49516 15852 49568 15904
rect 51816 15852 51868 15904
rect 52552 15988 52604 16040
rect 56784 16124 56836 16176
rect 56876 16124 56928 16176
rect 55404 16099 55456 16108
rect 55404 16065 55438 16099
rect 55438 16065 55456 16099
rect 53380 15920 53432 15972
rect 54024 15920 54076 15972
rect 55404 16056 55456 16065
rect 53104 15852 53156 15904
rect 57152 16031 57204 16040
rect 57152 15997 57161 16031
rect 57161 15997 57195 16031
rect 57195 15997 57204 16031
rect 57152 15988 57204 15997
rect 57796 16056 57848 16108
rect 58532 16124 58584 16176
rect 57704 15988 57756 16040
rect 58348 16099 58400 16108
rect 58348 16065 58357 16099
rect 58357 16065 58391 16099
rect 58391 16065 58400 16099
rect 58348 16056 58400 16065
rect 57888 15920 57940 15972
rect 55312 15852 55364 15904
rect 56600 15895 56652 15904
rect 56600 15861 56609 15895
rect 56609 15861 56643 15895
rect 56643 15861 56652 15895
rect 56600 15852 56652 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 47952 15648 48004 15700
rect 49884 15648 49936 15700
rect 50712 15648 50764 15700
rect 51632 15648 51684 15700
rect 52920 15648 52972 15700
rect 53472 15691 53524 15700
rect 53472 15657 53481 15691
rect 53481 15657 53515 15691
rect 53515 15657 53524 15691
rect 53472 15648 53524 15657
rect 53932 15648 53984 15700
rect 55404 15648 55456 15700
rect 56600 15648 56652 15700
rect 57152 15648 57204 15700
rect 57704 15648 57756 15700
rect 57980 15691 58032 15700
rect 57980 15657 57989 15691
rect 57989 15657 58023 15691
rect 58023 15657 58032 15691
rect 57980 15648 58032 15657
rect 58164 15648 58216 15700
rect 45928 15512 45980 15564
rect 49240 15580 49292 15632
rect 46572 15376 46624 15428
rect 48504 15376 48556 15428
rect 49240 15487 49292 15496
rect 49240 15453 49249 15487
rect 49249 15453 49283 15487
rect 49283 15453 49292 15487
rect 49240 15444 49292 15453
rect 49332 15487 49384 15496
rect 49332 15453 49341 15487
rect 49341 15453 49375 15487
rect 49375 15453 49384 15487
rect 49332 15444 49384 15453
rect 49424 15444 49476 15496
rect 50068 15444 50120 15496
rect 51816 15512 51868 15564
rect 49976 15376 50028 15428
rect 50804 15444 50856 15496
rect 51632 15487 51684 15496
rect 51632 15453 51641 15487
rect 51641 15453 51675 15487
rect 51675 15453 51684 15487
rect 51632 15444 51684 15453
rect 52736 15580 52788 15632
rect 51080 15376 51132 15428
rect 52828 15444 52880 15496
rect 53104 15580 53156 15632
rect 56508 15580 56560 15632
rect 54852 15512 54904 15564
rect 53472 15444 53524 15496
rect 53564 15487 53616 15496
rect 53564 15453 53573 15487
rect 53573 15453 53607 15487
rect 53607 15453 53616 15487
rect 53564 15444 53616 15453
rect 47492 15351 47544 15360
rect 47492 15317 47501 15351
rect 47501 15317 47535 15351
rect 47535 15317 47544 15351
rect 47492 15308 47544 15317
rect 47584 15308 47636 15360
rect 48044 15308 48096 15360
rect 49516 15308 49568 15360
rect 54024 15376 54076 15428
rect 55496 15512 55548 15564
rect 56784 15580 56836 15632
rect 56876 15580 56928 15632
rect 57796 15580 57848 15632
rect 57704 15487 57756 15496
rect 57704 15453 57713 15487
rect 57713 15453 57747 15487
rect 57747 15453 57756 15487
rect 57704 15444 57756 15453
rect 58072 15487 58124 15496
rect 58072 15453 58081 15487
rect 58081 15453 58115 15487
rect 58115 15453 58124 15487
rect 58072 15444 58124 15453
rect 58440 15376 58492 15428
rect 56324 15308 56376 15360
rect 56968 15308 57020 15360
rect 57520 15308 57572 15360
rect 57704 15308 57756 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 46572 15147 46624 15156
rect 46572 15113 46581 15147
rect 46581 15113 46615 15147
rect 46615 15113 46624 15147
rect 46572 15104 46624 15113
rect 48412 15104 48464 15156
rect 49056 15104 49108 15156
rect 49240 15147 49292 15156
rect 49240 15113 49249 15147
rect 49249 15113 49283 15147
rect 49283 15113 49292 15147
rect 49240 15104 49292 15113
rect 50068 15104 50120 15156
rect 50160 15104 50212 15156
rect 50620 15104 50672 15156
rect 10140 14968 10192 15020
rect 47584 15011 47636 15020
rect 47584 14977 47593 15011
rect 47593 14977 47627 15011
rect 47627 14977 47636 15011
rect 47584 14968 47636 14977
rect 47952 14968 48004 15020
rect 48136 15011 48188 15020
rect 48136 14977 48145 15011
rect 48145 14977 48179 15011
rect 48179 14977 48188 15011
rect 48136 14968 48188 14977
rect 48504 15011 48556 15020
rect 48504 14977 48513 15011
rect 48513 14977 48547 15011
rect 48547 14977 48556 15011
rect 48504 14968 48556 14977
rect 48688 15011 48740 15020
rect 48688 14977 48697 15011
rect 48697 14977 48731 15011
rect 48731 14977 48740 15011
rect 48688 14968 48740 14977
rect 48780 15011 48832 15020
rect 48780 14977 48789 15011
rect 48789 14977 48823 15011
rect 48823 14977 48832 15011
rect 48780 14968 48832 14977
rect 50436 15036 50488 15088
rect 50068 14968 50120 15020
rect 940 14900 992 14952
rect 47492 14900 47544 14952
rect 50528 14968 50580 15020
rect 50712 15011 50764 15020
rect 50712 14977 50721 15011
rect 50721 14977 50755 15011
rect 50755 14977 50764 15011
rect 50712 14968 50764 14977
rect 51080 15147 51132 15156
rect 51080 15113 51089 15147
rect 51089 15113 51123 15147
rect 51123 15113 51132 15147
rect 51080 15104 51132 15113
rect 51632 15104 51684 15156
rect 52828 15147 52880 15156
rect 52828 15113 52837 15147
rect 52837 15113 52871 15147
rect 52871 15113 52880 15147
rect 52828 15104 52880 15113
rect 53012 15104 53064 15156
rect 53196 15147 53248 15156
rect 53196 15113 53205 15147
rect 53205 15113 53239 15147
rect 53239 15113 53248 15147
rect 53196 15104 53248 15113
rect 53564 15147 53616 15156
rect 53564 15113 53573 15147
rect 53573 15113 53607 15147
rect 53607 15113 53616 15147
rect 53564 15104 53616 15113
rect 53656 15104 53708 15156
rect 54024 15147 54076 15156
rect 54024 15113 54033 15147
rect 54033 15113 54067 15147
rect 54067 15113 54076 15147
rect 54024 15104 54076 15113
rect 56968 15104 57020 15156
rect 57704 15147 57756 15156
rect 57704 15113 57713 15147
rect 57713 15113 57747 15147
rect 57747 15113 57756 15147
rect 57704 15104 57756 15113
rect 47124 14832 47176 14884
rect 51448 15011 51500 15020
rect 51448 14977 51457 15011
rect 51457 14977 51491 15011
rect 51491 14977 51500 15011
rect 51448 14968 51500 14977
rect 52736 15011 52788 15020
rect 52736 14977 52745 15011
rect 52745 14977 52779 15011
rect 52779 14977 52788 15011
rect 52736 14968 52788 14977
rect 52920 15011 52972 15020
rect 52920 14977 52929 15011
rect 52929 14977 52963 15011
rect 52963 14977 52972 15011
rect 52920 14968 52972 14977
rect 53380 15036 53432 15088
rect 53932 14968 53984 15020
rect 54116 15079 54168 15088
rect 54116 15045 54125 15079
rect 54125 15045 54159 15079
rect 54159 15045 54168 15079
rect 54116 15036 54168 15045
rect 55588 14968 55640 15020
rect 58440 15011 58492 15020
rect 58440 14977 58449 15011
rect 58449 14977 58483 15011
rect 58483 14977 58492 15011
rect 58440 14968 58492 14977
rect 53840 14900 53892 14952
rect 56140 14943 56192 14952
rect 56140 14909 56149 14943
rect 56149 14909 56183 14943
rect 56183 14909 56192 14943
rect 56140 14900 56192 14909
rect 57152 14943 57204 14952
rect 57152 14909 57161 14943
rect 57161 14909 57195 14943
rect 57195 14909 57204 14943
rect 57152 14900 57204 14909
rect 54024 14832 54076 14884
rect 50528 14764 50580 14816
rect 55496 14807 55548 14816
rect 55496 14773 55505 14807
rect 55505 14773 55539 14807
rect 55539 14773 55548 14807
rect 55496 14764 55548 14773
rect 57888 14807 57940 14816
rect 57888 14773 57897 14807
rect 57897 14773 57931 14807
rect 57931 14773 57940 14807
rect 57888 14764 57940 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 48504 14560 48556 14612
rect 48688 14560 48740 14612
rect 49148 14560 49200 14612
rect 50528 14603 50580 14612
rect 50528 14569 50537 14603
rect 50537 14569 50571 14603
rect 50571 14569 50580 14603
rect 50528 14560 50580 14569
rect 50620 14560 50672 14612
rect 50712 14560 50764 14612
rect 52736 14560 52788 14612
rect 57152 14560 57204 14612
rect 58900 14560 58952 14612
rect 56692 14535 56744 14544
rect 56692 14501 56701 14535
rect 56701 14501 56735 14535
rect 56735 14501 56744 14535
rect 56692 14492 56744 14501
rect 58072 14492 58124 14544
rect 49332 14399 49384 14408
rect 49332 14365 49341 14399
rect 49341 14365 49375 14399
rect 49375 14365 49384 14399
rect 49332 14356 49384 14365
rect 50436 14399 50488 14408
rect 50436 14365 50445 14399
rect 50445 14365 50479 14399
rect 50479 14365 50488 14399
rect 50436 14356 50488 14365
rect 52276 14399 52328 14408
rect 52276 14365 52285 14399
rect 52285 14365 52319 14399
rect 52319 14365 52328 14399
rect 52276 14356 52328 14365
rect 53380 14356 53432 14408
rect 53932 14356 53984 14408
rect 48504 14220 48556 14272
rect 52092 14220 52144 14272
rect 54024 14220 54076 14272
rect 54760 14220 54812 14272
rect 55036 14263 55088 14272
rect 55036 14229 55045 14263
rect 55045 14229 55079 14263
rect 55079 14229 55088 14263
rect 55036 14220 55088 14229
rect 55312 14399 55364 14408
rect 55312 14365 55321 14399
rect 55321 14365 55355 14399
rect 55355 14365 55364 14399
rect 55312 14356 55364 14365
rect 55220 14288 55272 14340
rect 56784 14288 56836 14340
rect 58164 14220 58216 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 48320 14016 48372 14068
rect 49332 14059 49384 14068
rect 49332 14025 49341 14059
rect 49341 14025 49375 14059
rect 49375 14025 49384 14059
rect 49332 14016 49384 14025
rect 51448 14059 51500 14068
rect 51448 14025 51457 14059
rect 51457 14025 51491 14059
rect 51491 14025 51500 14059
rect 51448 14016 51500 14025
rect 52920 14016 52972 14068
rect 53012 14016 53064 14068
rect 53656 14016 53708 14068
rect 53840 14016 53892 14068
rect 55036 14016 55088 14068
rect 55220 14016 55272 14068
rect 55496 14016 55548 14068
rect 55588 14016 55640 14068
rect 56140 14016 56192 14068
rect 56692 14016 56744 14068
rect 56784 14059 56836 14068
rect 56784 14025 56793 14059
rect 56793 14025 56827 14059
rect 56827 14025 56836 14059
rect 56784 14016 56836 14025
rect 58072 14016 58124 14068
rect 58164 14016 58216 14068
rect 58900 14016 58952 14068
rect 47124 13880 47176 13932
rect 47584 13923 47636 13932
rect 47584 13889 47593 13923
rect 47593 13889 47627 13923
rect 47627 13889 47636 13923
rect 47584 13880 47636 13889
rect 47952 13923 48004 13932
rect 47952 13889 47961 13923
rect 47961 13889 47995 13923
rect 47995 13889 48004 13923
rect 47952 13880 48004 13889
rect 49884 13880 49936 13932
rect 48504 13812 48556 13864
rect 49240 13812 49292 13864
rect 49332 13855 49384 13864
rect 49332 13821 49341 13855
rect 49341 13821 49375 13855
rect 49375 13821 49384 13855
rect 49332 13812 49384 13821
rect 49148 13787 49200 13796
rect 49148 13753 49157 13787
rect 49157 13753 49191 13787
rect 49191 13753 49200 13787
rect 49148 13744 49200 13753
rect 51264 13923 51316 13932
rect 51264 13889 51273 13923
rect 51273 13889 51307 13923
rect 51307 13889 51316 13923
rect 51264 13880 51316 13889
rect 51448 13880 51500 13932
rect 51540 13923 51592 13932
rect 51540 13889 51549 13923
rect 51549 13889 51583 13923
rect 51583 13889 51592 13923
rect 51540 13880 51592 13889
rect 51816 13923 51868 13932
rect 51816 13889 51825 13923
rect 51825 13889 51859 13923
rect 51859 13889 51868 13923
rect 51816 13880 51868 13889
rect 53104 13923 53156 13932
rect 53104 13889 53113 13923
rect 53113 13889 53147 13923
rect 53147 13889 53156 13923
rect 53104 13880 53156 13889
rect 52920 13812 52972 13864
rect 53932 13880 53984 13932
rect 54024 13923 54076 13932
rect 54024 13889 54033 13923
rect 54033 13889 54067 13923
rect 54067 13889 54076 13923
rect 54024 13880 54076 13889
rect 54760 13744 54812 13796
rect 53840 13676 53892 13728
rect 54852 13676 54904 13728
rect 56324 13812 56376 13864
rect 57888 13812 57940 13864
rect 57980 13744 58032 13796
rect 56600 13719 56652 13728
rect 56600 13685 56609 13719
rect 56609 13685 56643 13719
rect 56643 13685 56652 13719
rect 56600 13676 56652 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 47584 13472 47636 13524
rect 47952 13472 48004 13524
rect 49332 13472 49384 13524
rect 51540 13472 51592 13524
rect 53840 13515 53892 13524
rect 53840 13481 53849 13515
rect 53849 13481 53883 13515
rect 53883 13481 53892 13515
rect 53840 13472 53892 13481
rect 54024 13472 54076 13524
rect 54852 13472 54904 13524
rect 56600 13472 56652 13524
rect 58348 13515 58400 13524
rect 45928 13336 45980 13388
rect 46296 13379 46348 13388
rect 46296 13345 46305 13379
rect 46305 13345 46339 13379
rect 46339 13345 46348 13379
rect 46296 13336 46348 13345
rect 49976 13404 50028 13456
rect 56048 13404 56100 13456
rect 6736 13268 6788 13320
rect 48320 13311 48372 13320
rect 48320 13277 48329 13311
rect 48329 13277 48363 13311
rect 48363 13277 48372 13311
rect 48320 13268 48372 13277
rect 49148 13268 49200 13320
rect 940 13200 992 13252
rect 46848 13200 46900 13252
rect 51448 13311 51500 13320
rect 51448 13277 51457 13311
rect 51457 13277 51491 13311
rect 51491 13277 51500 13311
rect 51448 13268 51500 13277
rect 56600 13379 56652 13388
rect 56600 13345 56609 13379
rect 56609 13345 56643 13379
rect 56643 13345 56652 13379
rect 56600 13336 56652 13345
rect 52092 13311 52144 13320
rect 52092 13277 52101 13311
rect 52101 13277 52135 13311
rect 52135 13277 52144 13311
rect 52092 13268 52144 13277
rect 52184 13311 52236 13320
rect 52184 13277 52193 13311
rect 52193 13277 52227 13311
rect 52227 13277 52236 13311
rect 52184 13268 52236 13277
rect 53380 13268 53432 13320
rect 53564 13311 53616 13320
rect 53564 13277 53573 13311
rect 53573 13277 53607 13311
rect 53607 13277 53616 13311
rect 53564 13268 53616 13277
rect 53932 13311 53984 13320
rect 53932 13277 53941 13311
rect 53941 13277 53975 13311
rect 53975 13277 53984 13311
rect 53932 13268 53984 13277
rect 55956 13268 56008 13320
rect 58348 13481 58357 13515
rect 58357 13481 58391 13515
rect 58391 13481 58400 13515
rect 58348 13472 58400 13481
rect 47768 13175 47820 13184
rect 47768 13141 47777 13175
rect 47777 13141 47811 13175
rect 47811 13141 47820 13175
rect 47768 13132 47820 13141
rect 49976 13132 50028 13184
rect 50712 13132 50764 13184
rect 50896 13175 50948 13184
rect 50896 13141 50905 13175
rect 50905 13141 50939 13175
rect 50939 13141 50948 13175
rect 50896 13132 50948 13141
rect 52644 13132 52696 13184
rect 52920 13175 52972 13184
rect 52920 13141 52929 13175
rect 52929 13141 52963 13175
rect 52963 13141 52972 13175
rect 52920 13132 52972 13141
rect 54208 13200 54260 13252
rect 58900 13268 58952 13320
rect 56508 13132 56560 13184
rect 56692 13132 56744 13184
rect 58716 13132 58768 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 46848 12971 46900 12980
rect 46848 12937 46857 12971
rect 46857 12937 46891 12971
rect 46891 12937 46900 12971
rect 46848 12928 46900 12937
rect 47768 12928 47820 12980
rect 48320 12928 48372 12980
rect 49976 12971 50028 12980
rect 49976 12937 49985 12971
rect 49985 12937 50019 12971
rect 50019 12937 50028 12971
rect 49976 12928 50028 12937
rect 50896 12928 50948 12980
rect 51448 12928 51500 12980
rect 51816 12928 51868 12980
rect 52276 12928 52328 12980
rect 53564 12928 53616 12980
rect 54208 12928 54260 12980
rect 47032 12835 47084 12844
rect 47032 12801 47041 12835
rect 47041 12801 47075 12835
rect 47075 12801 47084 12835
rect 47032 12792 47084 12801
rect 47124 12835 47176 12844
rect 47124 12801 47133 12835
rect 47133 12801 47167 12835
rect 47167 12801 47176 12835
rect 47124 12792 47176 12801
rect 47676 12792 47728 12844
rect 47952 12825 48004 12844
rect 47952 12792 47961 12825
rect 47961 12792 47995 12825
rect 47995 12792 48004 12825
rect 50620 12903 50672 12912
rect 50620 12869 50629 12903
rect 50629 12869 50663 12903
rect 50663 12869 50672 12903
rect 50620 12860 50672 12869
rect 50068 12835 50120 12844
rect 50068 12801 50077 12835
rect 50077 12801 50111 12835
rect 50111 12801 50120 12835
rect 50068 12792 50120 12801
rect 50712 12792 50764 12844
rect 49700 12767 49752 12776
rect 49700 12733 49709 12767
rect 49709 12733 49743 12767
rect 49743 12733 49752 12767
rect 49700 12724 49752 12733
rect 51632 12860 51684 12912
rect 51172 12792 51224 12844
rect 55312 12860 55364 12912
rect 56508 12903 56560 12912
rect 53840 12792 53892 12844
rect 53932 12792 53984 12844
rect 54760 12835 54812 12844
rect 54760 12801 54769 12835
rect 54769 12801 54803 12835
rect 54803 12801 54812 12835
rect 54760 12792 54812 12801
rect 56508 12869 56531 12903
rect 56531 12869 56560 12903
rect 56508 12860 56560 12869
rect 58532 12971 58584 12980
rect 58532 12937 58541 12971
rect 58541 12937 58575 12971
rect 58575 12937 58584 12971
rect 58532 12928 58584 12937
rect 58072 12792 58124 12844
rect 51540 12767 51592 12776
rect 51540 12733 51549 12767
rect 51549 12733 51583 12767
rect 51583 12733 51592 12767
rect 51540 12724 51592 12733
rect 48504 12631 48556 12640
rect 48504 12597 48513 12631
rect 48513 12597 48547 12631
rect 48547 12597 48556 12631
rect 48504 12588 48556 12597
rect 51080 12656 51132 12708
rect 52644 12724 52696 12776
rect 52736 12767 52788 12776
rect 52736 12733 52745 12767
rect 52745 12733 52779 12767
rect 52779 12733 52788 12767
rect 52736 12724 52788 12733
rect 56140 12724 56192 12776
rect 54852 12656 54904 12708
rect 58348 12656 58400 12708
rect 54392 12631 54444 12640
rect 54392 12597 54401 12631
rect 54401 12597 54435 12631
rect 54435 12597 54444 12631
rect 54392 12588 54444 12597
rect 54484 12588 54536 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 49700 12384 49752 12436
rect 51540 12384 51592 12436
rect 52092 12427 52144 12436
rect 52092 12393 52101 12427
rect 52101 12393 52135 12427
rect 52135 12393 52144 12427
rect 52092 12384 52144 12393
rect 55956 12427 56008 12436
rect 55956 12393 55965 12427
rect 55965 12393 55999 12427
rect 55999 12393 56008 12427
rect 55956 12384 56008 12393
rect 56140 12427 56192 12436
rect 56140 12393 56149 12427
rect 56149 12393 56183 12427
rect 56183 12393 56192 12427
rect 56140 12384 56192 12393
rect 56600 12384 56652 12436
rect 46388 12248 46440 12300
rect 48504 12223 48556 12232
rect 48504 12189 48538 12223
rect 48538 12189 48556 12223
rect 48504 12180 48556 12189
rect 49608 12087 49660 12096
rect 49608 12053 49617 12087
rect 49617 12053 49651 12087
rect 49651 12053 49660 12087
rect 49608 12044 49660 12053
rect 49884 12223 49936 12232
rect 49884 12189 49893 12223
rect 49893 12189 49927 12223
rect 49927 12189 49936 12223
rect 49884 12180 49936 12189
rect 50988 12180 51040 12232
rect 52736 12248 52788 12300
rect 52092 12180 52144 12232
rect 52920 12180 52972 12232
rect 53840 12180 53892 12232
rect 54392 12180 54444 12232
rect 56048 12316 56100 12368
rect 50528 12155 50580 12164
rect 50528 12121 50562 12155
rect 50562 12121 50580 12155
rect 50528 12112 50580 12121
rect 51632 12044 51684 12096
rect 52092 12044 52144 12096
rect 56324 12180 56376 12232
rect 57980 12112 58032 12164
rect 58256 12180 58308 12232
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 49608 11840 49660 11892
rect 49884 11840 49936 11892
rect 2688 11747 2740 11756
rect 2688 11713 2697 11747
rect 2697 11713 2731 11747
rect 2731 11713 2740 11747
rect 2688 11704 2740 11713
rect 940 11636 992 11688
rect 52368 11636 52420 11688
rect 58624 11500 58676 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 48780 10752 48832 10804
rect 58900 10480 58952 10532
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 57980 10208 58032 10260
rect 10232 10004 10284 10056
rect 1584 9979 1636 9988
rect 1584 9945 1593 9979
rect 1593 9945 1627 9979
rect 1627 9945 1636 9979
rect 1584 9936 1636 9945
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 58900 9664 58952 9716
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 58348 9163 58400 9172
rect 58348 9129 58357 9163
rect 58357 9129 58391 9163
rect 58391 9129 58400 9163
rect 58348 9120 58400 9129
rect 58900 8848 58952 8900
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 58072 8576 58124 8628
rect 9312 8440 9364 8492
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 58900 8304 58952 8356
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 58900 7216 58952 7268
rect 49240 7148 49292 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 2688 6783 2740 6792
rect 2688 6749 2697 6783
rect 2697 6749 2731 6783
rect 2731 6749 2740 6783
rect 2688 6740 2740 6749
rect 940 6672 992 6724
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 4620 5176 4672 5228
rect 940 5108 992 5160
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 9036 3476 9088 3528
rect 940 3408 992 3460
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 12808 2635 12860 2644
rect 12808 2601 12817 2635
rect 12817 2601 12851 2635
rect 12851 2601 12860 2635
rect 12808 2592 12860 2601
rect 15384 2592 15436 2644
rect 42616 2635 42668 2644
rect 42616 2601 42625 2635
rect 42625 2601 42659 2635
rect 42659 2601 42668 2635
rect 42616 2592 42668 2601
rect 49792 2592 49844 2644
rect 2596 2363 2648 2372
rect 2596 2329 2605 2363
rect 2605 2329 2639 2363
rect 2639 2329 2648 2363
rect 2596 2320 2648 2329
rect 11796 2456 11848 2508
rect 12624 2431 12676 2440
rect 12624 2397 12633 2431
rect 12633 2397 12667 2431
rect 12667 2397 12676 2431
rect 12624 2388 12676 2397
rect 17592 2431 17644 2440
rect 17592 2397 17601 2431
rect 17601 2397 17635 2431
rect 17635 2397 17644 2431
rect 17592 2388 17644 2397
rect 22560 2431 22612 2440
rect 22560 2397 22569 2431
rect 22569 2397 22603 2431
rect 22603 2397 22612 2431
rect 22560 2388 22612 2397
rect 7564 2363 7616 2372
rect 7564 2329 7573 2363
rect 7573 2329 7607 2363
rect 7607 2329 7616 2363
rect 7564 2320 7616 2329
rect 9220 2320 9272 2372
rect 27712 2363 27764 2372
rect 27712 2329 27721 2363
rect 27721 2329 27755 2363
rect 27755 2329 27764 2363
rect 27712 2320 27764 2329
rect 45652 2456 45704 2508
rect 47676 2456 47728 2508
rect 4068 2295 4120 2304
rect 4068 2261 4077 2295
rect 4077 2261 4111 2295
rect 4111 2261 4120 2295
rect 4068 2252 4120 2261
rect 12440 2252 12492 2304
rect 32404 2320 32456 2372
rect 38660 2431 38712 2440
rect 38660 2397 38669 2431
rect 38669 2397 38703 2431
rect 38703 2397 38712 2431
rect 38660 2388 38712 2397
rect 42432 2431 42484 2440
rect 42432 2397 42441 2431
rect 42441 2397 42475 2431
rect 42475 2397 42484 2431
rect 42432 2388 42484 2397
rect 47216 2388 47268 2440
rect 52460 2388 52512 2440
rect 37372 2320 37424 2372
rect 57244 2363 57296 2372
rect 57244 2329 57253 2363
rect 57253 2329 57287 2363
rect 57287 2329 57296 2363
rect 57244 2320 57296 2329
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 4068 1980 4120 2032
rect 42248 1980 42300 2032
<< metal2 >>
rect 14922 59200 14978 60000
rect 44914 59200 44970 60000
rect 940 57384 992 57390
rect 940 57326 992 57332
rect 952 56953 980 57326
rect 3056 57248 3108 57254
rect 3056 57190 3108 57196
rect 938 56944 994 56953
rect 938 56879 994 56888
rect 940 55684 992 55690
rect 940 55626 992 55632
rect 952 55321 980 55626
rect 938 55312 994 55321
rect 938 55247 994 55256
rect 1584 54120 1636 54126
rect 1584 54062 1636 54068
rect 1596 53825 1624 54062
rect 2872 53984 2924 53990
rect 2872 53926 2924 53932
rect 1582 53816 1638 53825
rect 1582 53751 1638 53760
rect 1584 52488 1636 52494
rect 1582 52456 1584 52465
rect 1636 52456 1638 52465
rect 1582 52391 1638 52400
rect 2688 50924 2740 50930
rect 2688 50866 2740 50872
rect 940 50856 992 50862
rect 940 50798 992 50804
rect 952 50425 980 50798
rect 938 50416 994 50425
rect 938 50351 994 50360
rect 2228 49224 2280 49230
rect 2228 49166 2280 49172
rect 940 49156 992 49162
rect 940 49098 992 49104
rect 952 48793 980 49098
rect 938 48784 994 48793
rect 938 48719 994 48728
rect 940 47592 992 47598
rect 940 47534 992 47540
rect 952 47161 980 47534
rect 938 47152 994 47161
rect 938 47087 994 47096
rect 1584 45892 1636 45898
rect 1584 45834 1636 45840
rect 1596 45529 1624 45834
rect 1582 45520 1638 45529
rect 1582 45455 1638 45464
rect 1584 44328 1636 44334
rect 1584 44270 1636 44276
rect 1596 44169 1624 44270
rect 1582 44160 1638 44169
rect 1582 44095 1638 44104
rect 940 42628 992 42634
rect 940 42570 992 42576
rect 952 42265 980 42570
rect 938 42256 994 42265
rect 938 42191 994 42200
rect 1400 41132 1452 41138
rect 1400 41074 1452 41080
rect 1216 41064 1268 41070
rect 1216 41006 1268 41012
rect 1228 40633 1256 41006
rect 1214 40624 1270 40633
rect 1214 40559 1270 40568
rect 1412 40050 1440 41074
rect 1400 40044 1452 40050
rect 1400 39986 1452 39992
rect 1412 39642 1440 39986
rect 1952 39840 2004 39846
rect 1952 39782 2004 39788
rect 1400 39636 1452 39642
rect 1400 39578 1452 39584
rect 938 38992 994 39001
rect 938 38927 940 38936
rect 992 38927 994 38936
rect 940 38898 992 38904
rect 1964 38554 1992 39782
rect 1952 38548 2004 38554
rect 1952 38490 2004 38496
rect 1860 38344 1912 38350
rect 1860 38286 1912 38292
rect 1872 38026 1900 38286
rect 1872 37998 2084 38026
rect 1582 37360 1638 37369
rect 1582 37295 1638 37304
rect 1596 37262 1624 37295
rect 1584 37256 1636 37262
rect 1584 37198 1636 37204
rect 938 35728 994 35737
rect 938 35663 940 35672
rect 992 35663 994 35672
rect 940 35634 992 35640
rect 938 34096 994 34105
rect 938 34031 940 34040
rect 992 34031 994 34040
rect 940 34002 992 34008
rect 940 32836 992 32842
rect 940 32778 992 32784
rect 952 32473 980 32778
rect 1400 32768 1452 32774
rect 1400 32710 1452 32716
rect 1412 32570 1440 32710
rect 1400 32564 1452 32570
rect 1400 32506 1452 32512
rect 938 32464 994 32473
rect 938 32399 994 32408
rect 940 31272 992 31278
rect 940 31214 992 31220
rect 952 30841 980 31214
rect 938 30832 994 30841
rect 938 30767 994 30776
rect 940 29572 992 29578
rect 940 29514 992 29520
rect 952 29209 980 29514
rect 1400 29504 1452 29510
rect 1400 29446 1452 29452
rect 1412 29306 1440 29446
rect 1400 29300 1452 29306
rect 1400 29242 1452 29248
rect 938 29200 994 29209
rect 938 29135 994 29144
rect 2056 28762 2084 37998
rect 2240 36038 2268 49166
rect 2596 47660 2648 47666
rect 2596 47602 2648 47608
rect 2608 41970 2636 47602
rect 2516 41942 2636 41970
rect 2412 39364 2464 39370
rect 2412 39306 2464 39312
rect 2424 38826 2452 39306
rect 2412 38820 2464 38826
rect 2412 38762 2464 38768
rect 2424 37942 2452 38762
rect 2516 38282 2544 41942
rect 2700 40610 2728 50866
rect 2608 40582 2728 40610
rect 2608 39098 2636 40582
rect 2688 40520 2740 40526
rect 2688 40462 2740 40468
rect 2700 40186 2728 40462
rect 2688 40180 2740 40186
rect 2688 40122 2740 40128
rect 2596 39092 2648 39098
rect 2596 39034 2648 39040
rect 2504 38276 2556 38282
rect 2504 38218 2556 38224
rect 2608 38010 2636 39034
rect 2688 38548 2740 38554
rect 2688 38490 2740 38496
rect 2700 38350 2728 38490
rect 2688 38344 2740 38350
rect 2688 38286 2740 38292
rect 2884 38298 2912 53926
rect 2964 40384 3016 40390
rect 2964 40326 3016 40332
rect 2976 39370 3004 40326
rect 2964 39364 3016 39370
rect 2964 39306 3016 39312
rect 2596 38004 2648 38010
rect 2596 37946 2648 37952
rect 2412 37936 2464 37942
rect 2412 37878 2464 37884
rect 2424 36854 2452 37878
rect 2412 36848 2464 36854
rect 2412 36790 2464 36796
rect 2424 36106 2452 36790
rect 2700 36582 2728 38286
rect 2884 38270 3004 38298
rect 2872 38208 2924 38214
rect 2872 38150 2924 38156
rect 2884 38010 2912 38150
rect 2872 38004 2924 38010
rect 2872 37946 2924 37952
rect 2976 37806 3004 38270
rect 2964 37800 3016 37806
rect 2964 37742 3016 37748
rect 2780 37256 2832 37262
rect 2780 37198 2832 37204
rect 2688 36576 2740 36582
rect 2688 36518 2740 36524
rect 2412 36100 2464 36106
rect 2412 36042 2464 36048
rect 2228 36032 2280 36038
rect 2228 35974 2280 35980
rect 2424 34678 2452 36042
rect 2700 35494 2728 36518
rect 2792 36378 2820 37198
rect 2872 36576 2924 36582
rect 3068 36530 3096 57190
rect 4214 57148 4522 57157
rect 4214 57146 4220 57148
rect 4276 57146 4300 57148
rect 4356 57146 4380 57148
rect 4436 57146 4460 57148
rect 4516 57146 4522 57148
rect 4276 57094 4278 57146
rect 4458 57094 4460 57146
rect 4214 57092 4220 57094
rect 4276 57092 4300 57094
rect 4356 57092 4380 57094
rect 4436 57092 4460 57094
rect 4516 57092 4522 57094
rect 4214 57083 4522 57092
rect 4214 56060 4522 56069
rect 4214 56058 4220 56060
rect 4276 56058 4300 56060
rect 4356 56058 4380 56060
rect 4436 56058 4460 56060
rect 4516 56058 4522 56060
rect 4276 56006 4278 56058
rect 4458 56006 4460 56058
rect 4214 56004 4220 56006
rect 4276 56004 4300 56006
rect 4356 56004 4380 56006
rect 4436 56004 4460 56006
rect 4516 56004 4522 56006
rect 4214 55995 4522 56004
rect 4214 54972 4522 54981
rect 4214 54970 4220 54972
rect 4276 54970 4300 54972
rect 4356 54970 4380 54972
rect 4436 54970 4460 54972
rect 4516 54970 4522 54972
rect 4276 54918 4278 54970
rect 4458 54918 4460 54970
rect 4214 54916 4220 54918
rect 4276 54916 4300 54918
rect 4356 54916 4380 54918
rect 4436 54916 4460 54918
rect 4516 54916 4522 54918
rect 4214 54907 4522 54916
rect 4214 53884 4522 53893
rect 4214 53882 4220 53884
rect 4276 53882 4300 53884
rect 4356 53882 4380 53884
rect 4436 53882 4460 53884
rect 4516 53882 4522 53884
rect 4276 53830 4278 53882
rect 4458 53830 4460 53882
rect 4214 53828 4220 53830
rect 4276 53828 4300 53830
rect 4356 53828 4380 53830
rect 4436 53828 4460 53830
rect 4516 53828 4522 53830
rect 4214 53819 4522 53828
rect 4214 52796 4522 52805
rect 4214 52794 4220 52796
rect 4276 52794 4300 52796
rect 4356 52794 4380 52796
rect 4436 52794 4460 52796
rect 4516 52794 4522 52796
rect 4276 52742 4278 52794
rect 4458 52742 4460 52794
rect 4214 52740 4220 52742
rect 4276 52740 4300 52742
rect 4356 52740 4380 52742
rect 4436 52740 4460 52742
rect 4516 52740 4522 52742
rect 4214 52731 4522 52740
rect 5540 52488 5592 52494
rect 5540 52430 5592 52436
rect 4214 51708 4522 51717
rect 4214 51706 4220 51708
rect 4276 51706 4300 51708
rect 4356 51706 4380 51708
rect 4436 51706 4460 51708
rect 4516 51706 4522 51708
rect 4276 51654 4278 51706
rect 4458 51654 4460 51706
rect 4214 51652 4220 51654
rect 4276 51652 4300 51654
rect 4356 51652 4380 51654
rect 4436 51652 4460 51654
rect 4516 51652 4522 51654
rect 4214 51643 4522 51652
rect 4214 50620 4522 50629
rect 4214 50618 4220 50620
rect 4276 50618 4300 50620
rect 4356 50618 4380 50620
rect 4436 50618 4460 50620
rect 4516 50618 4522 50620
rect 4276 50566 4278 50618
rect 4458 50566 4460 50618
rect 4214 50564 4220 50566
rect 4276 50564 4300 50566
rect 4356 50564 4380 50566
rect 4436 50564 4460 50566
rect 4516 50564 4522 50566
rect 4214 50555 4522 50564
rect 4214 49532 4522 49541
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49467 4522 49476
rect 4214 48444 4522 48453
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48379 4522 48388
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 3792 44396 3844 44402
rect 3792 44338 3844 44344
rect 3516 39976 3568 39982
rect 3516 39918 3568 39924
rect 3240 39840 3292 39846
rect 3240 39782 3292 39788
rect 3252 39438 3280 39782
rect 3528 39642 3556 39918
rect 3516 39636 3568 39642
rect 3516 39578 3568 39584
rect 3804 39506 3832 44338
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 5552 41414 5580 52430
rect 6552 45960 6604 45966
rect 6552 45902 6604 45908
rect 5552 41386 5764 41414
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 3884 40112 3936 40118
rect 3884 40054 3936 40060
rect 3792 39500 3844 39506
rect 3792 39442 3844 39448
rect 3240 39432 3292 39438
rect 3240 39374 3292 39380
rect 3240 39296 3292 39302
rect 3240 39238 3292 39244
rect 3332 39296 3384 39302
rect 3332 39238 3384 39244
rect 3252 37806 3280 39238
rect 3344 37874 3372 39238
rect 3804 39098 3832 39442
rect 3792 39092 3844 39098
rect 3792 39034 3844 39040
rect 3700 38888 3752 38894
rect 3700 38830 3752 38836
rect 3516 38752 3568 38758
rect 3516 38694 3568 38700
rect 3424 38344 3476 38350
rect 3424 38286 3476 38292
rect 3436 38010 3464 38286
rect 3528 38010 3556 38694
rect 3424 38004 3476 38010
rect 3424 37946 3476 37952
rect 3516 38004 3568 38010
rect 3516 37946 3568 37952
rect 3332 37868 3384 37874
rect 3332 37810 3384 37816
rect 3240 37800 3292 37806
rect 2872 36518 2924 36524
rect 2780 36372 2832 36378
rect 2780 36314 2832 36320
rect 2792 36122 2820 36314
rect 2884 36242 2912 36518
rect 2976 36502 3096 36530
rect 3160 37760 3240 37788
rect 2872 36236 2924 36242
rect 2872 36178 2924 36184
rect 2792 36094 2912 36122
rect 2884 35698 2912 36094
rect 2872 35692 2924 35698
rect 2872 35634 2924 35640
rect 2688 35488 2740 35494
rect 2688 35430 2740 35436
rect 2596 35080 2648 35086
rect 2596 35022 2648 35028
rect 2608 34678 2636 35022
rect 2412 34672 2464 34678
rect 2412 34614 2464 34620
rect 2596 34672 2648 34678
rect 2596 34614 2648 34620
rect 2424 32502 2452 34614
rect 2608 33998 2636 34614
rect 2596 33992 2648 33998
rect 2596 33934 2648 33940
rect 2872 33992 2924 33998
rect 2872 33934 2924 33940
rect 2884 32570 2912 33934
rect 2872 32564 2924 32570
rect 2872 32506 2924 32512
rect 2412 32496 2464 32502
rect 2412 32438 2464 32444
rect 2424 30666 2452 32438
rect 2872 32360 2924 32366
rect 2872 32302 2924 32308
rect 2504 32224 2556 32230
rect 2504 32166 2556 32172
rect 2516 31890 2544 32166
rect 2884 32026 2912 32302
rect 2872 32020 2924 32026
rect 2872 31962 2924 31968
rect 2504 31884 2556 31890
rect 2504 31826 2556 31832
rect 2688 31340 2740 31346
rect 2688 31282 2740 31288
rect 2412 30660 2464 30666
rect 2412 30602 2464 30608
rect 2424 29238 2452 30602
rect 2700 30598 2728 31282
rect 2688 30592 2740 30598
rect 2688 30534 2740 30540
rect 2700 30258 2728 30534
rect 2688 30252 2740 30258
rect 2688 30194 2740 30200
rect 2976 30138 3004 36502
rect 3160 36106 3188 37760
rect 3240 37742 3292 37748
rect 3344 37330 3372 37810
rect 3712 37330 3740 38830
rect 3792 38344 3844 38350
rect 3792 38286 3844 38292
rect 3332 37324 3384 37330
rect 3252 37284 3332 37312
rect 3252 36310 3280 37284
rect 3332 37266 3384 37272
rect 3700 37324 3752 37330
rect 3700 37266 3752 37272
rect 3712 36718 3740 37266
rect 3608 36712 3660 36718
rect 3608 36654 3660 36660
rect 3700 36712 3752 36718
rect 3700 36654 3752 36660
rect 3332 36644 3384 36650
rect 3332 36586 3384 36592
rect 3240 36304 3292 36310
rect 3240 36246 3292 36252
rect 3148 36100 3200 36106
rect 3148 36042 3200 36048
rect 3160 35630 3188 36042
rect 3148 35624 3200 35630
rect 3148 35566 3200 35572
rect 3056 34944 3108 34950
rect 3056 34886 3108 34892
rect 3068 33998 3096 34886
rect 3160 34542 3188 35566
rect 3344 35290 3372 36586
rect 3620 36378 3648 36654
rect 3608 36372 3660 36378
rect 3608 36314 3660 36320
rect 3424 36168 3476 36174
rect 3424 36110 3476 36116
rect 3436 35834 3464 36110
rect 3424 35828 3476 35834
rect 3424 35770 3476 35776
rect 3424 35488 3476 35494
rect 3424 35430 3476 35436
rect 3332 35284 3384 35290
rect 3332 35226 3384 35232
rect 3436 35193 3464 35430
rect 3422 35184 3478 35193
rect 3344 35142 3422 35170
rect 3148 34536 3200 34542
rect 3148 34478 3200 34484
rect 3056 33992 3108 33998
rect 3056 33934 3108 33940
rect 3160 32366 3188 34478
rect 3344 33930 3372 35142
rect 3422 35119 3478 35128
rect 3804 35034 3832 38286
rect 3896 35290 3924 40054
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4620 39432 4672 39438
rect 4620 39374 4672 39380
rect 4068 39296 4120 39302
rect 4068 39238 4120 39244
rect 4080 38554 4108 39238
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4632 38554 4660 39374
rect 4804 39296 4856 39302
rect 4804 39238 4856 39244
rect 4068 38548 4120 38554
rect 4068 38490 4120 38496
rect 4620 38548 4672 38554
rect 4620 38490 4672 38496
rect 4816 38350 4844 39238
rect 5264 38888 5316 38894
rect 5264 38830 5316 38836
rect 5540 38888 5592 38894
rect 5540 38830 5592 38836
rect 5276 38554 5304 38830
rect 5264 38548 5316 38554
rect 5264 38490 5316 38496
rect 4252 38344 4304 38350
rect 4252 38286 4304 38292
rect 4804 38344 4856 38350
rect 4804 38286 4856 38292
rect 4264 37874 4292 38286
rect 4252 37868 4304 37874
rect 4252 37810 4304 37816
rect 4620 37800 4672 37806
rect 4620 37742 4672 37748
rect 4068 37664 4120 37670
rect 4068 37606 4120 37612
rect 3976 37188 4028 37194
rect 3976 37130 4028 37136
rect 3988 36378 4016 37130
rect 4080 36378 4108 37606
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4632 37126 4660 37742
rect 5552 37126 5580 38830
rect 5632 38344 5684 38350
rect 5632 38286 5684 38292
rect 4620 37120 4672 37126
rect 4620 37062 4672 37068
rect 5356 37120 5408 37126
rect 5356 37062 5408 37068
rect 5540 37120 5592 37126
rect 5540 37062 5592 37068
rect 5368 36854 5396 37062
rect 5356 36848 5408 36854
rect 5356 36790 5408 36796
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 3976 36372 4028 36378
rect 3976 36314 4028 36320
rect 4068 36372 4120 36378
rect 4068 36314 4120 36320
rect 3976 36168 4028 36174
rect 3976 36110 4028 36116
rect 4528 36168 4580 36174
rect 4528 36110 4580 36116
rect 3988 35494 4016 36110
rect 4540 35834 4568 36110
rect 4620 36100 4672 36106
rect 4620 36042 4672 36048
rect 4528 35828 4580 35834
rect 4528 35770 4580 35776
rect 4068 35692 4120 35698
rect 4068 35634 4120 35640
rect 3976 35488 4028 35494
rect 3976 35430 4028 35436
rect 3884 35284 3936 35290
rect 3884 35226 3936 35232
rect 3700 35012 3752 35018
rect 3804 35006 4016 35034
rect 3700 34954 3752 34960
rect 3712 34592 3740 34954
rect 3884 34604 3936 34610
rect 3712 34564 3884 34592
rect 3884 34546 3936 34552
rect 3424 34536 3476 34542
rect 3424 34478 3476 34484
rect 3436 34202 3464 34478
rect 3424 34196 3476 34202
rect 3424 34138 3476 34144
rect 3332 33924 3384 33930
rect 3332 33866 3384 33872
rect 3148 32360 3200 32366
rect 3200 32320 3280 32348
rect 3148 32302 3200 32308
rect 3148 31136 3200 31142
rect 3148 31078 3200 31084
rect 3160 30938 3188 31078
rect 3148 30932 3200 30938
rect 3148 30874 3200 30880
rect 3148 30796 3200 30802
rect 3148 30738 3200 30744
rect 3160 30326 3188 30738
rect 3148 30320 3200 30326
rect 3148 30262 3200 30268
rect 2976 30110 3188 30138
rect 3160 29510 3188 30110
rect 2964 29504 3016 29510
rect 2964 29446 3016 29452
rect 3148 29504 3200 29510
rect 3148 29446 3200 29452
rect 2976 29238 3004 29446
rect 2412 29232 2464 29238
rect 2412 29174 2464 29180
rect 2964 29232 3016 29238
rect 2964 29174 3016 29180
rect 3252 29170 3280 32320
rect 3344 31822 3372 33866
rect 3516 32768 3568 32774
rect 3516 32710 3568 32716
rect 3424 32292 3476 32298
rect 3424 32234 3476 32240
rect 3436 32026 3464 32234
rect 3528 32026 3556 32710
rect 3896 32366 3924 34546
rect 3792 32360 3844 32366
rect 3792 32302 3844 32308
rect 3884 32360 3936 32366
rect 3884 32302 3936 32308
rect 3424 32020 3476 32026
rect 3424 31962 3476 31968
rect 3516 32020 3568 32026
rect 3516 31962 3568 31968
rect 3332 31816 3384 31822
rect 3332 31758 3384 31764
rect 3344 30734 3372 31758
rect 3516 31680 3568 31686
rect 3804 31634 3832 32302
rect 3568 31628 3832 31634
rect 3516 31622 3832 31628
rect 3528 31606 3832 31622
rect 3896 31346 3924 32302
rect 3884 31340 3936 31346
rect 3884 31282 3936 31288
rect 3700 31272 3752 31278
rect 3700 31214 3752 31220
rect 3792 31272 3844 31278
rect 3792 31214 3844 31220
rect 3424 31136 3476 31142
rect 3424 31078 3476 31084
rect 3436 30802 3464 31078
rect 3712 30938 3740 31214
rect 3700 30932 3752 30938
rect 3700 30874 3752 30880
rect 3424 30796 3476 30802
rect 3424 30738 3476 30744
rect 3332 30728 3384 30734
rect 3332 30670 3384 30676
rect 3344 30122 3372 30670
rect 3700 30184 3752 30190
rect 3700 30126 3752 30132
rect 3332 30116 3384 30122
rect 3332 30058 3384 30064
rect 3608 30048 3660 30054
rect 3608 29990 3660 29996
rect 3620 29850 3648 29990
rect 3712 29850 3740 30126
rect 3608 29844 3660 29850
rect 3608 29786 3660 29792
rect 3700 29844 3752 29850
rect 3700 29786 3752 29792
rect 3240 29164 3292 29170
rect 3240 29106 3292 29112
rect 2044 28756 2096 28762
rect 2044 28698 2096 28704
rect 2688 28076 2740 28082
rect 2688 28018 2740 28024
rect 1584 28008 1636 28014
rect 1584 27950 1636 27956
rect 1596 27577 1624 27950
rect 1582 27568 1638 27577
rect 1582 27503 1638 27512
rect 2412 27396 2464 27402
rect 2412 27338 2464 27344
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 1412 26042 1440 26318
rect 1584 26308 1636 26314
rect 1584 26250 1636 26256
rect 1596 26217 1624 26250
rect 1582 26208 1638 26217
rect 1582 26143 1638 26152
rect 1400 26036 1452 26042
rect 1400 25978 1452 25984
rect 2424 25974 2452 27338
rect 2700 27334 2728 28018
rect 2780 27872 2832 27878
rect 2780 27814 2832 27820
rect 2688 27328 2740 27334
rect 2688 27270 2740 27276
rect 2700 26858 2728 27270
rect 2792 26926 2820 27814
rect 3252 27606 3280 29106
rect 3608 28960 3660 28966
rect 3608 28902 3660 28908
rect 3620 28558 3648 28902
rect 3608 28552 3660 28558
rect 3608 28494 3660 28500
rect 3700 28552 3752 28558
rect 3700 28494 3752 28500
rect 3424 28008 3476 28014
rect 3424 27950 3476 27956
rect 3436 27674 3464 27950
rect 3424 27668 3476 27674
rect 3424 27610 3476 27616
rect 3240 27600 3292 27606
rect 3240 27542 3292 27548
rect 3240 27464 3292 27470
rect 3240 27406 3292 27412
rect 3424 27464 3476 27470
rect 3424 27406 3476 27412
rect 2872 27396 2924 27402
rect 2872 27338 2924 27344
rect 2884 27130 2912 27338
rect 2872 27124 2924 27130
rect 2872 27066 2924 27072
rect 2780 26920 2832 26926
rect 2780 26862 2832 26868
rect 2688 26852 2740 26858
rect 2688 26794 2740 26800
rect 3252 26450 3280 27406
rect 3436 27130 3464 27406
rect 3424 27124 3476 27130
rect 3424 27066 3476 27072
rect 3332 26784 3384 26790
rect 3332 26726 3384 26732
rect 3240 26444 3292 26450
rect 3240 26386 3292 26392
rect 2412 25968 2464 25974
rect 2412 25910 2464 25916
rect 940 24744 992 24750
rect 940 24686 992 24692
rect 952 24313 980 24686
rect 938 24304 994 24313
rect 938 24239 994 24248
rect 2424 24138 2452 25910
rect 3148 25832 3200 25838
rect 3148 25774 3200 25780
rect 2688 24812 2740 24818
rect 2688 24754 2740 24760
rect 2412 24132 2464 24138
rect 2412 24074 2464 24080
rect 940 23044 992 23050
rect 940 22986 992 22992
rect 952 22681 980 22986
rect 1400 22976 1452 22982
rect 1400 22918 1452 22924
rect 1412 22778 1440 22918
rect 1400 22772 1452 22778
rect 1400 22714 1452 22720
rect 2424 22710 2452 24074
rect 2700 24070 2728 24754
rect 3056 24608 3108 24614
rect 3056 24550 3108 24556
rect 3068 24410 3096 24550
rect 3056 24404 3108 24410
rect 3056 24346 3108 24352
rect 3160 24274 3188 25774
rect 3240 25696 3292 25702
rect 3240 25638 3292 25644
rect 3252 25362 3280 25638
rect 3344 25430 3372 26726
rect 3424 25764 3476 25770
rect 3424 25706 3476 25712
rect 3436 25498 3464 25706
rect 3424 25492 3476 25498
rect 3424 25434 3476 25440
rect 3332 25424 3384 25430
rect 3332 25366 3384 25372
rect 3240 25356 3292 25362
rect 3240 25298 3292 25304
rect 3344 24410 3372 25366
rect 3712 25362 3740 28494
rect 3804 28490 3832 31214
rect 3896 30734 3924 31282
rect 3884 30728 3936 30734
rect 3884 30670 3936 30676
rect 3792 28484 3844 28490
rect 3792 28426 3844 28432
rect 3988 28218 4016 35006
rect 4080 34746 4108 35634
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4068 34740 4120 34746
rect 4068 34682 4120 34688
rect 4632 34474 4660 36042
rect 4988 36032 5040 36038
rect 4988 35974 5040 35980
rect 5000 35766 5028 35974
rect 4988 35760 5040 35766
rect 4988 35702 5040 35708
rect 4712 35488 4764 35494
rect 4712 35430 4764 35436
rect 4724 35290 4752 35430
rect 4712 35284 4764 35290
rect 4712 35226 4764 35232
rect 4988 35080 5040 35086
rect 4988 35022 5040 35028
rect 4620 34468 4672 34474
rect 4620 34410 4672 34416
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4804 33856 4856 33862
rect 4804 33798 4856 33804
rect 4816 33658 4844 33798
rect 5000 33658 5028 35022
rect 5172 34944 5224 34950
rect 5172 34886 5224 34892
rect 5184 33998 5212 34886
rect 5172 33992 5224 33998
rect 5172 33934 5224 33940
rect 4804 33652 4856 33658
rect 4804 33594 4856 33600
rect 4988 33652 5040 33658
rect 4988 33594 5040 33600
rect 5000 33454 5028 33594
rect 4988 33448 5040 33454
rect 4988 33390 5040 33396
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4804 32768 4856 32774
rect 4804 32710 4856 32716
rect 4816 32434 4844 32710
rect 4804 32428 4856 32434
rect 4804 32370 4856 32376
rect 4068 32224 4120 32230
rect 4068 32166 4120 32172
rect 4620 32224 4672 32230
rect 4620 32166 4672 32172
rect 4988 32224 5040 32230
rect 4988 32166 5040 32172
rect 4080 31686 4108 32166
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4632 32026 4660 32166
rect 5000 32026 5028 32166
rect 4620 32020 4672 32026
rect 4620 31962 4672 31968
rect 4988 32020 5040 32026
rect 4988 31962 5040 31968
rect 4988 31884 5040 31890
rect 4988 31826 5040 31832
rect 4896 31816 4948 31822
rect 4896 31758 4948 31764
rect 4344 31748 4396 31754
rect 4344 31690 4396 31696
rect 4068 31680 4120 31686
rect 4068 31622 4120 31628
rect 4356 31346 4384 31690
rect 4908 31482 4936 31758
rect 4896 31476 4948 31482
rect 4896 31418 4948 31424
rect 5000 31414 5028 31826
rect 4988 31408 5040 31414
rect 4988 31350 5040 31356
rect 5184 31346 5212 33934
rect 5264 33584 5316 33590
rect 5264 33526 5316 33532
rect 5276 31822 5304 33526
rect 5540 33312 5592 33318
rect 5540 33254 5592 33260
rect 5264 31816 5316 31822
rect 5264 31758 5316 31764
rect 5356 31748 5408 31754
rect 5356 31690 5408 31696
rect 4160 31340 4212 31346
rect 4080 31300 4160 31328
rect 4080 30394 4108 31300
rect 4160 31282 4212 31288
rect 4344 31340 4396 31346
rect 4344 31282 4396 31288
rect 5172 31340 5224 31346
rect 5172 31282 5224 31288
rect 4620 31136 4672 31142
rect 4620 31078 4672 31084
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30802 4660 31078
rect 4620 30796 4672 30802
rect 4620 30738 4672 30744
rect 5080 30660 5132 30666
rect 5080 30602 5132 30608
rect 4068 30388 4120 30394
rect 4068 30330 4120 30336
rect 4068 30252 4120 30258
rect 4068 30194 4120 30200
rect 4080 29850 4108 30194
rect 4896 30048 4948 30054
rect 4896 29990 4948 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4068 29844 4120 29850
rect 4068 29786 4120 29792
rect 4908 29714 4936 29990
rect 5092 29850 5120 30602
rect 5368 30258 5396 31690
rect 5448 30592 5500 30598
rect 5448 30534 5500 30540
rect 5172 30252 5224 30258
rect 5356 30252 5408 30258
rect 5172 30194 5224 30200
rect 5276 30212 5356 30240
rect 5080 29844 5132 29850
rect 5080 29786 5132 29792
rect 4896 29708 4948 29714
rect 4896 29650 4948 29656
rect 4804 29572 4856 29578
rect 4804 29514 4856 29520
rect 4712 29232 4764 29238
rect 4712 29174 4764 29180
rect 4252 29096 4304 29102
rect 4080 29044 4252 29050
rect 4080 29038 4304 29044
rect 4080 29022 4292 29038
rect 4080 28762 4108 29022
rect 4620 28960 4672 28966
rect 4620 28902 4672 28908
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4068 28756 4120 28762
rect 4068 28698 4120 28704
rect 4632 28558 4660 28902
rect 4724 28762 4752 29174
rect 4712 28756 4764 28762
rect 4712 28698 4764 28704
rect 4816 28626 4844 29514
rect 4988 29164 5040 29170
rect 4988 29106 5040 29112
rect 4896 28756 4948 28762
rect 4896 28698 4948 28704
rect 4804 28620 4856 28626
rect 4804 28562 4856 28568
rect 4068 28552 4120 28558
rect 4068 28494 4120 28500
rect 4160 28552 4212 28558
rect 4160 28494 4212 28500
rect 4620 28552 4672 28558
rect 4620 28494 4672 28500
rect 4080 28218 4108 28494
rect 3976 28212 4028 28218
rect 3976 28154 4028 28160
rect 4068 28212 4120 28218
rect 4068 28154 4120 28160
rect 4172 27946 4200 28494
rect 4908 28490 4936 28698
rect 5000 28490 5028 29106
rect 4896 28484 4948 28490
rect 4896 28426 4948 28432
rect 4988 28484 5040 28490
rect 4988 28426 5040 28432
rect 4712 28416 4764 28422
rect 4712 28358 4764 28364
rect 4160 27940 4212 27946
rect 4160 27882 4212 27888
rect 4620 27872 4672 27878
rect 4620 27814 4672 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4632 27674 4660 27814
rect 4620 27668 4672 27674
rect 4620 27610 4672 27616
rect 4160 27396 4212 27402
rect 4160 27338 4212 27344
rect 4172 27130 4200 27338
rect 4724 27130 4752 28358
rect 4804 28076 4856 28082
rect 4804 28018 4856 28024
rect 4816 27334 4844 28018
rect 4804 27328 4856 27334
rect 4804 27270 4856 27276
rect 4908 27146 4936 28426
rect 5000 28014 5028 28426
rect 4988 28008 5040 28014
rect 4988 27950 5040 27956
rect 4160 27124 4212 27130
rect 4160 27066 4212 27072
rect 4712 27124 4764 27130
rect 4712 27066 4764 27072
rect 4816 27118 4936 27146
rect 4816 27010 4844 27118
rect 4724 26982 4844 27010
rect 5000 26994 5028 27950
rect 4988 26988 5040 26994
rect 4620 26920 4672 26926
rect 4620 26862 4672 26868
rect 3792 26852 3844 26858
rect 3792 26794 3844 26800
rect 3804 25498 3832 26794
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4632 26382 4660 26862
rect 3976 26376 4028 26382
rect 3976 26318 4028 26324
rect 4620 26376 4672 26382
rect 4620 26318 4672 26324
rect 3884 26240 3936 26246
rect 3884 26182 3936 26188
rect 3896 25906 3924 26182
rect 3884 25900 3936 25906
rect 3884 25842 3936 25848
rect 3792 25492 3844 25498
rect 3792 25434 3844 25440
rect 3700 25356 3752 25362
rect 3700 25298 3752 25304
rect 3712 24954 3740 25298
rect 3700 24948 3752 24954
rect 3752 24908 3832 24936
rect 3700 24890 3752 24896
rect 3700 24744 3752 24750
rect 3700 24686 3752 24692
rect 3712 24410 3740 24686
rect 3332 24404 3384 24410
rect 3332 24346 3384 24352
rect 3700 24404 3752 24410
rect 3700 24346 3752 24352
rect 3148 24268 3200 24274
rect 3148 24210 3200 24216
rect 2872 24132 2924 24138
rect 2872 24074 2924 24080
rect 2688 24064 2740 24070
rect 2688 24006 2740 24012
rect 2700 23866 2728 24006
rect 2688 23860 2740 23866
rect 2688 23802 2740 23808
rect 2412 22704 2464 22710
rect 938 22672 994 22681
rect 2412 22646 2464 22652
rect 938 22607 994 22616
rect 940 21480 992 21486
rect 940 21422 992 21428
rect 952 21049 980 21422
rect 938 21040 994 21049
rect 938 20975 994 20984
rect 2424 20874 2452 22646
rect 2884 22166 2912 24074
rect 3160 22642 3188 24210
rect 3240 24200 3292 24206
rect 3240 24142 3292 24148
rect 3252 23866 3280 24142
rect 3344 24138 3372 24346
rect 3332 24132 3384 24138
rect 3332 24074 3384 24080
rect 3240 23860 3292 23866
rect 3240 23802 3292 23808
rect 3516 23248 3568 23254
rect 3516 23190 3568 23196
rect 3528 23066 3556 23190
rect 3436 23038 3556 23066
rect 3148 22636 3200 22642
rect 3148 22578 3200 22584
rect 2872 22160 2924 22166
rect 2872 22102 2924 22108
rect 2688 21548 2740 21554
rect 2688 21490 2740 21496
rect 2412 20868 2464 20874
rect 2412 20810 2464 20816
rect 940 19780 992 19786
rect 940 19722 992 19728
rect 952 19417 980 19722
rect 1400 19712 1452 19718
rect 1400 19654 1452 19660
rect 1412 19514 1440 19654
rect 1400 19508 1452 19514
rect 1400 19450 1452 19456
rect 2424 19446 2452 20810
rect 2700 20806 2728 21490
rect 2884 20874 2912 22102
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 3068 21146 3096 21286
rect 3056 21140 3108 21146
rect 3056 21082 3108 21088
rect 3160 20942 3188 22578
rect 3332 22568 3384 22574
rect 3332 22510 3384 22516
rect 3240 22432 3292 22438
rect 3240 22374 3292 22380
rect 3252 22234 3280 22374
rect 3344 22234 3372 22510
rect 3240 22228 3292 22234
rect 3240 22170 3292 22176
rect 3332 22228 3384 22234
rect 3332 22170 3384 22176
rect 3436 22094 3464 23038
rect 3516 22976 3568 22982
rect 3516 22918 3568 22924
rect 3528 22778 3556 22918
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3436 22066 3556 22094
rect 3528 20942 3556 22066
rect 3804 22030 3832 24908
rect 3988 23730 4016 26318
rect 4620 25900 4672 25906
rect 4620 25842 4672 25848
rect 4068 25832 4120 25838
rect 4068 25774 4120 25780
rect 4080 25498 4108 25774
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4632 25498 4660 25842
rect 4068 25492 4120 25498
rect 4068 25434 4120 25440
rect 4620 25492 4672 25498
rect 4620 25434 4672 25440
rect 4724 25294 4752 26982
rect 4988 26930 5040 26936
rect 5092 26858 5120 29786
rect 5184 29782 5212 30194
rect 5172 29776 5224 29782
rect 5172 29718 5224 29724
rect 5276 27402 5304 30212
rect 5356 30194 5408 30200
rect 5460 30138 5488 30534
rect 5552 30258 5580 33254
rect 5644 31482 5672 38286
rect 5736 37874 5764 41386
rect 6564 39506 6592 45902
rect 7564 42696 7616 42702
rect 7564 42638 7616 42644
rect 7576 40050 7604 42638
rect 8300 40112 8352 40118
rect 8300 40054 8352 40060
rect 7564 40044 7616 40050
rect 7564 39986 7616 39992
rect 6552 39500 6604 39506
rect 6552 39442 6604 39448
rect 6564 39098 6592 39442
rect 7748 39432 7800 39438
rect 7748 39374 7800 39380
rect 7196 39296 7248 39302
rect 7196 39238 7248 39244
rect 6552 39092 6604 39098
rect 6552 39034 6604 39040
rect 7208 38010 7236 39238
rect 7760 38486 7788 39374
rect 8312 39098 8340 40054
rect 8392 40044 8444 40050
rect 8392 39986 8444 39992
rect 8208 39092 8260 39098
rect 8208 39034 8260 39040
rect 8300 39092 8352 39098
rect 8300 39034 8352 39040
rect 8220 38978 8248 39034
rect 8404 38978 8432 39986
rect 9864 39976 9916 39982
rect 9864 39918 9916 39924
rect 10140 39976 10192 39982
rect 10140 39918 10192 39924
rect 9876 39642 9904 39918
rect 9864 39636 9916 39642
rect 9864 39578 9916 39584
rect 8668 39432 8720 39438
rect 8668 39374 8720 39380
rect 8680 39098 8708 39374
rect 9128 39296 9180 39302
rect 9128 39238 9180 39244
rect 8668 39092 8720 39098
rect 8668 39034 8720 39040
rect 8220 38950 8432 38978
rect 7932 38888 7984 38894
rect 7932 38830 7984 38836
rect 7944 38554 7972 38830
rect 8404 38554 8432 38950
rect 8484 38956 8536 38962
rect 8484 38898 8536 38904
rect 7932 38548 7984 38554
rect 7932 38490 7984 38496
rect 8392 38548 8444 38554
rect 8392 38490 8444 38496
rect 7748 38480 7800 38486
rect 8496 38434 8524 38898
rect 8760 38888 8812 38894
rect 8760 38830 8812 38836
rect 7748 38422 7800 38428
rect 7472 38412 7524 38418
rect 7472 38354 7524 38360
rect 8404 38406 8524 38434
rect 7484 38010 7512 38354
rect 7748 38344 7800 38350
rect 7748 38286 7800 38292
rect 7196 38004 7248 38010
rect 7196 37946 7248 37952
rect 7472 38004 7524 38010
rect 7472 37946 7524 37952
rect 5724 37868 5776 37874
rect 5724 37810 5776 37816
rect 5736 37466 5764 37810
rect 7288 37664 7340 37670
rect 7288 37606 7340 37612
rect 7300 37466 7328 37606
rect 5724 37460 5776 37466
rect 5724 37402 5776 37408
rect 7288 37460 7340 37466
rect 7288 37402 7340 37408
rect 7656 37324 7708 37330
rect 7656 37266 7708 37272
rect 6092 37188 6144 37194
rect 6092 37130 6144 37136
rect 5724 37120 5776 37126
rect 5724 37062 5776 37068
rect 5736 36786 5764 37062
rect 6104 36786 6132 37130
rect 7472 37120 7524 37126
rect 7472 37062 7524 37068
rect 7484 36922 7512 37062
rect 7668 36922 7696 37266
rect 7472 36916 7524 36922
rect 7472 36858 7524 36864
rect 7656 36916 7708 36922
rect 7656 36858 7708 36864
rect 5724 36780 5776 36786
rect 5724 36722 5776 36728
rect 6092 36780 6144 36786
rect 6092 36722 6144 36728
rect 5736 35630 5764 36722
rect 6104 35766 6132 36722
rect 7012 36644 7064 36650
rect 7012 36586 7064 36592
rect 6460 36100 6512 36106
rect 6460 36042 6512 36048
rect 6472 35834 6500 36042
rect 6184 35828 6236 35834
rect 6184 35770 6236 35776
rect 6460 35828 6512 35834
rect 6460 35770 6512 35776
rect 6092 35760 6144 35766
rect 6092 35702 6144 35708
rect 5724 35624 5776 35630
rect 5724 35566 5776 35572
rect 6196 35290 6224 35770
rect 6184 35284 6236 35290
rect 6184 35226 6236 35232
rect 6644 35080 6696 35086
rect 6644 35022 6696 35028
rect 6000 34604 6052 34610
rect 6000 34546 6052 34552
rect 6012 34202 6040 34546
rect 6000 34196 6052 34202
rect 6000 34138 6052 34144
rect 6552 34196 6604 34202
rect 6552 34138 6604 34144
rect 5908 33924 5960 33930
rect 5908 33866 5960 33872
rect 5920 33658 5948 33866
rect 6564 33658 6592 34138
rect 6656 33658 6684 35022
rect 6736 33856 6788 33862
rect 6736 33798 6788 33804
rect 5908 33652 5960 33658
rect 5908 33594 5960 33600
rect 6552 33652 6604 33658
rect 6552 33594 6604 33600
rect 6644 33652 6696 33658
rect 6644 33594 6696 33600
rect 6460 33584 6512 33590
rect 6460 33526 6512 33532
rect 6000 33516 6052 33522
rect 6000 33458 6052 33464
rect 6368 33516 6420 33522
rect 6368 33458 6420 33464
rect 6012 33318 6040 33458
rect 6380 33386 6408 33458
rect 6368 33380 6420 33386
rect 6368 33322 6420 33328
rect 6000 33312 6052 33318
rect 6000 33254 6052 33260
rect 6380 32774 6408 33322
rect 6472 32978 6500 33526
rect 6748 33522 6776 33798
rect 6736 33516 6788 33522
rect 6736 33458 6788 33464
rect 6460 32972 6512 32978
rect 6460 32914 6512 32920
rect 6368 32768 6420 32774
rect 6368 32710 6420 32716
rect 6380 32026 6408 32710
rect 6368 32020 6420 32026
rect 6368 31962 6420 31968
rect 6380 31804 6408 31962
rect 6460 31816 6512 31822
rect 6380 31776 6460 31804
rect 6276 31748 6328 31754
rect 6276 31690 6328 31696
rect 5632 31476 5684 31482
rect 5632 31418 5684 31424
rect 6288 31346 6316 31690
rect 6092 31340 6144 31346
rect 6092 31282 6144 31288
rect 6276 31340 6328 31346
rect 6276 31282 6328 31288
rect 5816 31272 5868 31278
rect 5816 31214 5868 31220
rect 5828 30734 5856 31214
rect 5908 31204 5960 31210
rect 5908 31146 5960 31152
rect 5816 30728 5868 30734
rect 5816 30670 5868 30676
rect 5920 30394 5948 31146
rect 5908 30388 5960 30394
rect 5908 30330 5960 30336
rect 5540 30252 5592 30258
rect 5540 30194 5592 30200
rect 5368 30110 5488 30138
rect 5368 28422 5396 30110
rect 5448 29300 5500 29306
rect 5448 29242 5500 29248
rect 5460 28626 5488 29242
rect 5448 28620 5500 28626
rect 5448 28562 5500 28568
rect 5552 28422 5580 30194
rect 5632 30116 5684 30122
rect 5632 30058 5684 30064
rect 5644 29102 5672 30058
rect 5920 29850 5948 30330
rect 5908 29844 5960 29850
rect 5908 29786 5960 29792
rect 5816 29572 5868 29578
rect 5816 29514 5868 29520
rect 5632 29096 5684 29102
rect 5632 29038 5684 29044
rect 5356 28416 5408 28422
rect 5356 28358 5408 28364
rect 5540 28416 5592 28422
rect 5540 28358 5592 28364
rect 5368 27878 5396 28358
rect 5356 27872 5408 27878
rect 5356 27814 5408 27820
rect 5644 27470 5672 29038
rect 5828 28762 5856 29514
rect 5908 29164 5960 29170
rect 5908 29106 5960 29112
rect 5920 28762 5948 29106
rect 6104 28762 6132 31282
rect 6184 30592 6236 30598
rect 6184 30534 6236 30540
rect 6196 30258 6224 30534
rect 6184 30252 6236 30258
rect 6184 30194 6236 30200
rect 6288 29238 6316 31282
rect 6380 31210 6408 31776
rect 6460 31758 6512 31764
rect 6368 31204 6420 31210
rect 6368 31146 6420 31152
rect 6368 30728 6420 30734
rect 6368 30670 6420 30676
rect 6380 30598 6408 30670
rect 6748 30598 6776 33458
rect 6828 32972 6880 32978
rect 6828 32914 6880 32920
rect 6368 30592 6420 30598
rect 6368 30534 6420 30540
rect 6736 30592 6788 30598
rect 6736 30534 6788 30540
rect 6276 29232 6328 29238
rect 6276 29174 6328 29180
rect 5816 28756 5868 28762
rect 5816 28698 5868 28704
rect 5908 28756 5960 28762
rect 5908 28698 5960 28704
rect 6092 28756 6144 28762
rect 6092 28698 6144 28704
rect 6380 28218 6408 30534
rect 6840 30326 6868 32914
rect 6920 32020 6972 32026
rect 6920 31962 6972 31968
rect 6932 31346 6960 31962
rect 6920 31340 6972 31346
rect 6920 31282 6972 31288
rect 7024 30938 7052 36586
rect 7288 36576 7340 36582
rect 7288 36518 7340 36524
rect 7300 36174 7328 36518
rect 7288 36168 7340 36174
rect 7288 36110 7340 36116
rect 7300 35222 7328 36110
rect 7288 35216 7340 35222
rect 7286 35184 7288 35193
rect 7340 35184 7342 35193
rect 7286 35119 7342 35128
rect 7760 33590 7788 38286
rect 8404 37874 8432 38406
rect 8772 38350 8800 38830
rect 8668 38344 8720 38350
rect 8668 38286 8720 38292
rect 8760 38344 8812 38350
rect 8760 38286 8812 38292
rect 8680 38010 8708 38286
rect 9036 38208 9088 38214
rect 9036 38150 9088 38156
rect 9048 38010 9076 38150
rect 8668 38004 8720 38010
rect 8668 37946 8720 37952
rect 9036 38004 9088 38010
rect 9036 37946 9088 37952
rect 8392 37868 8444 37874
rect 8392 37810 8444 37816
rect 8404 37262 8432 37810
rect 8668 37732 8720 37738
rect 8668 37674 8720 37680
rect 8680 37466 8708 37674
rect 8668 37460 8720 37466
rect 8668 37402 8720 37408
rect 8392 37256 8444 37262
rect 8392 37198 8444 37204
rect 8680 36854 8708 37402
rect 8760 37120 8812 37126
rect 8760 37062 8812 37068
rect 8944 37120 8996 37126
rect 8944 37062 8996 37068
rect 8668 36848 8720 36854
rect 8668 36790 8720 36796
rect 8392 36712 8444 36718
rect 8392 36654 8444 36660
rect 8208 36576 8260 36582
rect 8208 36518 8260 36524
rect 8220 36378 8248 36518
rect 8404 36378 8432 36654
rect 8208 36372 8260 36378
rect 8208 36314 8260 36320
rect 8392 36372 8444 36378
rect 8392 36314 8444 36320
rect 8772 36242 8800 37062
rect 8956 36378 8984 37062
rect 9140 36938 9168 39238
rect 9496 38344 9548 38350
rect 9496 38286 9548 38292
rect 9140 36910 9260 36938
rect 8944 36372 8996 36378
rect 8944 36314 8996 36320
rect 8760 36236 8812 36242
rect 8760 36178 8812 36184
rect 8392 36168 8444 36174
rect 8392 36110 8444 36116
rect 8208 35624 8260 35630
rect 8208 35566 8260 35572
rect 7472 33584 7524 33590
rect 7472 33526 7524 33532
rect 7748 33584 7800 33590
rect 7748 33526 7800 33532
rect 7104 33312 7156 33318
rect 7104 33254 7156 33260
rect 7116 32910 7144 33254
rect 7104 32904 7156 32910
rect 7104 32846 7156 32852
rect 7208 32830 7420 32858
rect 7208 32212 7236 32830
rect 7392 32774 7420 32830
rect 7288 32768 7340 32774
rect 7288 32710 7340 32716
rect 7380 32768 7432 32774
rect 7380 32710 7432 32716
rect 7300 32570 7328 32710
rect 7484 32570 7512 33526
rect 7564 33516 7616 33522
rect 7564 33458 7616 33464
rect 7840 33516 7892 33522
rect 7840 33458 7892 33464
rect 7576 33114 7604 33458
rect 7564 33108 7616 33114
rect 7564 33050 7616 33056
rect 7852 32910 7880 33458
rect 7840 32904 7892 32910
rect 7840 32846 7892 32852
rect 7288 32564 7340 32570
rect 7288 32506 7340 32512
rect 7472 32564 7524 32570
rect 7472 32506 7524 32512
rect 7116 32184 7236 32212
rect 7840 32224 7892 32230
rect 7116 31346 7144 32184
rect 7840 32166 7892 32172
rect 7852 32026 7880 32166
rect 7840 32020 7892 32026
rect 7840 31962 7892 31968
rect 7196 31748 7248 31754
rect 7196 31690 7248 31696
rect 7104 31340 7156 31346
rect 7104 31282 7156 31288
rect 7012 30932 7064 30938
rect 7012 30874 7064 30880
rect 6828 30320 6880 30326
rect 6828 30262 6880 30268
rect 6644 30252 6696 30258
rect 6644 30194 6696 30200
rect 6656 29850 6684 30194
rect 6644 29844 6696 29850
rect 6644 29786 6696 29792
rect 6736 29844 6788 29850
rect 6736 29786 6788 29792
rect 6748 29714 6776 29786
rect 6736 29708 6788 29714
rect 6736 29650 6788 29656
rect 6840 29594 6868 30262
rect 6564 29578 6868 29594
rect 6552 29572 6868 29578
rect 6604 29566 6868 29572
rect 6552 29514 6604 29520
rect 6736 29504 6788 29510
rect 6736 29446 6788 29452
rect 6920 29504 6972 29510
rect 6920 29446 6972 29452
rect 6748 29306 6776 29446
rect 6460 29300 6512 29306
rect 6460 29242 6512 29248
rect 6736 29300 6788 29306
rect 6736 29242 6788 29248
rect 6368 28212 6420 28218
rect 6368 28154 6420 28160
rect 6092 27872 6144 27878
rect 6092 27814 6144 27820
rect 5632 27464 5684 27470
rect 5632 27406 5684 27412
rect 5264 27396 5316 27402
rect 5264 27338 5316 27344
rect 5172 27328 5224 27334
rect 5172 27270 5224 27276
rect 5184 27062 5212 27270
rect 5172 27056 5224 27062
rect 5172 26998 5224 27004
rect 5080 26852 5132 26858
rect 5080 26794 5132 26800
rect 5172 26376 5224 26382
rect 5172 26318 5224 26324
rect 4804 26240 4856 26246
rect 4804 26182 4856 26188
rect 4816 25294 4844 26182
rect 5184 25294 5212 26318
rect 4068 25288 4120 25294
rect 4068 25230 4120 25236
rect 4712 25288 4764 25294
rect 4712 25230 4764 25236
rect 4804 25288 4856 25294
rect 4804 25230 4856 25236
rect 5172 25288 5224 25294
rect 5172 25230 5224 25236
rect 4080 23730 4108 25230
rect 4712 25152 4764 25158
rect 4712 25094 4764 25100
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4724 24206 4752 25094
rect 4896 24336 4948 24342
rect 4896 24278 4948 24284
rect 4344 24200 4396 24206
rect 4344 24142 4396 24148
rect 4712 24200 4764 24206
rect 4712 24142 4764 24148
rect 4356 23866 4384 24142
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4344 23860 4396 23866
rect 4344 23802 4396 23808
rect 3976 23724 4028 23730
rect 3976 23666 4028 23672
rect 4068 23724 4120 23730
rect 4068 23666 4120 23672
rect 3884 23656 3936 23662
rect 3884 23598 3936 23604
rect 3896 23118 3924 23598
rect 3988 23236 4016 23666
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23322 4660 24006
rect 4908 23866 4936 24278
rect 5276 24138 5304 27338
rect 6104 26994 6132 27814
rect 6276 27328 6328 27334
rect 6276 27270 6328 27276
rect 6288 27062 6316 27270
rect 6380 27062 6408 28154
rect 6472 27470 6500 29242
rect 6748 28762 6776 29242
rect 6932 29238 6960 29446
rect 6920 29232 6972 29238
rect 6920 29174 6972 29180
rect 6828 29096 6880 29102
rect 6828 29038 6880 29044
rect 6840 28762 6868 29038
rect 6736 28756 6788 28762
rect 6736 28698 6788 28704
rect 6828 28756 6880 28762
rect 6828 28698 6880 28704
rect 6552 28688 6604 28694
rect 6552 28630 6604 28636
rect 6564 27470 6592 28630
rect 6932 28558 6960 29174
rect 6920 28552 6972 28558
rect 6920 28494 6972 28500
rect 7116 28218 7144 31282
rect 7208 31142 7236 31690
rect 7196 31136 7248 31142
rect 7196 31078 7248 31084
rect 8220 30802 8248 35566
rect 8300 35012 8352 35018
rect 8300 34954 8352 34960
rect 8312 30938 8340 34954
rect 8404 31482 8432 36110
rect 8484 36032 8536 36038
rect 8484 35974 8536 35980
rect 8496 35086 8524 35974
rect 8772 35086 8800 36178
rect 8852 35624 8904 35630
rect 8852 35566 8904 35572
rect 8864 35290 8892 35566
rect 8852 35284 8904 35290
rect 8852 35226 8904 35232
rect 8484 35080 8536 35086
rect 8484 35022 8536 35028
rect 8760 35080 8812 35086
rect 8760 35022 8812 35028
rect 9128 35012 9180 35018
rect 9128 34954 9180 34960
rect 9036 33584 9088 33590
rect 9036 33526 9088 33532
rect 8576 32564 8628 32570
rect 8576 32506 8628 32512
rect 8392 31476 8444 31482
rect 8392 31418 8444 31424
rect 8484 31340 8536 31346
rect 8484 31282 8536 31288
rect 8496 31142 8524 31282
rect 8484 31136 8536 31142
rect 8484 31078 8536 31084
rect 8300 30932 8352 30938
rect 8300 30874 8352 30880
rect 8208 30796 8260 30802
rect 8208 30738 8260 30744
rect 7472 30728 7524 30734
rect 7472 30670 7524 30676
rect 7484 30054 7512 30670
rect 7472 30048 7524 30054
rect 7472 29990 7524 29996
rect 7484 29510 7512 29990
rect 7472 29504 7524 29510
rect 7472 29446 7524 29452
rect 7196 29028 7248 29034
rect 7196 28970 7248 28976
rect 7208 28558 7236 28970
rect 7288 28756 7340 28762
rect 7288 28698 7340 28704
rect 7196 28552 7248 28558
rect 7196 28494 7248 28500
rect 7104 28212 7156 28218
rect 7104 28154 7156 28160
rect 6828 27532 6880 27538
rect 6828 27474 6880 27480
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 6552 27464 6604 27470
rect 6552 27406 6604 27412
rect 6736 27328 6788 27334
rect 6736 27270 6788 27276
rect 6276 27056 6328 27062
rect 6276 26998 6328 27004
rect 6368 27056 6420 27062
rect 6368 26998 6420 27004
rect 5632 26988 5684 26994
rect 5632 26930 5684 26936
rect 6092 26988 6144 26994
rect 6092 26930 6144 26936
rect 5448 26308 5500 26314
rect 5448 26250 5500 26256
rect 5460 26042 5488 26250
rect 5448 26036 5500 26042
rect 5448 25978 5500 25984
rect 5644 25945 5672 26930
rect 5816 26784 5868 26790
rect 5816 26726 5868 26732
rect 5724 26580 5776 26586
rect 5724 26522 5776 26528
rect 5630 25936 5686 25945
rect 5630 25871 5686 25880
rect 5736 25498 5764 26522
rect 5828 25498 5856 26726
rect 6104 26518 6132 26930
rect 6184 26784 6236 26790
rect 6184 26726 6236 26732
rect 6552 26784 6604 26790
rect 6552 26726 6604 26732
rect 6092 26512 6144 26518
rect 6092 26454 6144 26460
rect 5724 25492 5776 25498
rect 5724 25434 5776 25440
rect 5816 25492 5868 25498
rect 5816 25434 5868 25440
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5448 25152 5500 25158
rect 5448 25094 5500 25100
rect 5540 25152 5592 25158
rect 5540 25094 5592 25100
rect 5460 24886 5488 25094
rect 5448 24880 5500 24886
rect 5448 24822 5500 24828
rect 5264 24132 5316 24138
rect 5264 24074 5316 24080
rect 4896 23860 4948 23866
rect 4896 23802 4948 23808
rect 4712 23520 4764 23526
rect 4712 23462 4764 23468
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 4620 23316 4672 23322
rect 4620 23258 4672 23264
rect 3988 23208 4200 23236
rect 3884 23112 3936 23118
rect 3936 23060 4108 23066
rect 3884 23054 4108 23060
rect 3896 23038 4108 23054
rect 3976 22772 4028 22778
rect 3976 22714 4028 22720
rect 3792 22024 3844 22030
rect 3792 21966 3844 21972
rect 3804 21690 3832 21966
rect 3792 21684 3844 21690
rect 3792 21626 3844 21632
rect 3700 21480 3752 21486
rect 3700 21422 3752 21428
rect 3712 21146 3740 21422
rect 3700 21140 3752 21146
rect 3700 21082 3752 21088
rect 3148 20936 3200 20942
rect 3148 20878 3200 20884
rect 3516 20936 3568 20942
rect 3516 20878 3568 20884
rect 2872 20868 2924 20874
rect 2872 20810 2924 20816
rect 2688 20800 2740 20806
rect 2688 20742 2740 20748
rect 2700 20466 2728 20742
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2412 19440 2464 19446
rect 938 19408 994 19417
rect 2412 19382 2464 19388
rect 3160 19378 3188 20878
rect 3988 20466 4016 22714
rect 4080 22166 4108 23038
rect 4172 22778 4200 23208
rect 4724 23186 4752 23462
rect 4712 23180 4764 23186
rect 4712 23122 4764 23128
rect 4712 22976 4764 22982
rect 4712 22918 4764 22924
rect 4160 22772 4212 22778
rect 4160 22714 4212 22720
rect 4724 22642 4752 22918
rect 4712 22636 4764 22642
rect 4712 22578 4764 22584
rect 4816 22506 4844 23462
rect 5356 22568 5408 22574
rect 5356 22510 5408 22516
rect 4804 22500 4856 22506
rect 4804 22442 4856 22448
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 22160 4120 22166
rect 4068 22102 4120 22108
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3884 20324 3936 20330
rect 3884 20266 3936 20272
rect 3896 20058 3924 20266
rect 3884 20052 3936 20058
rect 3884 19994 3936 20000
rect 3516 19712 3568 19718
rect 3516 19654 3568 19660
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3528 19378 3556 19654
rect 938 19343 994 19352
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2884 18970 2912 19246
rect 2872 18964 2924 18970
rect 2872 18906 2924 18912
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 1584 18216 1636 18222
rect 1584 18158 1636 18164
rect 1596 17921 1624 18158
rect 1582 17912 1638 17921
rect 1582 17847 1638 17856
rect 2240 17542 2268 18702
rect 2504 18352 2556 18358
rect 2504 18294 2556 18300
rect 2412 17604 2464 17610
rect 2412 17546 2464 17552
rect 2228 17536 2280 17542
rect 2228 17478 2280 17484
rect 2240 17202 2268 17478
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2424 16454 2452 17546
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 2412 16448 2464 16454
rect 2412 16390 2464 16396
rect 938 16144 994 16153
rect 938 16079 940 16088
rect 992 16079 994 16088
rect 940 16050 992 16056
rect 1688 16046 1716 16390
rect 1676 16040 1728 16046
rect 1676 15982 1728 15988
rect 940 14952 992 14958
rect 940 14894 992 14900
rect 952 14521 980 14894
rect 938 14512 994 14521
rect 938 14447 994 14456
rect 940 13252 992 13258
rect 940 13194 992 13200
rect 952 12889 980 13194
rect 938 12880 994 12889
rect 938 12815 994 12824
rect 940 11688 992 11694
rect 940 11630 992 11636
rect 952 11257 980 11630
rect 938 11248 994 11257
rect 938 11183 994 11192
rect 1584 9988 1636 9994
rect 1584 9930 1636 9936
rect 1596 9625 1624 9930
rect 1582 9616 1638 9625
rect 1582 9551 1638 9560
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1596 8265 1624 8366
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 2516 6914 2544 18294
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 2700 17882 2728 18226
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2688 17876 2740 17882
rect 2688 17818 2740 17824
rect 2884 17746 2912 18022
rect 2872 17740 2924 17746
rect 2872 17682 2924 17688
rect 3160 17678 3188 19314
rect 3240 19168 3292 19174
rect 3240 19110 3292 19116
rect 3252 18834 3280 19110
rect 3804 18970 3832 19654
rect 3988 19334 4016 20402
rect 4080 19854 4108 22102
rect 4632 22094 4660 22374
rect 4816 22234 4844 22442
rect 4804 22228 4856 22234
rect 4804 22170 4856 22176
rect 4632 22066 4844 22094
rect 4436 21956 4488 21962
rect 4436 21898 4488 21904
rect 4448 21486 4476 21898
rect 4816 21554 4844 22066
rect 5368 22030 5396 22510
rect 5356 22024 5408 22030
rect 5356 21966 5408 21972
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4804 21548 4856 21554
rect 4804 21490 4856 21496
rect 4436 21480 4488 21486
rect 4436 21422 4488 21428
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4724 21146 4752 21490
rect 4712 21140 4764 21146
rect 4712 21082 4764 21088
rect 4344 20936 4396 20942
rect 4344 20878 4396 20884
rect 4356 20602 4384 20878
rect 4620 20868 4672 20874
rect 4620 20810 4672 20816
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 4632 20398 4660 20810
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4620 20256 4672 20262
rect 4620 20198 4672 20204
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 4172 19854 4200 19994
rect 4632 19922 4660 20198
rect 4620 19916 4672 19922
rect 4620 19858 4672 19864
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 4160 19848 4212 19854
rect 4160 19790 4212 19796
rect 4528 19848 4580 19854
rect 4724 19802 4752 21082
rect 5368 20942 5396 21966
rect 5356 20936 5408 20942
rect 5356 20878 5408 20884
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 5092 20058 5120 20402
rect 5080 20052 5132 20058
rect 5080 19994 5132 20000
rect 4580 19796 4752 19802
rect 4528 19790 4752 19796
rect 4540 19774 4752 19790
rect 4620 19712 4672 19718
rect 4620 19654 4672 19660
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 3988 19306 4108 19334
rect 4080 19174 4108 19306
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 3792 18964 3844 18970
rect 3792 18906 3844 18912
rect 3240 18828 3292 18834
rect 3240 18770 3292 18776
rect 4080 18766 4108 19110
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 3620 18426 3648 18702
rect 3792 18624 3844 18630
rect 3792 18566 3844 18572
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3516 18216 3568 18222
rect 3516 18158 3568 18164
rect 3528 17882 3556 18158
rect 3804 17882 3832 18566
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3792 17876 3844 17882
rect 3792 17818 3844 17824
rect 4080 17678 4108 18702
rect 4528 18624 4580 18630
rect 4528 18566 4580 18572
rect 4540 18358 4568 18566
rect 4528 18352 4580 18358
rect 4528 18294 4580 18300
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17882 4660 19654
rect 4724 18902 4752 19654
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4712 18896 4764 18902
rect 4712 18838 4764 18844
rect 4712 18080 4764 18086
rect 4712 18022 4764 18028
rect 4620 17876 4672 17882
rect 4620 17818 4672 17824
rect 4724 17814 4752 18022
rect 4712 17808 4764 17814
rect 4712 17750 4764 17756
rect 3148 17672 3200 17678
rect 4068 17672 4120 17678
rect 3148 17614 3200 17620
rect 3988 17620 4068 17626
rect 3988 17614 4120 17620
rect 3160 16658 3188 17614
rect 3988 17598 4108 17614
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3436 16794 3464 16934
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 3988 16590 4016 17598
rect 4160 17128 4212 17134
rect 4080 17076 4160 17082
rect 4080 17070 4212 17076
rect 4080 17054 4200 17070
rect 4080 16590 4108 17054
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 4068 16584 4120 16590
rect 4068 16526 4120 16532
rect 3804 16250 3832 16526
rect 4528 16448 4580 16454
rect 4580 16408 4660 16436
rect 4528 16390 4580 16396
rect 3792 16244 3844 16250
rect 3792 16186 3844 16192
rect 4632 16046 4660 16408
rect 4724 16114 4752 17750
rect 4816 16998 4844 18906
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4908 17882 4936 18770
rect 5368 18340 5396 19382
rect 5448 18352 5500 18358
rect 5368 18312 5448 18340
rect 4896 17876 4948 17882
rect 4896 17818 4948 17824
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 5368 16522 5396 18312
rect 5448 18294 5500 18300
rect 5552 17338 5580 25094
rect 5644 22030 5672 25230
rect 5736 24954 5764 25434
rect 5724 24948 5776 24954
rect 5724 24890 5776 24896
rect 5736 24206 5764 24890
rect 5724 24200 5776 24206
rect 5724 24142 5776 24148
rect 5724 22160 5776 22166
rect 5724 22102 5776 22108
rect 5632 22024 5684 22030
rect 5632 21966 5684 21972
rect 5736 21622 5764 22102
rect 6000 22024 6052 22030
rect 6000 21966 6052 21972
rect 5724 21616 5776 21622
rect 5724 21558 5776 21564
rect 6012 21554 6040 21966
rect 6000 21548 6052 21554
rect 6000 21490 6052 21496
rect 5908 20460 5960 20466
rect 5908 20402 5960 20408
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5828 20058 5856 20198
rect 5816 20052 5868 20058
rect 5816 19994 5868 20000
rect 5920 19990 5948 20402
rect 5908 19984 5960 19990
rect 5908 19926 5960 19932
rect 5908 18624 5960 18630
rect 5908 18566 5960 18572
rect 5920 18222 5948 18566
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 6196 17338 6224 26726
rect 6564 26586 6592 26726
rect 6552 26580 6604 26586
rect 6552 26522 6604 26528
rect 6748 24410 6776 27270
rect 6736 24404 6788 24410
rect 6736 24346 6788 24352
rect 6552 24200 6604 24206
rect 6552 24142 6604 24148
rect 6368 24064 6420 24070
rect 6368 24006 6420 24012
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6288 19922 6316 20198
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 6380 18766 6408 24006
rect 6564 23118 6592 24142
rect 6840 23322 6868 27474
rect 7300 27112 7328 28698
rect 7484 27470 7512 29446
rect 8588 28994 8616 32506
rect 8852 32428 8904 32434
rect 8852 32370 8904 32376
rect 8760 31340 8812 31346
rect 8760 31282 8812 31288
rect 8772 31142 8800 31282
rect 8864 31210 8892 32370
rect 9048 31414 9076 33526
rect 9036 31408 9088 31414
rect 9036 31350 9088 31356
rect 8852 31204 8904 31210
rect 8852 31146 8904 31152
rect 8760 31136 8812 31142
rect 8760 31078 8812 31084
rect 8944 31136 8996 31142
rect 8944 31078 8996 31084
rect 8956 30734 8984 31078
rect 8944 30728 8996 30734
rect 8944 30670 8996 30676
rect 9140 29714 9168 34954
rect 9232 30938 9260 36910
rect 9508 36854 9536 38286
rect 9496 36848 9548 36854
rect 9496 36790 9548 36796
rect 9864 34536 9916 34542
rect 9864 34478 9916 34484
rect 9312 33992 9364 33998
rect 9312 33934 9364 33940
rect 9324 33658 9352 33934
rect 9404 33924 9456 33930
rect 9404 33866 9456 33872
rect 9312 33652 9364 33658
rect 9312 33594 9364 33600
rect 9312 33516 9364 33522
rect 9312 33458 9364 33464
rect 9324 32570 9352 33458
rect 9416 33386 9444 33866
rect 9876 33862 9904 34478
rect 9772 33856 9824 33862
rect 9772 33798 9824 33804
rect 9864 33856 9916 33862
rect 9864 33798 9916 33804
rect 9404 33380 9456 33386
rect 9404 33322 9456 33328
rect 9784 33318 9812 33798
rect 9876 33658 9904 33798
rect 9864 33652 9916 33658
rect 9864 33594 9916 33600
rect 9772 33312 9824 33318
rect 9772 33254 9824 33260
rect 9312 32564 9364 32570
rect 9312 32506 9364 32512
rect 10152 31686 10180 39918
rect 11704 39840 11756 39846
rect 11704 39782 11756 39788
rect 10232 38752 10284 38758
rect 10232 38694 10284 38700
rect 10244 38282 10272 38694
rect 10508 38412 10560 38418
rect 10508 38354 10560 38360
rect 10232 38276 10284 38282
rect 10232 38218 10284 38224
rect 10520 36786 10548 38354
rect 10508 36780 10560 36786
rect 10508 36722 10560 36728
rect 10232 36712 10284 36718
rect 10232 36654 10284 36660
rect 10244 36378 10272 36654
rect 10232 36372 10284 36378
rect 10232 36314 10284 36320
rect 10520 35698 10548 36722
rect 10508 35692 10560 35698
rect 10508 35634 10560 35640
rect 10324 33380 10376 33386
rect 10324 33322 10376 33328
rect 10336 32502 10364 33322
rect 10416 33312 10468 33318
rect 10416 33254 10468 33260
rect 10324 32496 10376 32502
rect 10324 32438 10376 32444
rect 10232 32360 10284 32366
rect 10232 32302 10284 32308
rect 10244 32026 10272 32302
rect 10232 32020 10284 32026
rect 10232 31962 10284 31968
rect 10428 31754 10456 33254
rect 10600 31816 10652 31822
rect 10600 31758 10652 31764
rect 10416 31748 10468 31754
rect 10416 31690 10468 31696
rect 10140 31680 10192 31686
rect 10140 31622 10192 31628
rect 10048 31408 10100 31414
rect 10048 31350 10100 31356
rect 9680 31136 9732 31142
rect 9680 31078 9732 31084
rect 9220 30932 9272 30938
rect 9220 30874 9272 30880
rect 9692 30870 9720 31078
rect 9680 30864 9732 30870
rect 9680 30806 9732 30812
rect 10060 30666 10088 31350
rect 10152 30938 10180 31622
rect 10612 30954 10640 31758
rect 11716 31754 11744 39782
rect 12440 32496 12492 32502
rect 12440 32438 12492 32444
rect 12348 32224 12400 32230
rect 12348 32166 12400 32172
rect 11716 31726 11836 31754
rect 11704 31680 11756 31686
rect 11704 31622 11756 31628
rect 10968 31340 11020 31346
rect 10968 31282 11020 31288
rect 11520 31340 11572 31346
rect 11520 31282 11572 31288
rect 10140 30932 10192 30938
rect 10140 30874 10192 30880
rect 10428 30926 10640 30954
rect 9772 30660 9824 30666
rect 9772 30602 9824 30608
rect 10048 30660 10100 30666
rect 10048 30602 10100 30608
rect 9312 30592 9364 30598
rect 9312 30534 9364 30540
rect 9220 30048 9272 30054
rect 9220 29990 9272 29996
rect 9128 29708 9180 29714
rect 9128 29650 9180 29656
rect 8944 29640 8996 29646
rect 8944 29582 8996 29588
rect 8956 29306 8984 29582
rect 8944 29300 8996 29306
rect 8944 29242 8996 29248
rect 8588 28966 8800 28994
rect 8392 28484 8444 28490
rect 8392 28426 8444 28432
rect 8404 28150 8432 28426
rect 8772 28218 8800 28966
rect 9128 28416 9180 28422
rect 9128 28358 9180 28364
rect 9140 28218 9168 28358
rect 8760 28212 8812 28218
rect 8760 28154 8812 28160
rect 9128 28212 9180 28218
rect 9128 28154 9180 28160
rect 8392 28144 8444 28150
rect 8392 28086 8444 28092
rect 7656 27872 7708 27878
rect 7656 27814 7708 27820
rect 7472 27464 7524 27470
rect 7472 27406 7524 27412
rect 7668 27402 7696 27814
rect 8404 27538 8432 28086
rect 8484 28076 8536 28082
rect 8484 28018 8536 28024
rect 8392 27532 8444 27538
rect 8392 27474 8444 27480
rect 7656 27396 7708 27402
rect 7656 27338 7708 27344
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 7300 27084 7420 27112
rect 7196 26988 7248 26994
rect 7248 26948 7328 26976
rect 7196 26930 7248 26936
rect 7104 26784 7156 26790
rect 7104 26726 7156 26732
rect 7116 26450 7144 26726
rect 7104 26444 7156 26450
rect 7104 26386 7156 26392
rect 7196 25696 7248 25702
rect 7196 25638 7248 25644
rect 7208 25294 7236 25638
rect 7300 25430 7328 26948
rect 7288 25424 7340 25430
rect 7288 25366 7340 25372
rect 7196 25288 7248 25294
rect 7196 25230 7248 25236
rect 7288 25288 7340 25294
rect 7392 25242 7420 27084
rect 7472 27056 7524 27062
rect 7472 26998 7524 27004
rect 7484 26450 7512 26998
rect 8220 26994 8248 27270
rect 7840 26988 7892 26994
rect 7840 26930 7892 26936
rect 8208 26988 8260 26994
rect 8208 26930 8260 26936
rect 7852 26586 7880 26930
rect 7840 26580 7892 26586
rect 7840 26522 7892 26528
rect 7472 26444 7524 26450
rect 7472 26386 7524 26392
rect 8392 26444 8444 26450
rect 8392 26386 8444 26392
rect 7564 26308 7616 26314
rect 7564 26250 7616 26256
rect 7472 25696 7524 25702
rect 7472 25638 7524 25644
rect 7484 25498 7512 25638
rect 7472 25492 7524 25498
rect 7472 25434 7524 25440
rect 7340 25236 7420 25242
rect 7288 25230 7420 25236
rect 7300 25214 7420 25230
rect 7300 24750 7328 25214
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7012 24200 7064 24206
rect 7012 24142 7064 24148
rect 7024 23526 7052 24142
rect 7300 23866 7328 24686
rect 7380 24200 7432 24206
rect 7380 24142 7432 24148
rect 7288 23860 7340 23866
rect 7288 23802 7340 23808
rect 7012 23520 7064 23526
rect 7012 23462 7064 23468
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 7024 23118 7052 23462
rect 6552 23112 6604 23118
rect 6552 23054 6604 23060
rect 7012 23112 7064 23118
rect 7012 23054 7064 23060
rect 6644 22976 6696 22982
rect 6644 22918 6696 22924
rect 6656 22094 6684 22918
rect 7012 22568 7064 22574
rect 7012 22510 7064 22516
rect 6564 22066 6684 22094
rect 6460 21548 6512 21554
rect 6460 21490 6512 21496
rect 6472 21146 6500 21490
rect 6460 21140 6512 21146
rect 6460 21082 6512 21088
rect 6472 20602 6500 21082
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 6564 19666 6592 22066
rect 6644 21956 6696 21962
rect 6644 21898 6696 21904
rect 6656 21690 6684 21898
rect 7024 21690 7052 22510
rect 7300 22094 7328 23802
rect 7392 23322 7420 24142
rect 7576 24138 7604 26250
rect 7748 26240 7800 26246
rect 7748 26182 7800 26188
rect 7760 26042 7788 26182
rect 7748 26036 7800 26042
rect 7748 25978 7800 25984
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 7852 24682 7880 25842
rect 7932 25288 7984 25294
rect 7932 25230 7984 25236
rect 7840 24676 7892 24682
rect 7840 24618 7892 24624
rect 7656 24336 7708 24342
rect 7656 24278 7708 24284
rect 7564 24132 7616 24138
rect 7564 24074 7616 24080
rect 7380 23316 7432 23322
rect 7380 23258 7432 23264
rect 7380 22636 7432 22642
rect 7380 22578 7432 22584
rect 7392 22234 7420 22578
rect 7380 22228 7432 22234
rect 7380 22170 7432 22176
rect 7116 22066 7328 22094
rect 6644 21684 6696 21690
rect 6644 21626 6696 21632
rect 7012 21684 7064 21690
rect 7012 21626 7064 21632
rect 7024 21554 7052 21626
rect 7012 21548 7064 21554
rect 7012 21490 7064 21496
rect 6920 20868 6972 20874
rect 6920 20810 6972 20816
rect 6932 20602 6960 20810
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6736 20256 6788 20262
rect 6736 20198 6788 20204
rect 6748 19854 6776 20198
rect 7116 20058 7144 22066
rect 7576 21622 7604 24074
rect 7668 23866 7696 24278
rect 7852 24138 7880 24618
rect 7840 24132 7892 24138
rect 7840 24074 7892 24080
rect 7944 23866 7972 25230
rect 8024 25220 8076 25226
rect 8024 25162 8076 25168
rect 7656 23860 7708 23866
rect 7932 23860 7984 23866
rect 7656 23802 7708 23808
rect 7852 23820 7932 23848
rect 7852 23118 7880 23820
rect 7932 23802 7984 23808
rect 7932 23520 7984 23526
rect 7932 23462 7984 23468
rect 7944 23322 7972 23462
rect 7932 23316 7984 23322
rect 7932 23258 7984 23264
rect 7840 23112 7892 23118
rect 7840 23054 7892 23060
rect 8036 22778 8064 25162
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 8312 24206 8340 25094
rect 8208 24200 8260 24206
rect 8208 24142 8260 24148
rect 8300 24200 8352 24206
rect 8300 24142 8352 24148
rect 8220 23866 8248 24142
rect 8208 23860 8260 23866
rect 8208 23802 8260 23808
rect 8116 23656 8168 23662
rect 8116 23598 8168 23604
rect 8128 23322 8156 23598
rect 8116 23316 8168 23322
rect 8116 23258 8168 23264
rect 8404 23118 8432 26386
rect 8496 26024 8524 28018
rect 8668 28008 8720 28014
rect 8944 28008 8996 28014
rect 8720 27968 8944 27996
rect 8668 27950 8720 27956
rect 8944 27950 8996 27956
rect 8852 27532 8904 27538
rect 8852 27474 8904 27480
rect 8496 25996 8708 26024
rect 8680 25906 8708 25996
rect 8484 25900 8536 25906
rect 8484 25842 8536 25848
rect 8576 25900 8628 25906
rect 8576 25842 8628 25848
rect 8668 25900 8720 25906
rect 8668 25842 8720 25848
rect 8496 25294 8524 25842
rect 8588 25362 8616 25842
rect 8760 25696 8812 25702
rect 8760 25638 8812 25644
rect 8772 25498 8800 25638
rect 8760 25492 8812 25498
rect 8760 25434 8812 25440
rect 8576 25356 8628 25362
rect 8576 25298 8628 25304
rect 8484 25288 8536 25294
rect 8484 25230 8536 25236
rect 8864 25226 8892 27474
rect 9232 26518 9260 29990
rect 9324 28966 9352 30534
rect 9784 29646 9812 30602
rect 9864 30592 9916 30598
rect 9864 30534 9916 30540
rect 9956 30592 10008 30598
rect 9956 30534 10008 30540
rect 9876 30394 9904 30534
rect 9864 30388 9916 30394
rect 9864 30330 9916 30336
rect 9772 29640 9824 29646
rect 9772 29582 9824 29588
rect 9312 28960 9364 28966
rect 9312 28902 9364 28908
rect 9324 28422 9352 28902
rect 9312 28416 9364 28422
rect 9312 28358 9364 28364
rect 9220 26512 9272 26518
rect 9220 26454 9272 26460
rect 9034 25936 9090 25945
rect 9034 25871 9036 25880
rect 9088 25871 9090 25880
rect 9036 25842 9088 25848
rect 8852 25220 8904 25226
rect 8852 25162 8904 25168
rect 8484 24336 8536 24342
rect 8484 24278 8536 24284
rect 8496 23866 8524 24278
rect 8484 23860 8536 23866
rect 8484 23802 8536 23808
rect 8392 23112 8444 23118
rect 8392 23054 8444 23060
rect 8404 22778 8432 23054
rect 8024 22772 8076 22778
rect 8024 22714 8076 22720
rect 8392 22772 8444 22778
rect 8392 22714 8444 22720
rect 8036 22522 8064 22714
rect 8036 22494 8156 22522
rect 8024 22432 8076 22438
rect 8024 22374 8076 22380
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 8036 21536 8064 22374
rect 8128 22094 8156 22494
rect 8576 22432 8628 22438
rect 8576 22374 8628 22380
rect 8588 22234 8616 22374
rect 8576 22228 8628 22234
rect 8576 22170 8628 22176
rect 8128 22066 8340 22094
rect 8208 21956 8260 21962
rect 8208 21898 8260 21904
rect 8220 21690 8248 21898
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8208 21548 8260 21554
rect 8036 21508 8208 21536
rect 8208 21490 8260 21496
rect 8312 21434 8340 22066
rect 8116 21412 8168 21418
rect 8116 21354 8168 21360
rect 8220 21406 8340 21434
rect 8128 21146 8156 21354
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 8024 20868 8076 20874
rect 8024 20810 8076 20816
rect 8036 20262 8064 20810
rect 8128 20602 8156 21082
rect 8220 20602 8248 21406
rect 8864 20874 8892 25162
rect 8576 20868 8628 20874
rect 8576 20810 8628 20816
rect 8852 20868 8904 20874
rect 8852 20810 8904 20816
rect 8116 20596 8168 20602
rect 8116 20538 8168 20544
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8588 20534 8616 20810
rect 8576 20528 8628 20534
rect 8576 20470 8628 20476
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 7932 20256 7984 20262
rect 7932 20198 7984 20204
rect 8024 20256 8076 20262
rect 8024 20198 8076 20204
rect 7104 20052 7156 20058
rect 7104 19994 7156 20000
rect 7944 19854 7972 20198
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 7932 19848 7984 19854
rect 7932 19790 7984 19796
rect 8312 19786 8340 20402
rect 8300 19780 8352 19786
rect 8300 19722 8352 19728
rect 6472 19638 6592 19666
rect 6368 18760 6420 18766
rect 6368 18702 6420 18708
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 5540 17332 5592 17338
rect 5540 17274 5592 17280
rect 6184 17332 6236 17338
rect 6184 17274 6236 17280
rect 6184 17128 6236 17134
rect 6184 17070 6236 17076
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5460 16794 5488 16934
rect 6196 16794 6224 17070
rect 5448 16788 5500 16794
rect 5448 16730 5500 16736
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6288 16658 6316 18158
rect 6472 17202 6500 19638
rect 8864 19514 8892 20810
rect 9048 20262 9076 25842
rect 9128 25696 9180 25702
rect 9128 25638 9180 25644
rect 9140 25430 9168 25638
rect 9128 25424 9180 25430
rect 9128 25366 9180 25372
rect 9232 22642 9260 26454
rect 9324 22710 9352 28358
rect 9784 26994 9812 29582
rect 9968 29578 9996 30534
rect 9956 29572 10008 29578
rect 9956 29514 10008 29520
rect 9968 29238 9996 29514
rect 9956 29232 10008 29238
rect 9956 29174 10008 29180
rect 9864 28688 9916 28694
rect 9864 28630 9916 28636
rect 9876 28082 9904 28630
rect 9968 28558 9996 29174
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 9864 28076 9916 28082
rect 9864 28018 9916 28024
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 9680 26580 9732 26586
rect 9680 26522 9732 26528
rect 9692 26042 9720 26522
rect 9680 26036 9732 26042
rect 9680 25978 9732 25984
rect 9692 25362 9720 25978
rect 9772 25968 9824 25974
rect 9772 25910 9824 25916
rect 9784 25498 9812 25910
rect 9772 25492 9824 25498
rect 9772 25434 9824 25440
rect 9680 25356 9732 25362
rect 9680 25298 9732 25304
rect 9876 25226 9904 28018
rect 9968 27130 9996 28494
rect 9956 27124 10008 27130
rect 9956 27066 10008 27072
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9864 25220 9916 25226
rect 9864 25162 9916 25168
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9692 24410 9720 24550
rect 9968 24410 9996 26726
rect 10060 24886 10088 30602
rect 10324 30592 10376 30598
rect 10324 30534 10376 30540
rect 10336 30394 10364 30534
rect 10324 30388 10376 30394
rect 10324 30330 10376 30336
rect 10428 30122 10456 30926
rect 10600 30592 10652 30598
rect 10600 30534 10652 30540
rect 10612 30326 10640 30534
rect 10980 30326 11008 31282
rect 11060 30388 11112 30394
rect 11060 30330 11112 30336
rect 10600 30320 10652 30326
rect 10600 30262 10652 30268
rect 10968 30320 11020 30326
rect 10968 30262 11020 30268
rect 10692 30252 10744 30258
rect 10692 30194 10744 30200
rect 10876 30242 10928 30248
rect 10416 30116 10468 30122
rect 10416 30058 10468 30064
rect 10232 29776 10284 29782
rect 10232 29718 10284 29724
rect 10244 28218 10272 29718
rect 10704 29458 10732 30194
rect 10876 30184 10928 30190
rect 10888 29646 10916 30184
rect 11072 30054 11100 30330
rect 11532 30190 11560 31282
rect 11716 30870 11744 31622
rect 11704 30864 11756 30870
rect 11704 30806 11756 30812
rect 11520 30184 11572 30190
rect 11520 30126 11572 30132
rect 11060 30048 11112 30054
rect 11060 29990 11112 29996
rect 10876 29640 10928 29646
rect 10876 29582 10928 29588
rect 11152 29504 11204 29510
rect 10704 29430 11100 29458
rect 11152 29446 11204 29452
rect 10704 29170 10732 29430
rect 11072 29238 11100 29430
rect 10968 29232 11020 29238
rect 10968 29174 11020 29180
rect 11060 29232 11112 29238
rect 11060 29174 11112 29180
rect 10508 29164 10560 29170
rect 10508 29106 10560 29112
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10692 29164 10744 29170
rect 10692 29106 10744 29112
rect 10520 28762 10548 29106
rect 10612 28994 10640 29106
rect 10980 28994 11008 29174
rect 11060 29096 11112 29102
rect 11164 29084 11192 29446
rect 11428 29232 11480 29238
rect 11428 29174 11480 29180
rect 11112 29056 11192 29084
rect 11060 29038 11112 29044
rect 10612 28966 11008 28994
rect 10612 28762 10640 28966
rect 10508 28756 10560 28762
rect 10508 28698 10560 28704
rect 10600 28756 10652 28762
rect 10600 28698 10652 28704
rect 11244 28756 11296 28762
rect 11244 28698 11296 28704
rect 11060 28552 11112 28558
rect 11060 28494 11112 28500
rect 10232 28212 10284 28218
rect 10232 28154 10284 28160
rect 10140 28008 10192 28014
rect 10140 27950 10192 27956
rect 10152 26586 10180 27950
rect 10244 27470 10272 28154
rect 11072 28014 11100 28494
rect 11060 28008 11112 28014
rect 11060 27950 11112 27956
rect 11256 27878 11284 28698
rect 11336 28552 11388 28558
rect 11336 28494 11388 28500
rect 11348 28150 11376 28494
rect 11336 28144 11388 28150
rect 11336 28086 11388 28092
rect 10324 27872 10376 27878
rect 10324 27814 10376 27820
rect 11244 27872 11296 27878
rect 11244 27814 11296 27820
rect 10232 27464 10284 27470
rect 10232 27406 10284 27412
rect 10140 26580 10192 26586
rect 10140 26522 10192 26528
rect 10336 26246 10364 27814
rect 11348 27674 11376 28086
rect 10968 27668 11020 27674
rect 10968 27610 11020 27616
rect 11336 27668 11388 27674
rect 11336 27610 11388 27616
rect 10416 27532 10468 27538
rect 10468 27492 10548 27520
rect 10416 27474 10468 27480
rect 10416 26988 10468 26994
rect 10416 26930 10468 26936
rect 10140 26240 10192 26246
rect 10140 26182 10192 26188
rect 10324 26240 10376 26246
rect 10324 26182 10376 26188
rect 10152 25702 10180 26182
rect 10336 25770 10364 26182
rect 10428 26042 10456 26930
rect 10520 26790 10548 27492
rect 10508 26784 10560 26790
rect 10508 26726 10560 26732
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10416 26036 10468 26042
rect 10416 25978 10468 25984
rect 10416 25900 10468 25906
rect 10416 25842 10468 25848
rect 10324 25764 10376 25770
rect 10324 25706 10376 25712
rect 10140 25696 10192 25702
rect 10140 25638 10192 25644
rect 10428 25498 10456 25842
rect 10416 25492 10468 25498
rect 10416 25434 10468 25440
rect 10232 25220 10284 25226
rect 10232 25162 10284 25168
rect 10048 24880 10100 24886
rect 10048 24822 10100 24828
rect 9680 24404 9732 24410
rect 9680 24346 9732 24352
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 9312 22704 9364 22710
rect 9312 22646 9364 22652
rect 9692 22642 9720 24346
rect 10048 24200 10100 24206
rect 10048 24142 10100 24148
rect 10140 24200 10192 24206
rect 10140 24142 10192 24148
rect 9772 24064 9824 24070
rect 9772 24006 9824 24012
rect 9220 22636 9272 22642
rect 9220 22578 9272 22584
rect 9680 22636 9732 22642
rect 9680 22578 9732 22584
rect 9232 22234 9260 22578
rect 9784 22522 9812 24006
rect 10060 23866 10088 24142
rect 10152 23866 10180 24142
rect 10048 23860 10100 23866
rect 10048 23802 10100 23808
rect 10140 23860 10192 23866
rect 10140 23802 10192 23808
rect 10140 23724 10192 23730
rect 10140 23666 10192 23672
rect 10152 23118 10180 23666
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 9968 22778 9996 23054
rect 10140 22976 10192 22982
rect 10140 22918 10192 22924
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 9600 22494 9812 22522
rect 9956 22568 10008 22574
rect 9956 22510 10008 22516
rect 9600 22250 9628 22494
rect 9680 22432 9732 22438
rect 9732 22392 9812 22420
rect 9680 22374 9732 22380
rect 9220 22228 9272 22234
rect 9600 22222 9720 22250
rect 9220 22170 9272 22176
rect 9036 20256 9088 20262
rect 9036 20198 9088 20204
rect 8852 19508 8904 19514
rect 8852 19450 8904 19456
rect 6828 19304 6880 19310
rect 6828 19246 6880 19252
rect 6840 18970 6868 19246
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 6828 18964 6880 18970
rect 6828 18906 6880 18912
rect 8404 18834 8432 19110
rect 6828 18828 6880 18834
rect 6828 18770 6880 18776
rect 8392 18828 8444 18834
rect 8392 18770 8444 18776
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6656 17610 6684 18702
rect 6840 18426 6868 18770
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 7024 18358 7052 18566
rect 8312 18358 8340 18566
rect 7012 18352 7064 18358
rect 7012 18294 7064 18300
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 6920 18284 6972 18290
rect 6920 18226 6972 18232
rect 6932 17678 6960 18226
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6644 17604 6696 17610
rect 6644 17546 6696 17552
rect 6656 17202 6684 17546
rect 6932 17270 6960 17614
rect 8680 17338 8708 17682
rect 9048 17610 9076 20198
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9324 19378 9352 19790
rect 9312 19372 9364 19378
rect 9312 19314 9364 19320
rect 9220 18080 9272 18086
rect 9220 18022 9272 18028
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 9232 17542 9260 18022
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 6460 17196 6512 17202
rect 6460 17138 6512 17144
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 6276 16652 6328 16658
rect 6276 16594 6328 16600
rect 6932 16590 6960 17206
rect 8116 17128 8168 17134
rect 8116 17070 8168 17076
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 7472 16992 7524 16998
rect 7472 16934 7524 16940
rect 7484 16794 7512 16934
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 5356 16516 5408 16522
rect 5356 16458 5408 16464
rect 6380 16250 6408 16526
rect 6736 16448 6788 16454
rect 6736 16390 6788 16396
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6748 16114 6776 16390
rect 6932 16250 6960 16526
rect 8128 16250 8156 17070
rect 9048 16454 9076 17070
rect 9036 16448 9088 16454
rect 9036 16390 9088 16396
rect 6920 16244 6972 16250
rect 6920 16186 6972 16192
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 2688 15904 2740 15910
rect 2688 15846 2740 15852
rect 2700 11762 2728 15846
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 2688 11756 2740 11762
rect 2688 11698 2740 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 2516 6886 2728 6914
rect 2700 6798 2728 6886
rect 2688 6792 2740 6798
rect 2688 6734 2740 6740
rect 940 6724 992 6730
rect 940 6666 992 6672
rect 952 6361 980 6666
rect 938 6352 994 6361
rect 938 6287 994 6296
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5234 4660 15982
rect 6748 13326 6776 16050
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 952 4729 980 5102
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 938 4720 994 4729
rect 938 4655 994 4664
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 9048 3534 9076 16390
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 940 3460 992 3466
rect 940 3402 992 3408
rect 952 3097 980 3402
rect 938 3088 994 3097
rect 938 3023 994 3032
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 9232 2378 9260 17478
rect 9324 8498 9352 19314
rect 9692 18290 9720 22222
rect 9784 21026 9812 22392
rect 9968 22234 9996 22510
rect 9956 22228 10008 22234
rect 9956 22170 10008 22176
rect 10152 22030 10180 22918
rect 10140 22024 10192 22030
rect 10140 21966 10192 21972
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9864 21412 9916 21418
rect 9864 21354 9916 21360
rect 9876 21146 9904 21354
rect 9968 21146 9996 21830
rect 10048 21344 10100 21350
rect 10048 21286 10100 21292
rect 10060 21146 10088 21286
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9956 21140 10008 21146
rect 9956 21082 10008 21088
rect 10048 21140 10100 21146
rect 10048 21082 10100 21088
rect 9784 20998 9904 21026
rect 9772 20868 9824 20874
rect 9772 20810 9824 20816
rect 9784 18834 9812 20810
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9680 18284 9732 18290
rect 9680 18226 9732 18232
rect 9784 16658 9812 18770
rect 9876 17882 9904 20998
rect 9956 20936 10008 20942
rect 10244 20890 10272 25162
rect 10324 25152 10376 25158
rect 10324 25094 10376 25100
rect 10336 24070 10364 25094
rect 10520 24290 10548 26726
rect 10612 26518 10640 26726
rect 10600 26512 10652 26518
rect 10600 26454 10652 26460
rect 10980 26382 11008 27610
rect 11244 27396 11296 27402
rect 11244 27338 11296 27344
rect 11336 27396 11388 27402
rect 11336 27338 11388 27344
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 10876 26308 10928 26314
rect 10876 26250 10928 26256
rect 10888 26042 10916 26250
rect 10980 26042 11008 26318
rect 10876 26036 10928 26042
rect 10876 25978 10928 25984
rect 10968 26036 11020 26042
rect 10968 25978 11020 25984
rect 11152 25900 11204 25906
rect 11152 25842 11204 25848
rect 11164 25702 11192 25842
rect 11152 25696 11204 25702
rect 11152 25638 11204 25644
rect 11164 25430 11192 25638
rect 11152 25424 11204 25430
rect 11152 25366 11204 25372
rect 10600 24608 10652 24614
rect 10600 24550 10652 24556
rect 10428 24262 10548 24290
rect 10324 24064 10376 24070
rect 10324 24006 10376 24012
rect 10336 22030 10364 24006
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10428 21146 10456 24262
rect 10508 24200 10560 24206
rect 10508 24142 10560 24148
rect 10520 23866 10548 24142
rect 10612 24070 10640 24550
rect 10600 24064 10652 24070
rect 10600 24006 10652 24012
rect 10508 23860 10560 23866
rect 10508 23802 10560 23808
rect 10612 21962 10640 24006
rect 10968 23724 11020 23730
rect 10968 23666 11020 23672
rect 10980 23526 11008 23666
rect 10968 23520 11020 23526
rect 10968 23462 11020 23468
rect 10784 22636 10836 22642
rect 10784 22578 10836 22584
rect 10796 22166 10824 22578
rect 10980 22438 11008 23462
rect 10968 22432 11020 22438
rect 10968 22374 11020 22380
rect 10980 22166 11008 22374
rect 10784 22160 10836 22166
rect 10784 22102 10836 22108
rect 10968 22160 11020 22166
rect 10968 22102 11020 22108
rect 10600 21956 10652 21962
rect 10600 21898 10652 21904
rect 10416 21140 10468 21146
rect 10416 21082 10468 21088
rect 9956 20878 10008 20884
rect 9968 18902 9996 20878
rect 10060 20862 10272 20890
rect 10060 20806 10088 20862
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 10140 20800 10192 20806
rect 10140 20742 10192 20748
rect 10060 20058 10088 20742
rect 10152 20398 10180 20742
rect 10140 20392 10192 20398
rect 10140 20334 10192 20340
rect 10324 20392 10376 20398
rect 10324 20334 10376 20340
rect 10048 20052 10100 20058
rect 10048 19994 10100 20000
rect 9956 18896 10008 18902
rect 9956 18838 10008 18844
rect 9968 18154 9996 18838
rect 9956 18148 10008 18154
rect 9956 18090 10008 18096
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9968 17678 9996 18090
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 10060 16794 10088 17478
rect 10048 16788 10100 16794
rect 10048 16730 10100 16736
rect 9772 16652 9824 16658
rect 9772 16594 9824 16600
rect 10152 15026 10180 20334
rect 10336 19446 10364 20334
rect 10612 20330 10640 21898
rect 10692 21480 10744 21486
rect 10692 21422 10744 21428
rect 10704 20602 10732 21422
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 10692 20596 10744 20602
rect 10692 20538 10744 20544
rect 10980 20398 11008 20810
rect 11256 20534 11284 27338
rect 11348 27130 11376 27338
rect 11336 27124 11388 27130
rect 11336 27066 11388 27072
rect 11336 26376 11388 26382
rect 11336 26318 11388 26324
rect 11348 25906 11376 26318
rect 11336 25900 11388 25906
rect 11336 25842 11388 25848
rect 11336 24744 11388 24750
rect 11336 24686 11388 24692
rect 11348 23866 11376 24686
rect 11440 24070 11468 29174
rect 11532 29034 11560 30126
rect 11612 29572 11664 29578
rect 11612 29514 11664 29520
rect 11624 29306 11652 29514
rect 11612 29300 11664 29306
rect 11612 29242 11664 29248
rect 11520 29028 11572 29034
rect 11520 28970 11572 28976
rect 11716 26994 11744 30806
rect 11520 26988 11572 26994
rect 11520 26930 11572 26936
rect 11704 26988 11756 26994
rect 11704 26930 11756 26936
rect 11532 26042 11560 26930
rect 11704 26784 11756 26790
rect 11704 26726 11756 26732
rect 11612 26308 11664 26314
rect 11612 26250 11664 26256
rect 11520 26036 11572 26042
rect 11520 25978 11572 25984
rect 11624 25974 11652 26250
rect 11612 25968 11664 25974
rect 11612 25910 11664 25916
rect 11428 24064 11480 24070
rect 11428 24006 11480 24012
rect 11336 23860 11388 23866
rect 11336 23802 11388 23808
rect 11348 22574 11376 23802
rect 11336 22568 11388 22574
rect 11336 22510 11388 22516
rect 11520 22094 11572 22098
rect 11716 22094 11744 26726
rect 11808 24664 11836 31726
rect 11888 29640 11940 29646
rect 11888 29582 11940 29588
rect 11900 28762 11928 29582
rect 11888 28756 11940 28762
rect 11888 28698 11940 28704
rect 12360 27470 12388 32166
rect 12452 29578 12480 32438
rect 13452 31748 13504 31754
rect 13452 31690 13504 31696
rect 12532 31340 12584 31346
rect 12532 31282 12584 31288
rect 12440 29572 12492 29578
rect 12440 29514 12492 29520
rect 12544 28626 12572 31282
rect 13464 31278 13492 31690
rect 13452 31272 13504 31278
rect 13452 31214 13504 31220
rect 12900 30592 12952 30598
rect 12900 30534 12952 30540
rect 12624 30320 12676 30326
rect 12624 30262 12676 30268
rect 12532 28620 12584 28626
rect 12532 28562 12584 28568
rect 12636 27470 12664 30262
rect 12912 28014 12940 30534
rect 13360 28960 13412 28966
rect 13360 28902 13412 28908
rect 12992 28552 13044 28558
rect 12992 28494 13044 28500
rect 12900 28008 12952 28014
rect 12900 27950 12952 27956
rect 12912 27470 12940 27950
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 12624 27464 12676 27470
rect 12624 27406 12676 27412
rect 12808 27464 12860 27470
rect 12808 27406 12860 27412
rect 12900 27464 12952 27470
rect 12900 27406 12952 27412
rect 11980 27328 12032 27334
rect 11980 27270 12032 27276
rect 11888 26036 11940 26042
rect 11888 25978 11940 25984
rect 11900 25498 11928 25978
rect 11888 25492 11940 25498
rect 11888 25434 11940 25440
rect 11888 24676 11940 24682
rect 11808 24636 11888 24664
rect 11888 24618 11940 24624
rect 11992 23662 12020 27270
rect 12820 27130 12848 27406
rect 12808 27124 12860 27130
rect 12808 27066 12860 27072
rect 12624 26308 12676 26314
rect 12624 26250 12676 26256
rect 12348 26240 12400 26246
rect 12348 26182 12400 26188
rect 12072 25900 12124 25906
rect 12072 25842 12124 25848
rect 12084 25362 12112 25842
rect 12164 25764 12216 25770
rect 12164 25706 12216 25712
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 12176 23798 12204 25706
rect 12360 25702 12388 26182
rect 12636 26042 12664 26250
rect 12624 26036 12676 26042
rect 12624 25978 12676 25984
rect 12624 25764 12676 25770
rect 12624 25706 12676 25712
rect 12348 25696 12400 25702
rect 12348 25638 12400 25644
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12544 25158 12572 25434
rect 12532 25152 12584 25158
rect 12532 25094 12584 25100
rect 12544 24954 12572 25094
rect 12636 24954 12664 25706
rect 12716 25220 12768 25226
rect 12716 25162 12768 25168
rect 12532 24948 12584 24954
rect 12532 24890 12584 24896
rect 12624 24948 12676 24954
rect 12624 24890 12676 24896
rect 12728 24750 12756 25162
rect 12716 24744 12768 24750
rect 12716 24686 12768 24692
rect 12532 24676 12584 24682
rect 12532 24618 12584 24624
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12164 23792 12216 23798
rect 12164 23734 12216 23740
rect 11980 23656 12032 23662
rect 11980 23598 12032 23604
rect 12268 23594 12296 23802
rect 12256 23588 12308 23594
rect 12256 23530 12308 23536
rect 11888 23520 11940 23526
rect 11888 23462 11940 23468
rect 12072 23520 12124 23526
rect 12072 23462 12124 23468
rect 11900 23322 11928 23462
rect 11888 23316 11940 23322
rect 11888 23258 11940 23264
rect 11900 22778 11928 23258
rect 11888 22772 11940 22778
rect 11888 22714 11940 22720
rect 11900 22438 11928 22714
rect 11888 22432 11940 22438
rect 11888 22374 11940 22380
rect 11900 22234 11928 22374
rect 11888 22228 11940 22234
rect 11888 22170 11940 22176
rect 11520 22092 11744 22094
rect 11572 22066 11744 22092
rect 11520 22034 11572 22040
rect 11980 21412 12032 21418
rect 11980 21354 12032 21360
rect 11992 21010 12020 21354
rect 11980 21004 12032 21010
rect 11980 20946 12032 20952
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 10968 20392 11020 20398
rect 10968 20334 11020 20340
rect 10600 20324 10652 20330
rect 10600 20266 10652 20272
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 10876 19712 10928 19718
rect 10876 19654 10928 19660
rect 10888 19514 10916 19654
rect 10876 19508 10928 19514
rect 10876 19450 10928 19456
rect 10324 19440 10376 19446
rect 10324 19382 10376 19388
rect 10336 18630 10364 19382
rect 10980 19378 11008 19722
rect 11256 19378 11284 20470
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 10968 19372 11020 19378
rect 10968 19314 11020 19320
rect 11244 19372 11296 19378
rect 11244 19314 11296 19320
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11072 18834 11100 19110
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10336 17678 10364 18566
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10232 17536 10284 17542
rect 10232 17478 10284 17484
rect 10244 17134 10272 17478
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10244 10062 10272 17070
rect 10336 16454 10364 17614
rect 11072 17338 11100 18158
rect 11256 17338 11284 19314
rect 11440 18970 11468 19790
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11428 18964 11480 18970
rect 11428 18906 11480 18912
rect 11060 17332 11112 17338
rect 11060 17274 11112 17280
rect 11244 17332 11296 17338
rect 11244 17274 11296 17280
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10232 10056 10284 10062
rect 10232 9998 10284 10004
rect 9312 8492 9364 8498
rect 9312 8434 9364 8440
rect 11808 2514 11836 19654
rect 11992 19514 12020 20946
rect 11980 19508 12032 19514
rect 11980 19450 12032 19456
rect 11992 17882 12020 19450
rect 12084 18698 12112 23462
rect 12452 22642 12480 24346
rect 12544 24070 12572 24618
rect 12728 24206 12756 24686
rect 12912 24410 12940 27406
rect 13004 24818 13032 28494
rect 13372 28422 13400 28902
rect 13360 28416 13412 28422
rect 13360 28358 13412 28364
rect 13084 28076 13136 28082
rect 13084 28018 13136 28024
rect 13096 25498 13124 28018
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 13188 25770 13216 27406
rect 13360 27328 13412 27334
rect 13360 27270 13412 27276
rect 13372 26790 13400 27270
rect 13360 26784 13412 26790
rect 13360 26726 13412 26732
rect 13372 26246 13400 26726
rect 13360 26240 13412 26246
rect 13360 26182 13412 26188
rect 13176 25764 13228 25770
rect 13176 25706 13228 25712
rect 13084 25492 13136 25498
rect 13084 25434 13136 25440
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 13096 24954 13124 25230
rect 13084 24948 13136 24954
rect 13084 24890 13136 24896
rect 12992 24812 13044 24818
rect 12992 24754 13044 24760
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 12716 24200 12768 24206
rect 12716 24142 12768 24148
rect 12900 24200 12952 24206
rect 12900 24142 12952 24148
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 12532 24064 12584 24070
rect 12532 24006 12584 24012
rect 12544 23526 12572 24006
rect 12636 23594 12664 24074
rect 12716 24064 12768 24070
rect 12716 24006 12768 24012
rect 12624 23588 12676 23594
rect 12624 23530 12676 23536
rect 12532 23520 12584 23526
rect 12532 23462 12584 23468
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12440 22432 12492 22438
rect 12440 22374 12492 22380
rect 12452 21962 12480 22374
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 12176 21146 12204 21286
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 12164 18080 12216 18086
rect 12164 18022 12216 18028
rect 11980 17876 12032 17882
rect 11980 17818 12032 17824
rect 12176 17610 12204 18022
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12544 6914 12572 23462
rect 12728 22642 12756 24006
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12820 22642 12848 23666
rect 12912 22982 12940 24142
rect 13004 24138 13032 24754
rect 13176 24608 13228 24614
rect 13176 24550 13228 24556
rect 12992 24132 13044 24138
rect 12992 24074 13044 24080
rect 13004 23730 13032 24074
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12900 22976 12952 22982
rect 12900 22918 12952 22924
rect 12716 22636 12768 22642
rect 12716 22578 12768 22584
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 12912 19334 12940 22918
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 13004 22094 13032 22578
rect 13004 22066 13124 22094
rect 13096 21894 13124 22066
rect 13084 21888 13136 21894
rect 13084 21830 13136 21836
rect 13188 20602 13216 24550
rect 13372 24206 13400 26182
rect 13464 25770 13492 31214
rect 13728 30660 13780 30666
rect 13728 30602 13780 30608
rect 13452 25764 13504 25770
rect 13452 25706 13504 25712
rect 13636 25492 13688 25498
rect 13636 25434 13688 25440
rect 13452 25152 13504 25158
rect 13452 25094 13504 25100
rect 13464 24886 13492 25094
rect 13452 24880 13504 24886
rect 13452 24822 13504 24828
rect 13648 24410 13676 25434
rect 13636 24404 13688 24410
rect 13636 24346 13688 24352
rect 13360 24200 13412 24206
rect 13360 24142 13412 24148
rect 13636 24064 13688 24070
rect 13636 24006 13688 24012
rect 13648 23866 13676 24006
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 13740 20942 13768 30602
rect 14936 25906 14964 59200
rect 19574 57692 19882 57701
rect 19574 57690 19580 57692
rect 19636 57690 19660 57692
rect 19716 57690 19740 57692
rect 19796 57690 19820 57692
rect 19876 57690 19882 57692
rect 19636 57638 19638 57690
rect 19818 57638 19820 57690
rect 19574 57636 19580 57638
rect 19636 57636 19660 57638
rect 19716 57636 19740 57638
rect 19796 57636 19820 57638
rect 19876 57636 19882 57638
rect 19574 57627 19882 57636
rect 44928 57526 44956 59200
rect 50294 57692 50602 57701
rect 50294 57690 50300 57692
rect 50356 57690 50380 57692
rect 50436 57690 50460 57692
rect 50516 57690 50540 57692
rect 50596 57690 50602 57692
rect 50356 57638 50358 57690
rect 50538 57638 50540 57690
rect 50294 57636 50300 57638
rect 50356 57636 50380 57638
rect 50436 57636 50460 57638
rect 50516 57636 50540 57638
rect 50596 57636 50602 57638
rect 50294 57627 50602 57636
rect 44916 57520 44968 57526
rect 44916 57462 44968 57468
rect 46480 57384 46532 57390
rect 46480 57326 46532 57332
rect 34934 57148 35242 57157
rect 34934 57146 34940 57148
rect 34996 57146 35020 57148
rect 35076 57146 35100 57148
rect 35156 57146 35180 57148
rect 35236 57146 35242 57148
rect 34996 57094 34998 57146
rect 35178 57094 35180 57146
rect 34934 57092 34940 57094
rect 34996 57092 35020 57094
rect 35076 57092 35100 57094
rect 35156 57092 35180 57094
rect 35236 57092 35242 57094
rect 34934 57083 35242 57092
rect 19574 56604 19882 56613
rect 19574 56602 19580 56604
rect 19636 56602 19660 56604
rect 19716 56602 19740 56604
rect 19796 56602 19820 56604
rect 19876 56602 19882 56604
rect 19636 56550 19638 56602
rect 19818 56550 19820 56602
rect 19574 56548 19580 56550
rect 19636 56548 19660 56550
rect 19716 56548 19740 56550
rect 19796 56548 19820 56550
rect 19876 56548 19882 56550
rect 19574 56539 19882 56548
rect 34934 56060 35242 56069
rect 34934 56058 34940 56060
rect 34996 56058 35020 56060
rect 35076 56058 35100 56060
rect 35156 56058 35180 56060
rect 35236 56058 35242 56060
rect 34996 56006 34998 56058
rect 35178 56006 35180 56058
rect 34934 56004 34940 56006
rect 34996 56004 35020 56006
rect 35076 56004 35100 56006
rect 35156 56004 35180 56006
rect 35236 56004 35242 56006
rect 34934 55995 35242 56004
rect 15844 55616 15896 55622
rect 15844 55558 15896 55564
rect 15856 31278 15884 55558
rect 19574 55516 19882 55525
rect 19574 55514 19580 55516
rect 19636 55514 19660 55516
rect 19716 55514 19740 55516
rect 19796 55514 19820 55516
rect 19876 55514 19882 55516
rect 19636 55462 19638 55514
rect 19818 55462 19820 55514
rect 19574 55460 19580 55462
rect 19636 55460 19660 55462
rect 19716 55460 19740 55462
rect 19796 55460 19820 55462
rect 19876 55460 19882 55462
rect 19574 55451 19882 55460
rect 34934 54972 35242 54981
rect 34934 54970 34940 54972
rect 34996 54970 35020 54972
rect 35076 54970 35100 54972
rect 35156 54970 35180 54972
rect 35236 54970 35242 54972
rect 34996 54918 34998 54970
rect 35178 54918 35180 54970
rect 34934 54916 34940 54918
rect 34996 54916 35020 54918
rect 35076 54916 35100 54918
rect 35156 54916 35180 54918
rect 35236 54916 35242 54918
rect 34934 54907 35242 54916
rect 19574 54428 19882 54437
rect 19574 54426 19580 54428
rect 19636 54426 19660 54428
rect 19716 54426 19740 54428
rect 19796 54426 19820 54428
rect 19876 54426 19882 54428
rect 19636 54374 19638 54426
rect 19818 54374 19820 54426
rect 19574 54372 19580 54374
rect 19636 54372 19660 54374
rect 19716 54372 19740 54374
rect 19796 54372 19820 54374
rect 19876 54372 19882 54374
rect 19574 54363 19882 54372
rect 34934 53884 35242 53893
rect 34934 53882 34940 53884
rect 34996 53882 35020 53884
rect 35076 53882 35100 53884
rect 35156 53882 35180 53884
rect 35236 53882 35242 53884
rect 34996 53830 34998 53882
rect 35178 53830 35180 53882
rect 34934 53828 34940 53830
rect 34996 53828 35020 53830
rect 35076 53828 35100 53830
rect 35156 53828 35180 53830
rect 35236 53828 35242 53830
rect 34934 53819 35242 53828
rect 19574 53340 19882 53349
rect 19574 53338 19580 53340
rect 19636 53338 19660 53340
rect 19716 53338 19740 53340
rect 19796 53338 19820 53340
rect 19876 53338 19882 53340
rect 19636 53286 19638 53338
rect 19818 53286 19820 53338
rect 19574 53284 19580 53286
rect 19636 53284 19660 53286
rect 19716 53284 19740 53286
rect 19796 53284 19820 53286
rect 19876 53284 19882 53286
rect 19574 53275 19882 53284
rect 34934 52796 35242 52805
rect 34934 52794 34940 52796
rect 34996 52794 35020 52796
rect 35076 52794 35100 52796
rect 35156 52794 35180 52796
rect 35236 52794 35242 52796
rect 34996 52742 34998 52794
rect 35178 52742 35180 52794
rect 34934 52740 34940 52742
rect 34996 52740 35020 52742
rect 35076 52740 35100 52742
rect 35156 52740 35180 52742
rect 35236 52740 35242 52742
rect 34934 52731 35242 52740
rect 19574 52252 19882 52261
rect 19574 52250 19580 52252
rect 19636 52250 19660 52252
rect 19716 52250 19740 52252
rect 19796 52250 19820 52252
rect 19876 52250 19882 52252
rect 19636 52198 19638 52250
rect 19818 52198 19820 52250
rect 19574 52196 19580 52198
rect 19636 52196 19660 52198
rect 19716 52196 19740 52198
rect 19796 52196 19820 52198
rect 19876 52196 19882 52198
rect 19574 52187 19882 52196
rect 34934 51708 35242 51717
rect 34934 51706 34940 51708
rect 34996 51706 35020 51708
rect 35076 51706 35100 51708
rect 35156 51706 35180 51708
rect 35236 51706 35242 51708
rect 34996 51654 34998 51706
rect 35178 51654 35180 51706
rect 34934 51652 34940 51654
rect 34996 51652 35020 51654
rect 35076 51652 35100 51654
rect 35156 51652 35180 51654
rect 35236 51652 35242 51654
rect 34934 51643 35242 51652
rect 19574 51164 19882 51173
rect 19574 51162 19580 51164
rect 19636 51162 19660 51164
rect 19716 51162 19740 51164
rect 19796 51162 19820 51164
rect 19876 51162 19882 51164
rect 19636 51110 19638 51162
rect 19818 51110 19820 51162
rect 19574 51108 19580 51110
rect 19636 51108 19660 51110
rect 19716 51108 19740 51110
rect 19796 51108 19820 51110
rect 19876 51108 19882 51110
rect 19574 51099 19882 51108
rect 34934 50620 35242 50629
rect 34934 50618 34940 50620
rect 34996 50618 35020 50620
rect 35076 50618 35100 50620
rect 35156 50618 35180 50620
rect 35236 50618 35242 50620
rect 34996 50566 34998 50618
rect 35178 50566 35180 50618
rect 34934 50564 34940 50566
rect 34996 50564 35020 50566
rect 35076 50564 35100 50566
rect 35156 50564 35180 50566
rect 35236 50564 35242 50566
rect 34934 50555 35242 50564
rect 19574 50076 19882 50085
rect 19574 50074 19580 50076
rect 19636 50074 19660 50076
rect 19716 50074 19740 50076
rect 19796 50074 19820 50076
rect 19876 50074 19882 50076
rect 19636 50022 19638 50074
rect 19818 50022 19820 50074
rect 19574 50020 19580 50022
rect 19636 50020 19660 50022
rect 19716 50020 19740 50022
rect 19796 50020 19820 50022
rect 19876 50020 19882 50022
rect 19574 50011 19882 50020
rect 34934 49532 35242 49541
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49467 35242 49476
rect 19574 48988 19882 48997
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48923 19882 48932
rect 34934 48444 35242 48453
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48379 35242 48388
rect 19574 47900 19882 47909
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47835 19882 47844
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 17132 35692 17184 35698
rect 17132 35634 17184 35640
rect 15844 31272 15896 31278
rect 15844 31214 15896 31220
rect 15384 30184 15436 30190
rect 15384 30126 15436 30132
rect 15016 29776 15068 29782
rect 15016 29718 15068 29724
rect 15028 29306 15056 29718
rect 15396 29510 15424 30126
rect 15856 29850 15884 31214
rect 17144 30666 17172 35634
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 41604 33992 41656 33998
rect 41604 33934 41656 33940
rect 45652 33992 45704 33998
rect 45652 33934 45704 33940
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 38384 33108 38436 33114
rect 38384 33050 38436 33056
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 38396 32570 38424 33050
rect 41616 32978 41644 33934
rect 41880 33924 41932 33930
rect 41880 33866 41932 33872
rect 44180 33924 44232 33930
rect 44180 33866 44232 33872
rect 41892 33658 41920 33866
rect 42616 33856 42668 33862
rect 42616 33798 42668 33804
rect 43260 33856 43312 33862
rect 43260 33798 43312 33804
rect 41880 33652 41932 33658
rect 41880 33594 41932 33600
rect 41604 32972 41656 32978
rect 41604 32914 41656 32920
rect 40592 32836 40644 32842
rect 40592 32778 40644 32784
rect 40604 32570 40632 32778
rect 41420 32768 41472 32774
rect 41420 32710 41472 32716
rect 38384 32564 38436 32570
rect 38384 32506 38436 32512
rect 40592 32564 40644 32570
rect 40592 32506 40644 32512
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 37740 31952 37792 31958
rect 37740 31894 37792 31900
rect 36268 31816 36320 31822
rect 36268 31758 36320 31764
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 17132 30660 17184 30666
rect 17132 30602 17184 30608
rect 36280 30598 36308 31758
rect 36728 31748 36780 31754
rect 36728 31690 36780 31696
rect 36740 31482 36768 31690
rect 36728 31476 36780 31482
rect 36728 31418 36780 31424
rect 37752 31346 37780 31894
rect 38396 31822 38424 32506
rect 39028 32428 39080 32434
rect 39028 32370 39080 32376
rect 39212 32428 39264 32434
rect 39212 32370 39264 32376
rect 39488 32428 39540 32434
rect 39488 32370 39540 32376
rect 38844 31884 38896 31890
rect 38844 31826 38896 31832
rect 38384 31816 38436 31822
rect 38384 31758 38436 31764
rect 37740 31340 37792 31346
rect 37740 31282 37792 31288
rect 38200 31340 38252 31346
rect 38200 31282 38252 31288
rect 38212 30938 38240 31282
rect 38200 30932 38252 30938
rect 38200 30874 38252 30880
rect 38292 30660 38344 30666
rect 38292 30602 38344 30608
rect 36268 30592 36320 30598
rect 36268 30534 36320 30540
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 31024 30116 31076 30122
rect 31024 30058 31076 30064
rect 31036 29850 31064 30058
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 15844 29844 15896 29850
rect 15844 29786 15896 29792
rect 31024 29844 31076 29850
rect 31024 29786 31076 29792
rect 15856 29714 15884 29786
rect 36280 29714 36308 30534
rect 38304 30122 38332 30602
rect 37372 30116 37424 30122
rect 37372 30058 37424 30064
rect 38292 30116 38344 30122
rect 38292 30058 38344 30064
rect 15844 29708 15896 29714
rect 15844 29650 15896 29656
rect 36268 29708 36320 29714
rect 36268 29650 36320 29656
rect 37188 29708 37240 29714
rect 37188 29650 37240 29656
rect 15384 29504 15436 29510
rect 15384 29446 15436 29452
rect 15016 29300 15068 29306
rect 15016 29242 15068 29248
rect 14924 25900 14976 25906
rect 14924 25842 14976 25848
rect 13820 24336 13872 24342
rect 13820 24278 13872 24284
rect 13832 23866 13860 24278
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 12452 6886 12572 6914
rect 12820 19306 12940 19334
rect 11796 2508 11848 2514
rect 11796 2450 11848 2456
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 7564 2372 7616 2378
rect 7564 2314 7616 2320
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 2608 800 2636 2314
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4080 2038 4108 2246
rect 4068 2032 4120 2038
rect 4068 1974 4120 1980
rect 7576 800 7604 2314
rect 12452 2310 12480 6886
rect 12820 2650 12848 19306
rect 15396 2650 15424 29446
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 36280 28762 36308 29650
rect 37200 29306 37228 29650
rect 37188 29300 37240 29306
rect 37188 29242 37240 29248
rect 37384 29170 37412 30058
rect 37648 29572 37700 29578
rect 37648 29514 37700 29520
rect 37464 29504 37516 29510
rect 37464 29446 37516 29452
rect 37372 29164 37424 29170
rect 37372 29106 37424 29112
rect 37476 29034 37504 29446
rect 37660 29238 37688 29514
rect 37648 29232 37700 29238
rect 37648 29174 37700 29180
rect 37832 29096 37884 29102
rect 37832 29038 37884 29044
rect 37464 29028 37516 29034
rect 37464 28970 37516 28976
rect 36268 28756 36320 28762
rect 36268 28698 36320 28704
rect 37464 28756 37516 28762
rect 37464 28698 37516 28704
rect 37476 28490 37504 28698
rect 37464 28484 37516 28490
rect 37464 28426 37516 28432
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 25320 27396 25372 27402
rect 25320 27338 25372 27344
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 25332 27062 25360 27338
rect 25320 27056 25372 27062
rect 25320 26998 25372 27004
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 25332 25498 25360 26998
rect 37280 26920 37332 26926
rect 37280 26862 37332 26868
rect 36268 26784 36320 26790
rect 36268 26726 36320 26732
rect 36728 26784 36780 26790
rect 36728 26726 36780 26732
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35440 26444 35492 26450
rect 35440 26386 35492 26392
rect 31116 25764 31168 25770
rect 31116 25706 31168 25712
rect 25320 25492 25372 25498
rect 25320 25434 25372 25440
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19984 21412 20036 21418
rect 19984 21354 20036 21360
rect 18236 20936 18288 20942
rect 18236 20878 18288 20884
rect 18248 20466 18276 20878
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19996 20602 20024 21354
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 18236 20460 18288 20466
rect 18236 20402 18288 20408
rect 31128 20262 31156 25706
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35452 24274 35480 26386
rect 35716 26308 35768 26314
rect 35716 26250 35768 26256
rect 35728 26042 35756 26250
rect 36280 26042 36308 26726
rect 36740 26314 36768 26726
rect 36728 26308 36780 26314
rect 36728 26250 36780 26256
rect 35716 26036 35768 26042
rect 35716 25978 35768 25984
rect 36268 26036 36320 26042
rect 36268 25978 36320 25984
rect 36544 25832 36596 25838
rect 36544 25774 36596 25780
rect 36556 25498 36584 25774
rect 36544 25492 36596 25498
rect 36544 25434 36596 25440
rect 36740 24614 36768 26250
rect 37096 26240 37148 26246
rect 37096 26182 37148 26188
rect 37108 26042 37136 26182
rect 37292 26042 37320 26862
rect 37476 26790 37504 28426
rect 37464 26784 37516 26790
rect 37464 26726 37516 26732
rect 37844 26382 37872 29038
rect 38016 28960 38068 28966
rect 38016 28902 38068 28908
rect 38028 28694 38056 28902
rect 38396 28762 38424 31758
rect 38476 31680 38528 31686
rect 38476 31622 38528 31628
rect 38660 31680 38712 31686
rect 38660 31622 38712 31628
rect 38488 31346 38516 31622
rect 38672 31482 38700 31622
rect 38856 31482 38884 31826
rect 38660 31476 38712 31482
rect 38660 31418 38712 31424
rect 38844 31476 38896 31482
rect 38844 31418 38896 31424
rect 38476 31340 38528 31346
rect 38476 31282 38528 31288
rect 38660 31340 38712 31346
rect 38660 31282 38712 31288
rect 38672 30938 38700 31282
rect 38660 30932 38712 30938
rect 38660 30874 38712 30880
rect 38856 30734 38884 31418
rect 39040 31346 39068 32370
rect 39224 31872 39252 32370
rect 39304 32224 39356 32230
rect 39304 32166 39356 32172
rect 39396 32224 39448 32230
rect 39396 32166 39448 32172
rect 39132 31844 39252 31872
rect 39028 31340 39080 31346
rect 39028 31282 39080 31288
rect 39132 31210 39160 31844
rect 39316 31754 39344 32166
rect 39408 32026 39436 32166
rect 39396 32020 39448 32026
rect 39396 31962 39448 31968
rect 39224 31726 39344 31754
rect 39396 31748 39448 31754
rect 39120 31204 39172 31210
rect 39120 31146 39172 31152
rect 38844 30728 38896 30734
rect 38844 30670 38896 30676
rect 39224 30258 39252 31726
rect 39396 31690 39448 31696
rect 39408 31346 39436 31690
rect 39500 31482 39528 32370
rect 40592 32360 40644 32366
rect 40592 32302 40644 32308
rect 40604 32026 40632 32302
rect 41236 32224 41288 32230
rect 41236 32166 41288 32172
rect 40592 32020 40644 32026
rect 40592 31962 40644 31968
rect 41248 31890 41276 32166
rect 40040 31884 40092 31890
rect 40040 31826 40092 31832
rect 41236 31884 41288 31890
rect 41236 31826 41288 31832
rect 39948 31816 40000 31822
rect 39948 31758 40000 31764
rect 39488 31476 39540 31482
rect 39488 31418 39540 31424
rect 39396 31340 39448 31346
rect 39396 31282 39448 31288
rect 39408 31210 39436 31282
rect 39396 31204 39448 31210
rect 39396 31146 39448 31152
rect 39960 30938 39988 31758
rect 40052 31754 40080 31826
rect 41432 31754 41460 32710
rect 41616 31890 41644 32914
rect 42628 32910 42656 33798
rect 43272 33590 43300 33798
rect 43260 33584 43312 33590
rect 43260 33526 43312 33532
rect 42892 33516 42944 33522
rect 42892 33458 42944 33464
rect 42904 32910 42932 33458
rect 43260 33448 43312 33454
rect 43260 33390 43312 33396
rect 43272 33046 43300 33390
rect 43812 33380 43864 33386
rect 43812 33322 43864 33328
rect 43260 33040 43312 33046
rect 43260 32982 43312 32988
rect 43272 32910 43300 32982
rect 42616 32904 42668 32910
rect 42616 32846 42668 32852
rect 42708 32904 42760 32910
rect 42708 32846 42760 32852
rect 42892 32904 42944 32910
rect 42892 32846 42944 32852
rect 43260 32904 43312 32910
rect 43260 32846 43312 32852
rect 43536 32904 43588 32910
rect 43536 32846 43588 32852
rect 43720 32904 43772 32910
rect 43720 32846 43772 32852
rect 42156 32768 42208 32774
rect 42156 32710 42208 32716
rect 42168 32570 42196 32710
rect 42720 32570 42748 32846
rect 42800 32836 42852 32842
rect 42800 32778 42852 32784
rect 42812 32570 42840 32778
rect 42904 32570 42932 32846
rect 43548 32774 43576 32846
rect 43076 32768 43128 32774
rect 43076 32710 43128 32716
rect 43536 32768 43588 32774
rect 43536 32710 43588 32716
rect 42156 32564 42208 32570
rect 42156 32506 42208 32512
rect 42708 32564 42760 32570
rect 42708 32506 42760 32512
rect 42800 32564 42852 32570
rect 42800 32506 42852 32512
rect 42892 32564 42944 32570
rect 42892 32506 42944 32512
rect 43088 32434 43116 32710
rect 43732 32502 43760 32846
rect 43824 32842 43852 33322
rect 44086 33144 44142 33153
rect 44086 33079 44088 33088
rect 44140 33079 44142 33088
rect 44088 33050 44140 33056
rect 43812 32836 43864 32842
rect 43812 32778 43864 32784
rect 43824 32502 43852 32778
rect 43720 32496 43772 32502
rect 43720 32438 43772 32444
rect 43812 32496 43864 32502
rect 43812 32438 43864 32444
rect 44192 32450 44220 33866
rect 45468 33856 45520 33862
rect 45468 33798 45520 33804
rect 44640 33584 44692 33590
rect 44640 33526 44692 33532
rect 44272 33108 44324 33114
rect 44272 33050 44324 33056
rect 44284 32570 44312 33050
rect 44652 32994 44680 33526
rect 44824 33312 44876 33318
rect 44824 33254 44876 33260
rect 44560 32966 44680 32994
rect 44456 32836 44508 32842
rect 44456 32778 44508 32784
rect 44272 32564 44324 32570
rect 44272 32506 44324 32512
rect 42892 32428 42944 32434
rect 42892 32370 42944 32376
rect 43076 32428 43128 32434
rect 44192 32422 44404 32450
rect 43076 32370 43128 32376
rect 42064 32360 42116 32366
rect 42064 32302 42116 32308
rect 42076 32026 42104 32302
rect 42064 32020 42116 32026
rect 42064 31962 42116 31968
rect 41604 31884 41656 31890
rect 41604 31826 41656 31832
rect 40052 31726 40264 31754
rect 40236 31346 40264 31726
rect 41420 31748 41472 31754
rect 41420 31690 41472 31696
rect 40224 31340 40276 31346
rect 40224 31282 40276 31288
rect 40132 31136 40184 31142
rect 40132 31078 40184 31084
rect 39948 30932 40000 30938
rect 39948 30874 40000 30880
rect 39580 30796 39632 30802
rect 39580 30738 39632 30744
rect 39212 30252 39264 30258
rect 39212 30194 39264 30200
rect 39396 30252 39448 30258
rect 39396 30194 39448 30200
rect 39488 30252 39540 30258
rect 39488 30194 39540 30200
rect 38660 30048 38712 30054
rect 38660 29990 38712 29996
rect 38936 30048 38988 30054
rect 38936 29990 38988 29996
rect 38672 29782 38700 29990
rect 38660 29776 38712 29782
rect 38660 29718 38712 29724
rect 38948 29510 38976 29990
rect 39408 29714 39436 30194
rect 39396 29708 39448 29714
rect 39396 29650 39448 29656
rect 38936 29504 38988 29510
rect 38936 29446 38988 29452
rect 39212 29164 39264 29170
rect 39212 29106 39264 29112
rect 39028 29096 39080 29102
rect 39028 29038 39080 29044
rect 38660 29028 38712 29034
rect 38660 28970 38712 28976
rect 38384 28756 38436 28762
rect 38384 28698 38436 28704
rect 38016 28688 38068 28694
rect 38016 28630 38068 28636
rect 38568 28552 38620 28558
rect 38568 28494 38620 28500
rect 38476 28416 38528 28422
rect 38476 28358 38528 28364
rect 38488 28218 38516 28358
rect 38580 28218 38608 28494
rect 38672 28490 38700 28970
rect 39040 28762 39068 29038
rect 39028 28756 39080 28762
rect 39028 28698 39080 28704
rect 38660 28484 38712 28490
rect 38660 28426 38712 28432
rect 38476 28212 38528 28218
rect 38476 28154 38528 28160
rect 38568 28212 38620 28218
rect 38568 28154 38620 28160
rect 38108 28076 38160 28082
rect 38108 28018 38160 28024
rect 37924 27872 37976 27878
rect 37924 27814 37976 27820
rect 37936 27470 37964 27814
rect 37924 27464 37976 27470
rect 37924 27406 37976 27412
rect 38016 27464 38068 27470
rect 38016 27406 38068 27412
rect 38028 27130 38056 27406
rect 38016 27124 38068 27130
rect 38016 27066 38068 27072
rect 38120 27062 38148 28018
rect 38672 27470 38700 28426
rect 39224 28218 39252 29106
rect 39408 29016 39436 29650
rect 39500 29510 39528 30194
rect 39592 29714 39620 30738
rect 40144 30734 40172 31078
rect 41328 30796 41380 30802
rect 41328 30738 41380 30744
rect 40040 30728 40092 30734
rect 40040 30670 40092 30676
rect 40132 30728 40184 30734
rect 40132 30670 40184 30676
rect 40052 30394 40080 30670
rect 40040 30388 40092 30394
rect 40040 30330 40092 30336
rect 39764 30048 39816 30054
rect 39764 29990 39816 29996
rect 39580 29708 39632 29714
rect 39580 29650 39632 29656
rect 39592 29510 39620 29650
rect 39776 29646 39804 29990
rect 39948 29844 40000 29850
rect 39948 29786 40000 29792
rect 39764 29640 39816 29646
rect 39764 29582 39816 29588
rect 39960 29594 39988 29786
rect 40052 29714 40080 30330
rect 40408 30252 40460 30258
rect 40408 30194 40460 30200
rect 40040 29708 40092 29714
rect 40040 29650 40092 29656
rect 39960 29566 40172 29594
rect 39488 29504 39540 29510
rect 39488 29446 39540 29452
rect 39580 29504 39632 29510
rect 39580 29446 39632 29452
rect 40040 29504 40092 29510
rect 40040 29446 40092 29452
rect 39488 29028 39540 29034
rect 39408 28988 39488 29016
rect 39488 28970 39540 28976
rect 39304 28416 39356 28422
rect 39304 28358 39356 28364
rect 39212 28212 39264 28218
rect 39212 28154 39264 28160
rect 39224 27538 39252 28154
rect 39212 27532 39264 27538
rect 39212 27474 39264 27480
rect 38476 27464 38528 27470
rect 38660 27464 38712 27470
rect 38528 27424 38608 27452
rect 38476 27406 38528 27412
rect 38580 27130 38608 27424
rect 38660 27406 38712 27412
rect 38672 27334 38700 27406
rect 39316 27334 39344 28358
rect 40052 28218 40080 29446
rect 40144 29306 40172 29566
rect 40132 29300 40184 29306
rect 40132 29242 40184 29248
rect 40040 28212 40092 28218
rect 40040 28154 40092 28160
rect 40420 28082 40448 30194
rect 41340 29850 41368 30738
rect 41432 30326 41460 31690
rect 41616 31278 41644 31826
rect 42904 31686 42932 32370
rect 43088 32026 43116 32370
rect 43628 32360 43680 32366
rect 43628 32302 43680 32308
rect 44180 32360 44232 32366
rect 44180 32302 44232 32308
rect 43076 32020 43128 32026
rect 43076 31962 43128 31968
rect 43352 31952 43404 31958
rect 43352 31894 43404 31900
rect 42892 31680 42944 31686
rect 42892 31622 42944 31628
rect 41604 31272 41656 31278
rect 41604 31214 41656 31220
rect 42524 31272 42576 31278
rect 42524 31214 42576 31220
rect 41972 30796 42024 30802
rect 41972 30738 42024 30744
rect 41420 30320 41472 30326
rect 41420 30262 41472 30268
rect 41328 29844 41380 29850
rect 41328 29786 41380 29792
rect 41432 29578 41460 30262
rect 41984 30190 42012 30738
rect 42536 30190 42564 31214
rect 43168 31204 43220 31210
rect 43168 31146 43220 31152
rect 43180 30734 43208 31146
rect 42984 30728 43036 30734
rect 42984 30670 43036 30676
rect 43168 30728 43220 30734
rect 43168 30670 43220 30676
rect 42800 30660 42852 30666
rect 42800 30602 42852 30608
rect 42812 30258 42840 30602
rect 42800 30252 42852 30258
rect 42800 30194 42852 30200
rect 41972 30184 42024 30190
rect 41972 30126 42024 30132
rect 42524 30184 42576 30190
rect 42524 30126 42576 30132
rect 41984 29646 42012 30126
rect 42536 29646 42564 30126
rect 41972 29640 42024 29646
rect 41972 29582 42024 29588
rect 42524 29640 42576 29646
rect 42524 29582 42576 29588
rect 40960 29572 41012 29578
rect 40960 29514 41012 29520
rect 41420 29572 41472 29578
rect 41420 29514 41472 29520
rect 40972 29238 41000 29514
rect 40960 29232 41012 29238
rect 40960 29174 41012 29180
rect 40684 28960 40736 28966
rect 40684 28902 40736 28908
rect 40696 28762 40724 28902
rect 40684 28756 40736 28762
rect 40684 28698 40736 28704
rect 41326 28112 41382 28121
rect 40040 28076 40092 28082
rect 40040 28018 40092 28024
rect 40224 28076 40276 28082
rect 40224 28018 40276 28024
rect 40408 28076 40460 28082
rect 40408 28018 40460 28024
rect 40684 28076 40736 28082
rect 41984 28082 42012 29582
rect 42248 28960 42300 28966
rect 42248 28902 42300 28908
rect 42260 28626 42288 28902
rect 42248 28620 42300 28626
rect 42248 28562 42300 28568
rect 42536 28558 42564 29582
rect 42800 29096 42852 29102
rect 42800 29038 42852 29044
rect 42812 28762 42840 29038
rect 42800 28756 42852 28762
rect 42800 28698 42852 28704
rect 42800 28620 42852 28626
rect 42800 28562 42852 28568
rect 42524 28552 42576 28558
rect 42524 28494 42576 28500
rect 41326 28047 41328 28056
rect 40684 28018 40736 28024
rect 41380 28047 41382 28056
rect 41972 28076 42024 28082
rect 41328 28018 41380 28024
rect 41972 28018 42024 28024
rect 39672 28008 39724 28014
rect 39672 27950 39724 27956
rect 39684 27674 39712 27950
rect 40052 27674 40080 28018
rect 40236 27962 40264 28018
rect 40144 27934 40264 27962
rect 40316 28008 40368 28014
rect 40316 27950 40368 27956
rect 40420 27962 40448 28018
rect 39672 27668 39724 27674
rect 39672 27610 39724 27616
rect 40040 27668 40092 27674
rect 40040 27610 40092 27616
rect 39396 27464 39448 27470
rect 39396 27406 39448 27412
rect 39856 27464 39908 27470
rect 39856 27406 39908 27412
rect 38660 27328 38712 27334
rect 38660 27270 38712 27276
rect 39212 27328 39264 27334
rect 39212 27270 39264 27276
rect 39304 27328 39356 27334
rect 39304 27270 39356 27276
rect 38568 27124 38620 27130
rect 38568 27066 38620 27072
rect 38108 27056 38160 27062
rect 38108 26998 38160 27004
rect 38120 26382 38148 26998
rect 38672 26858 38700 27270
rect 38752 26988 38804 26994
rect 38752 26930 38804 26936
rect 38844 26988 38896 26994
rect 38844 26930 38896 26936
rect 38660 26852 38712 26858
rect 38660 26794 38712 26800
rect 37832 26376 37884 26382
rect 37832 26318 37884 26324
rect 38108 26376 38160 26382
rect 38108 26318 38160 26324
rect 37844 26042 37872 26318
rect 38764 26314 38792 26930
rect 38752 26308 38804 26314
rect 38752 26250 38804 26256
rect 38856 26246 38884 26930
rect 39120 26784 39172 26790
rect 39120 26726 39172 26732
rect 39132 26518 39160 26726
rect 39224 26518 39252 27270
rect 39408 27062 39436 27406
rect 39396 27056 39448 27062
rect 39396 26998 39448 27004
rect 39120 26512 39172 26518
rect 39120 26454 39172 26460
rect 39212 26512 39264 26518
rect 39212 26454 39264 26460
rect 39224 26382 39252 26454
rect 39212 26376 39264 26382
rect 39212 26318 39264 26324
rect 39120 26308 39172 26314
rect 39120 26250 39172 26256
rect 37924 26240 37976 26246
rect 37924 26182 37976 26188
rect 38844 26240 38896 26246
rect 38844 26182 38896 26188
rect 37936 26042 37964 26182
rect 37096 26036 37148 26042
rect 37096 25978 37148 25984
rect 37280 26036 37332 26042
rect 37280 25978 37332 25984
rect 37832 26036 37884 26042
rect 37832 25978 37884 25984
rect 37924 26036 37976 26042
rect 37924 25978 37976 25984
rect 37108 25906 37136 25978
rect 38856 25974 38884 26182
rect 39132 26042 39160 26250
rect 39120 26036 39172 26042
rect 39120 25978 39172 25984
rect 37372 25968 37424 25974
rect 37372 25910 37424 25916
rect 37648 25968 37700 25974
rect 37648 25910 37700 25916
rect 38844 25968 38896 25974
rect 38844 25910 38896 25916
rect 36912 25900 36964 25906
rect 36912 25842 36964 25848
rect 37096 25900 37148 25906
rect 37096 25842 37148 25848
rect 36924 25498 36952 25842
rect 36912 25492 36964 25498
rect 36912 25434 36964 25440
rect 36820 25288 36872 25294
rect 36820 25230 36872 25236
rect 36832 24818 36860 25230
rect 36820 24812 36872 24818
rect 36820 24754 36872 24760
rect 35900 24608 35952 24614
rect 35900 24550 35952 24556
rect 36728 24608 36780 24614
rect 36728 24550 36780 24556
rect 34520 24268 34572 24274
rect 34520 24210 34572 24216
rect 35440 24268 35492 24274
rect 35440 24210 35492 24216
rect 34532 21418 34560 24210
rect 35912 24138 35940 24550
rect 35440 24132 35492 24138
rect 35440 24074 35492 24080
rect 35900 24132 35952 24138
rect 35900 24074 35952 24080
rect 35452 23866 35480 24074
rect 35440 23860 35492 23866
rect 35440 23802 35492 23808
rect 36832 23730 36860 24754
rect 37004 24064 37056 24070
rect 37004 24006 37056 24012
rect 37016 23866 37044 24006
rect 37004 23860 37056 23866
rect 37004 23802 37056 23808
rect 37108 23730 37136 25842
rect 37384 24818 37412 25910
rect 37464 25492 37516 25498
rect 37464 25434 37516 25440
rect 37476 25294 37504 25434
rect 37660 25430 37688 25910
rect 37740 25900 37792 25906
rect 37740 25842 37792 25848
rect 39212 25900 39264 25906
rect 39212 25842 39264 25848
rect 37752 25702 37780 25842
rect 37740 25696 37792 25702
rect 37740 25638 37792 25644
rect 38568 25492 38620 25498
rect 38568 25434 38620 25440
rect 37648 25424 37700 25430
rect 37648 25366 37700 25372
rect 37660 25294 37688 25366
rect 37464 25288 37516 25294
rect 37464 25230 37516 25236
rect 37648 25288 37700 25294
rect 37648 25230 37700 25236
rect 37832 25288 37884 25294
rect 37832 25230 37884 25236
rect 37372 24812 37424 24818
rect 37372 24754 37424 24760
rect 37188 24744 37240 24750
rect 37188 24686 37240 24692
rect 37200 24410 37228 24686
rect 37384 24682 37412 24754
rect 37372 24676 37424 24682
rect 37372 24618 37424 24624
rect 37280 24608 37332 24614
rect 37280 24550 37332 24556
rect 37188 24404 37240 24410
rect 37188 24346 37240 24352
rect 37292 23866 37320 24550
rect 37844 24274 37872 25230
rect 38476 24812 38528 24818
rect 38476 24754 38528 24760
rect 38016 24608 38068 24614
rect 38016 24550 38068 24556
rect 37832 24268 37884 24274
rect 37832 24210 37884 24216
rect 37556 24200 37608 24206
rect 37556 24142 37608 24148
rect 37280 23860 37332 23866
rect 37280 23802 37332 23808
rect 36820 23724 36872 23730
rect 36820 23666 36872 23672
rect 37096 23724 37148 23730
rect 37096 23666 37148 23672
rect 37568 23526 37596 24142
rect 38028 23866 38056 24550
rect 38384 24064 38436 24070
rect 38384 24006 38436 24012
rect 38396 23866 38424 24006
rect 38488 23866 38516 24754
rect 38580 24206 38608 25434
rect 38936 25288 38988 25294
rect 38936 25230 38988 25236
rect 38948 24954 38976 25230
rect 39224 25158 39252 25842
rect 39408 25702 39436 26998
rect 39868 26994 39896 27406
rect 40144 26994 40172 27934
rect 40224 27872 40276 27878
rect 40224 27814 40276 27820
rect 40236 27470 40264 27814
rect 40328 27674 40356 27950
rect 40420 27934 40540 27962
rect 40408 27872 40460 27878
rect 40408 27814 40460 27820
rect 40316 27668 40368 27674
rect 40316 27610 40368 27616
rect 40224 27464 40276 27470
rect 40224 27406 40276 27412
rect 39856 26988 39908 26994
rect 39856 26930 39908 26936
rect 39948 26988 40000 26994
rect 39948 26930 40000 26936
rect 40132 26988 40184 26994
rect 40132 26930 40184 26936
rect 39960 26518 39988 26930
rect 40224 26920 40276 26926
rect 40224 26862 40276 26868
rect 40236 26586 40264 26862
rect 40224 26580 40276 26586
rect 40224 26522 40276 26528
rect 39948 26512 40000 26518
rect 39948 26454 40000 26460
rect 39396 25696 39448 25702
rect 39396 25638 39448 25644
rect 40040 25288 40092 25294
rect 40040 25230 40092 25236
rect 39212 25152 39264 25158
rect 39212 25094 39264 25100
rect 40052 24954 40080 25230
rect 38936 24948 38988 24954
rect 38936 24890 38988 24896
rect 40040 24948 40092 24954
rect 40040 24890 40092 24896
rect 39028 24812 39080 24818
rect 39028 24754 39080 24760
rect 39764 24812 39816 24818
rect 39764 24754 39816 24760
rect 39040 24410 39068 24754
rect 39028 24404 39080 24410
rect 39028 24346 39080 24352
rect 39776 24206 39804 24754
rect 40052 24410 40080 24890
rect 40040 24404 40092 24410
rect 40040 24346 40092 24352
rect 38568 24200 38620 24206
rect 38568 24142 38620 24148
rect 39120 24200 39172 24206
rect 39120 24142 39172 24148
rect 39396 24200 39448 24206
rect 39396 24142 39448 24148
rect 39764 24200 39816 24206
rect 39764 24142 39816 24148
rect 38580 23866 38608 24142
rect 39132 23866 39160 24142
rect 38016 23860 38068 23866
rect 38016 23802 38068 23808
rect 38384 23860 38436 23866
rect 38384 23802 38436 23808
rect 38476 23860 38528 23866
rect 38476 23802 38528 23808
rect 38568 23860 38620 23866
rect 38568 23802 38620 23808
rect 39120 23860 39172 23866
rect 39120 23802 39172 23808
rect 39408 23798 39436 24142
rect 39396 23792 39448 23798
rect 39396 23734 39448 23740
rect 39396 23656 39448 23662
rect 39396 23598 39448 23604
rect 37556 23520 37608 23526
rect 37556 23462 37608 23468
rect 37740 23520 37792 23526
rect 37740 23462 37792 23468
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 37752 23050 37780 23462
rect 39408 23322 39436 23598
rect 40236 23322 40264 26522
rect 40420 26466 40448 27814
rect 40512 27538 40540 27934
rect 40500 27532 40552 27538
rect 40500 27474 40552 27480
rect 40696 27470 40724 28018
rect 40684 27464 40736 27470
rect 40684 27406 40736 27412
rect 40696 26790 40724 27406
rect 42156 27328 42208 27334
rect 42156 27270 42208 27276
rect 42168 27062 42196 27270
rect 42156 27056 42208 27062
rect 42156 26998 42208 27004
rect 40684 26784 40736 26790
rect 40684 26726 40736 26732
rect 40592 26580 40644 26586
rect 40592 26522 40644 26528
rect 40328 26450 40448 26466
rect 40316 26444 40448 26450
rect 40368 26438 40448 26444
rect 40316 26386 40368 26392
rect 40408 26376 40460 26382
rect 40408 26318 40460 26324
rect 40420 25974 40448 26318
rect 40408 25968 40460 25974
rect 40408 25910 40460 25916
rect 40420 25498 40448 25910
rect 40408 25492 40460 25498
rect 40408 25434 40460 25440
rect 40604 25362 40632 26522
rect 40592 25356 40644 25362
rect 40592 25298 40644 25304
rect 40696 24818 40724 26726
rect 41696 26512 41748 26518
rect 41696 26454 41748 26460
rect 40776 26240 40828 26246
rect 40776 26182 40828 26188
rect 40788 25430 40816 26182
rect 41420 25696 41472 25702
rect 41420 25638 41472 25644
rect 41604 25696 41656 25702
rect 41604 25638 41656 25644
rect 41432 25498 41460 25638
rect 41420 25492 41472 25498
rect 41420 25434 41472 25440
rect 40776 25424 40828 25430
rect 40776 25366 40828 25372
rect 41512 25424 41564 25430
rect 41512 25366 41564 25372
rect 41052 25220 41104 25226
rect 41052 25162 41104 25168
rect 40960 25152 41012 25158
rect 40960 25094 41012 25100
rect 40972 24818 41000 25094
rect 41064 24954 41092 25162
rect 41052 24948 41104 24954
rect 41052 24890 41104 24896
rect 41524 24818 41552 25366
rect 41616 25294 41644 25638
rect 41708 25294 41736 26454
rect 42168 26246 42196 26998
rect 42432 26988 42484 26994
rect 42432 26930 42484 26936
rect 42340 26784 42392 26790
rect 42340 26726 42392 26732
rect 42352 26450 42380 26726
rect 42444 26586 42472 26930
rect 42432 26580 42484 26586
rect 42432 26522 42484 26528
rect 42340 26444 42392 26450
rect 42340 26386 42392 26392
rect 42156 26240 42208 26246
rect 42156 26182 42208 26188
rect 41604 25288 41656 25294
rect 41604 25230 41656 25236
rect 41696 25288 41748 25294
rect 41696 25230 41748 25236
rect 41880 25288 41932 25294
rect 41880 25230 41932 25236
rect 41616 24818 41644 25230
rect 41788 25220 41840 25226
rect 41788 25162 41840 25168
rect 40684 24812 40736 24818
rect 40684 24754 40736 24760
rect 40960 24812 41012 24818
rect 40960 24754 41012 24760
rect 41512 24812 41564 24818
rect 41512 24754 41564 24760
rect 41604 24812 41656 24818
rect 41604 24754 41656 24760
rect 41328 24200 41380 24206
rect 41328 24142 41380 24148
rect 40868 23520 40920 23526
rect 40868 23462 40920 23468
rect 39396 23316 39448 23322
rect 39396 23258 39448 23264
rect 40224 23316 40276 23322
rect 40224 23258 40276 23264
rect 39396 23112 39448 23118
rect 39396 23054 39448 23060
rect 37740 23044 37792 23050
rect 37740 22986 37792 22992
rect 39408 22778 39436 23054
rect 39764 23044 39816 23050
rect 39764 22986 39816 22992
rect 40132 23044 40184 23050
rect 40132 22986 40184 22992
rect 39396 22772 39448 22778
rect 39396 22714 39448 22720
rect 39776 22574 39804 22986
rect 40144 22778 40172 22986
rect 40880 22778 40908 23462
rect 41236 23112 41288 23118
rect 41236 23054 41288 23060
rect 40132 22772 40184 22778
rect 40132 22714 40184 22720
rect 40868 22772 40920 22778
rect 40868 22714 40920 22720
rect 41248 22574 41276 23054
rect 39764 22568 39816 22574
rect 39764 22510 39816 22516
rect 41236 22568 41288 22574
rect 41236 22510 41288 22516
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 41340 22098 41368 24142
rect 41604 24132 41656 24138
rect 41604 24074 41656 24080
rect 41616 23866 41644 24074
rect 41604 23860 41656 23866
rect 41604 23802 41656 23808
rect 41328 22092 41380 22098
rect 41328 22034 41380 22040
rect 34520 21412 34572 21418
rect 34520 21354 34572 21360
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 31116 20256 31168 20262
rect 31116 20198 31168 20204
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 41800 19854 41828 25162
rect 41892 24954 41920 25230
rect 41880 24948 41932 24954
rect 41880 24890 41932 24896
rect 42168 24274 42196 26182
rect 42248 25492 42300 25498
rect 42248 25434 42300 25440
rect 42260 24614 42288 25434
rect 42536 25362 42564 28494
rect 42616 26988 42668 26994
rect 42616 26930 42668 26936
rect 42628 25498 42656 26930
rect 42812 26586 42840 28562
rect 42996 27674 43024 30670
rect 43076 30592 43128 30598
rect 43076 30534 43128 30540
rect 43088 30394 43116 30534
rect 43076 30388 43128 30394
rect 43076 30330 43128 30336
rect 43076 28416 43128 28422
rect 43076 28358 43128 28364
rect 42984 27668 43036 27674
rect 42984 27610 43036 27616
rect 42892 27328 42944 27334
rect 42892 27270 42944 27276
rect 42904 27130 42932 27270
rect 43088 27130 43116 28358
rect 42892 27124 42944 27130
rect 42892 27066 42944 27072
rect 42984 27124 43036 27130
rect 42984 27066 43036 27072
rect 43076 27124 43128 27130
rect 43076 27066 43128 27072
rect 42996 27010 43024 27066
rect 43180 27010 43208 30670
rect 43364 30258 43392 31894
rect 43640 31822 43668 32302
rect 44192 31958 44220 32302
rect 44180 31952 44232 31958
rect 44180 31894 44232 31900
rect 43628 31816 43680 31822
rect 43628 31758 43680 31764
rect 44376 31754 44404 32422
rect 44468 32298 44496 32778
rect 44560 32502 44588 32966
rect 44836 32910 44864 33254
rect 44640 32904 44692 32910
rect 44640 32846 44692 32852
rect 44824 32904 44876 32910
rect 44824 32846 44876 32852
rect 44548 32496 44600 32502
rect 44548 32438 44600 32444
rect 44456 32292 44508 32298
rect 44456 32234 44508 32240
rect 44560 31958 44588 32438
rect 44652 32230 44680 32846
rect 44732 32768 44784 32774
rect 44732 32710 44784 32716
rect 44744 32230 44772 32710
rect 44916 32564 44968 32570
rect 44916 32506 44968 32512
rect 44928 32434 44956 32506
rect 45480 32434 45508 33798
rect 45664 33658 45692 33934
rect 46388 33856 46440 33862
rect 46388 33798 46440 33804
rect 45652 33652 45704 33658
rect 45652 33594 45704 33600
rect 46400 33522 46428 33798
rect 46492 33522 46520 57326
rect 50294 56604 50602 56613
rect 50294 56602 50300 56604
rect 50356 56602 50380 56604
rect 50436 56602 50460 56604
rect 50516 56602 50540 56604
rect 50596 56602 50602 56604
rect 50356 56550 50358 56602
rect 50538 56550 50540 56602
rect 50294 56548 50300 56550
rect 50356 56548 50380 56550
rect 50436 56548 50460 56550
rect 50516 56548 50540 56550
rect 50596 56548 50602 56550
rect 50294 56539 50602 56548
rect 50294 55516 50602 55525
rect 50294 55514 50300 55516
rect 50356 55514 50380 55516
rect 50436 55514 50460 55516
rect 50516 55514 50540 55516
rect 50596 55514 50602 55516
rect 50356 55462 50358 55514
rect 50538 55462 50540 55514
rect 50294 55460 50300 55462
rect 50356 55460 50380 55462
rect 50436 55460 50460 55462
rect 50516 55460 50540 55462
rect 50596 55460 50602 55462
rect 50294 55451 50602 55460
rect 50294 54428 50602 54437
rect 50294 54426 50300 54428
rect 50356 54426 50380 54428
rect 50436 54426 50460 54428
rect 50516 54426 50540 54428
rect 50596 54426 50602 54428
rect 50356 54374 50358 54426
rect 50538 54374 50540 54426
rect 50294 54372 50300 54374
rect 50356 54372 50380 54374
rect 50436 54372 50460 54374
rect 50516 54372 50540 54374
rect 50596 54372 50602 54374
rect 50294 54363 50602 54372
rect 50294 53340 50602 53349
rect 50294 53338 50300 53340
rect 50356 53338 50380 53340
rect 50436 53338 50460 53340
rect 50516 53338 50540 53340
rect 50596 53338 50602 53340
rect 50356 53286 50358 53338
rect 50538 53286 50540 53338
rect 50294 53284 50300 53286
rect 50356 53284 50380 53286
rect 50436 53284 50460 53286
rect 50516 53284 50540 53286
rect 50596 53284 50602 53286
rect 50294 53275 50602 53284
rect 58900 53100 58952 53106
rect 58900 53042 58952 53048
rect 58912 52873 58940 53042
rect 58992 52896 59044 52902
rect 58898 52864 58954 52873
rect 58992 52838 59044 52844
rect 58898 52799 58954 52808
rect 58624 52692 58676 52698
rect 58624 52634 58676 52640
rect 50294 52252 50602 52261
rect 50294 52250 50300 52252
rect 50356 52250 50380 52252
rect 50436 52250 50460 52252
rect 50516 52250 50540 52252
rect 50596 52250 50602 52252
rect 50356 52198 50358 52250
rect 50538 52198 50540 52250
rect 50294 52196 50300 52198
rect 50356 52196 50380 52198
rect 50436 52196 50460 52198
rect 50516 52196 50540 52198
rect 50596 52196 50602 52198
rect 50294 52187 50602 52196
rect 50294 51164 50602 51173
rect 50294 51162 50300 51164
rect 50356 51162 50380 51164
rect 50436 51162 50460 51164
rect 50516 51162 50540 51164
rect 50596 51162 50602 51164
rect 50356 51110 50358 51162
rect 50538 51110 50540 51162
rect 50294 51108 50300 51110
rect 50356 51108 50380 51110
rect 50436 51108 50460 51110
rect 50516 51108 50540 51110
rect 50596 51108 50602 51110
rect 50294 51099 50602 51108
rect 50294 50076 50602 50085
rect 50294 50074 50300 50076
rect 50356 50074 50380 50076
rect 50436 50074 50460 50076
rect 50516 50074 50540 50076
rect 50596 50074 50602 50076
rect 50356 50022 50358 50074
rect 50538 50022 50540 50074
rect 50294 50020 50300 50022
rect 50356 50020 50380 50022
rect 50436 50020 50460 50022
rect 50516 50020 50540 50022
rect 50596 50020 50602 50022
rect 50294 50011 50602 50020
rect 58348 49088 58400 49094
rect 58348 49030 58400 49036
rect 50294 48988 50602 48997
rect 50294 48986 50300 48988
rect 50356 48986 50380 48988
rect 50436 48986 50460 48988
rect 50516 48986 50540 48988
rect 50596 48986 50602 48988
rect 50356 48934 50358 48986
rect 50538 48934 50540 48986
rect 50294 48932 50300 48934
rect 50356 48932 50380 48934
rect 50436 48932 50460 48934
rect 50516 48932 50540 48934
rect 50596 48932 50602 48934
rect 50294 48923 50602 48932
rect 57796 48000 57848 48006
rect 57796 47942 57848 47948
rect 50294 47900 50602 47909
rect 50294 47898 50300 47900
rect 50356 47898 50380 47900
rect 50436 47898 50460 47900
rect 50516 47898 50540 47900
rect 50596 47898 50602 47900
rect 50356 47846 50358 47898
rect 50538 47846 50540 47898
rect 50294 47844 50300 47846
rect 50356 47844 50380 47846
rect 50436 47844 50460 47846
rect 50516 47844 50540 47846
rect 50596 47844 50602 47846
rect 50294 47835 50602 47844
rect 50294 46812 50602 46821
rect 50294 46810 50300 46812
rect 50356 46810 50380 46812
rect 50436 46810 50460 46812
rect 50516 46810 50540 46812
rect 50596 46810 50602 46812
rect 50356 46758 50358 46810
rect 50538 46758 50540 46810
rect 50294 46756 50300 46758
rect 50356 46756 50380 46758
rect 50436 46756 50460 46758
rect 50516 46756 50540 46758
rect 50596 46756 50602 46758
rect 50294 46747 50602 46756
rect 50294 45724 50602 45733
rect 50294 45722 50300 45724
rect 50356 45722 50380 45724
rect 50436 45722 50460 45724
rect 50516 45722 50540 45724
rect 50596 45722 50602 45724
rect 50356 45670 50358 45722
rect 50538 45670 50540 45722
rect 50294 45668 50300 45670
rect 50356 45668 50380 45670
rect 50436 45668 50460 45670
rect 50516 45668 50540 45670
rect 50596 45668 50602 45670
rect 50294 45659 50602 45668
rect 57520 44736 57572 44742
rect 57520 44678 57572 44684
rect 50294 44636 50602 44645
rect 50294 44634 50300 44636
rect 50356 44634 50380 44636
rect 50436 44634 50460 44636
rect 50516 44634 50540 44636
rect 50596 44634 50602 44636
rect 50356 44582 50358 44634
rect 50538 44582 50540 44634
rect 50294 44580 50300 44582
rect 50356 44580 50380 44582
rect 50436 44580 50460 44582
rect 50516 44580 50540 44582
rect 50596 44580 50602 44582
rect 50294 44571 50602 44580
rect 57532 43722 57560 44678
rect 57520 43716 57572 43722
rect 57520 43658 57572 43664
rect 50294 43548 50602 43557
rect 50294 43546 50300 43548
rect 50356 43546 50380 43548
rect 50436 43546 50460 43548
rect 50516 43546 50540 43548
rect 50596 43546 50602 43548
rect 50356 43494 50358 43546
rect 50538 43494 50540 43546
rect 50294 43492 50300 43494
rect 50356 43492 50380 43494
rect 50436 43492 50460 43494
rect 50516 43492 50540 43494
rect 50596 43492 50602 43494
rect 50294 43483 50602 43492
rect 57428 43240 57480 43246
rect 57428 43182 57480 43188
rect 56692 43104 56744 43110
rect 56692 43046 56744 43052
rect 56784 43104 56836 43110
rect 56784 43046 56836 43052
rect 56704 42770 56732 43046
rect 56692 42764 56744 42770
rect 56692 42706 56744 42712
rect 55680 42628 55732 42634
rect 55680 42570 55732 42576
rect 50294 42460 50602 42469
rect 50294 42458 50300 42460
rect 50356 42458 50380 42460
rect 50436 42458 50460 42460
rect 50516 42458 50540 42460
rect 50596 42458 50602 42460
rect 50356 42406 50358 42458
rect 50538 42406 50540 42458
rect 50294 42404 50300 42406
rect 50356 42404 50380 42406
rect 50436 42404 50460 42406
rect 50516 42404 50540 42406
rect 50596 42404 50602 42406
rect 50294 42395 50602 42404
rect 50294 41372 50602 41381
rect 50294 41370 50300 41372
rect 50356 41370 50380 41372
rect 50436 41370 50460 41372
rect 50516 41370 50540 41372
rect 50596 41370 50602 41372
rect 50356 41318 50358 41370
rect 50538 41318 50540 41370
rect 50294 41316 50300 41318
rect 50356 41316 50380 41318
rect 50436 41316 50460 41318
rect 50516 41316 50540 41318
rect 50596 41316 50602 41318
rect 50294 41307 50602 41316
rect 47308 40452 47360 40458
rect 47308 40394 47360 40400
rect 46388 33516 46440 33522
rect 46388 33458 46440 33464
rect 46480 33516 46532 33522
rect 46480 33458 46532 33464
rect 46020 33448 46072 33454
rect 46020 33390 46072 33396
rect 46032 33114 46060 33390
rect 46110 33144 46166 33153
rect 46020 33108 46072 33114
rect 46110 33079 46112 33088
rect 46020 33050 46072 33056
rect 46164 33079 46166 33088
rect 46112 33050 46164 33056
rect 45652 32564 45704 32570
rect 45652 32506 45704 32512
rect 44916 32428 44968 32434
rect 44916 32370 44968 32376
rect 45468 32428 45520 32434
rect 45468 32370 45520 32376
rect 45560 32360 45612 32366
rect 45388 32308 45560 32314
rect 45388 32302 45612 32308
rect 45388 32286 45600 32302
rect 44640 32224 44692 32230
rect 44640 32166 44692 32172
rect 44732 32224 44784 32230
rect 44732 32166 44784 32172
rect 44652 32026 44680 32166
rect 44640 32020 44692 32026
rect 44640 31962 44692 31968
rect 44548 31952 44600 31958
rect 44548 31894 44600 31900
rect 44640 31816 44692 31822
rect 44640 31758 44692 31764
rect 44364 31748 44416 31754
rect 44364 31690 44416 31696
rect 44088 31272 44140 31278
rect 44088 31214 44140 31220
rect 44100 30938 44128 31214
rect 44088 30932 44140 30938
rect 44088 30874 44140 30880
rect 43720 30728 43772 30734
rect 43720 30670 43772 30676
rect 43732 30394 43760 30670
rect 43720 30388 43772 30394
rect 43720 30330 43772 30336
rect 43352 30252 43404 30258
rect 43352 30194 43404 30200
rect 44180 30252 44232 30258
rect 44180 30194 44232 30200
rect 43996 30184 44048 30190
rect 43996 30126 44048 30132
rect 43444 30048 43496 30054
rect 43444 29990 43496 29996
rect 43536 30048 43588 30054
rect 43536 29990 43588 29996
rect 43456 29782 43484 29990
rect 43548 29850 43576 29990
rect 43536 29844 43588 29850
rect 43536 29786 43588 29792
rect 43444 29776 43496 29782
rect 43444 29718 43496 29724
rect 44008 29646 44036 30126
rect 44192 29850 44220 30194
rect 44180 29844 44232 29850
rect 44180 29786 44232 29792
rect 43996 29640 44048 29646
rect 43996 29582 44048 29588
rect 43628 29572 43680 29578
rect 43628 29514 43680 29520
rect 44548 29572 44600 29578
rect 44548 29514 44600 29520
rect 43536 29504 43588 29510
rect 43536 29446 43588 29452
rect 43548 29238 43576 29446
rect 43536 29232 43588 29238
rect 43536 29174 43588 29180
rect 43260 28484 43312 28490
rect 43260 28426 43312 28432
rect 43272 28218 43300 28426
rect 43640 28218 43668 29514
rect 44088 29028 44140 29034
rect 44088 28970 44140 28976
rect 43260 28212 43312 28218
rect 43260 28154 43312 28160
rect 43628 28212 43680 28218
rect 43628 28154 43680 28160
rect 43444 28076 43496 28082
rect 43444 28018 43496 28024
rect 43456 27674 43484 28018
rect 43628 28008 43680 28014
rect 43548 27956 43628 27962
rect 43548 27950 43680 27956
rect 43548 27934 43668 27950
rect 43444 27668 43496 27674
rect 43444 27610 43496 27616
rect 43548 27334 43576 27934
rect 43720 27668 43772 27674
rect 43720 27610 43772 27616
rect 43536 27328 43588 27334
rect 43536 27270 43588 27276
rect 43548 27062 43576 27270
rect 43732 27062 43760 27610
rect 43904 27532 43956 27538
rect 43904 27474 43956 27480
rect 42996 26982 43208 27010
rect 43352 27056 43404 27062
rect 43352 26998 43404 27004
rect 43536 27056 43588 27062
rect 43536 26998 43588 27004
rect 43720 27056 43772 27062
rect 43720 26998 43772 27004
rect 43260 26988 43312 26994
rect 43260 26930 43312 26936
rect 42800 26580 42852 26586
rect 42800 26522 42852 26528
rect 42892 25900 42944 25906
rect 42892 25842 42944 25848
rect 42708 25696 42760 25702
rect 42708 25638 42760 25644
rect 42616 25492 42668 25498
rect 42616 25434 42668 25440
rect 42524 25356 42576 25362
rect 42524 25298 42576 25304
rect 42720 24954 42748 25638
rect 42800 25220 42852 25226
rect 42800 25162 42852 25168
rect 42812 24954 42840 25162
rect 42904 25158 42932 25842
rect 42892 25152 42944 25158
rect 42892 25094 42944 25100
rect 42708 24948 42760 24954
rect 42708 24890 42760 24896
rect 42800 24948 42852 24954
rect 42800 24890 42852 24896
rect 42904 24886 42932 25094
rect 42892 24880 42944 24886
rect 42892 24822 42944 24828
rect 42248 24608 42300 24614
rect 42248 24550 42300 24556
rect 42156 24268 42208 24274
rect 42156 24210 42208 24216
rect 42260 23662 42288 24550
rect 42708 24200 42760 24206
rect 42708 24142 42760 24148
rect 42248 23656 42300 23662
rect 42248 23598 42300 23604
rect 42260 22982 42288 23598
rect 42720 23322 42748 24142
rect 42708 23316 42760 23322
rect 42708 23258 42760 23264
rect 42248 22976 42300 22982
rect 42248 22918 42300 22924
rect 41788 19848 41840 19854
rect 41788 19790 41840 19796
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 38660 18080 38712 18086
rect 38660 18022 38712 18028
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 38672 2446 38700 18022
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12636 1306 12664 2382
rect 17604 1306 17632 2382
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 22572 1306 22600 2382
rect 27712 2372 27764 2378
rect 27712 2314 27764 2320
rect 32404 2372 32456 2378
rect 32404 2314 32456 2320
rect 37372 2372 37424 2378
rect 37372 2314 37424 2320
rect 27724 1442 27752 2314
rect 12544 1278 12664 1306
rect 17512 1278 17632 1306
rect 22480 1278 22600 1306
rect 27448 1414 27752 1442
rect 12544 800 12572 1278
rect 17512 800 17540 1278
rect 22480 800 22508 1278
rect 27448 800 27476 1414
rect 32416 800 32444 2314
rect 37384 800 37412 2314
rect 42260 2038 42288 22918
rect 42432 22432 42484 22438
rect 42432 22374 42484 22380
rect 42444 22234 42472 22374
rect 42720 22234 42748 23258
rect 43272 22778 43300 26930
rect 43364 26246 43392 26998
rect 43916 26994 43944 27474
rect 43996 27056 44048 27062
rect 43996 26998 44048 27004
rect 43904 26988 43956 26994
rect 43904 26930 43956 26936
rect 44008 26382 44036 26998
rect 43904 26376 43956 26382
rect 43904 26318 43956 26324
rect 43996 26376 44048 26382
rect 43996 26318 44048 26324
rect 43352 26240 43404 26246
rect 43352 26182 43404 26188
rect 43812 24812 43864 24818
rect 43812 24754 43864 24760
rect 43824 24410 43852 24754
rect 43812 24404 43864 24410
rect 43812 24346 43864 24352
rect 43444 24064 43496 24070
rect 43444 24006 43496 24012
rect 43456 23798 43484 24006
rect 43824 23866 43852 24346
rect 43916 24274 43944 26318
rect 44100 25770 44128 28970
rect 44456 26376 44508 26382
rect 44454 26344 44456 26353
rect 44508 26344 44510 26353
rect 44376 26302 44454 26330
rect 44088 25764 44140 25770
rect 44088 25706 44140 25712
rect 44088 25492 44140 25498
rect 44088 25434 44140 25440
rect 44100 25294 44128 25434
rect 44088 25288 44140 25294
rect 44088 25230 44140 25236
rect 43996 24676 44048 24682
rect 43996 24618 44048 24624
rect 43904 24268 43956 24274
rect 43904 24210 43956 24216
rect 43916 24138 43944 24210
rect 43904 24132 43956 24138
rect 43904 24074 43956 24080
rect 44008 24120 44036 24618
rect 44100 24342 44128 25230
rect 44376 24818 44404 26302
rect 44454 26279 44510 26288
rect 44456 25900 44508 25906
rect 44456 25842 44508 25848
rect 44468 24818 44496 25842
rect 44560 24818 44588 29514
rect 44652 28762 44680 31758
rect 45388 31754 45416 32286
rect 45560 32224 45612 32230
rect 45560 32166 45612 32172
rect 45192 31748 45416 31754
rect 45244 31726 45416 31748
rect 45192 31690 45244 31696
rect 45204 31346 45232 31690
rect 45572 31482 45600 32166
rect 45664 31822 45692 32506
rect 46204 32292 46256 32298
rect 46204 32234 46256 32240
rect 45652 31816 45704 31822
rect 45652 31758 45704 31764
rect 45560 31476 45612 31482
rect 45560 31418 45612 31424
rect 45192 31340 45244 31346
rect 45192 31282 45244 31288
rect 45100 30048 45152 30054
rect 45100 29990 45152 29996
rect 44824 29640 44876 29646
rect 44824 29582 44876 29588
rect 44732 29096 44784 29102
rect 44732 29038 44784 29044
rect 44640 28756 44692 28762
rect 44640 28698 44692 28704
rect 44652 28218 44680 28698
rect 44640 28212 44692 28218
rect 44640 28154 44692 28160
rect 44640 28008 44692 28014
rect 44640 27950 44692 27956
rect 44180 24812 44232 24818
rect 44180 24754 44232 24760
rect 44364 24812 44416 24818
rect 44364 24754 44416 24760
rect 44456 24812 44508 24818
rect 44456 24754 44508 24760
rect 44548 24812 44600 24818
rect 44548 24754 44600 24760
rect 44088 24336 44140 24342
rect 44088 24278 44140 24284
rect 44088 24132 44140 24138
rect 44008 24092 44088 24120
rect 43812 23860 43864 23866
rect 43812 23802 43864 23808
rect 43444 23792 43496 23798
rect 43444 23734 43496 23740
rect 43260 22772 43312 22778
rect 43260 22714 43312 22720
rect 43168 22636 43220 22642
rect 43168 22578 43220 22584
rect 42984 22568 43036 22574
rect 42984 22510 43036 22516
rect 42432 22228 42484 22234
rect 42708 22228 42760 22234
rect 42432 22170 42484 22176
rect 42628 22188 42708 22216
rect 42628 22030 42656 22188
rect 42708 22170 42760 22176
rect 42616 22024 42668 22030
rect 42616 21966 42668 21972
rect 42892 22024 42944 22030
rect 42892 21966 42944 21972
rect 42904 21690 42932 21966
rect 42996 21690 43024 22510
rect 43180 21962 43208 22578
rect 43456 22574 43484 23734
rect 44008 23730 44036 24092
rect 44088 24074 44140 24080
rect 43996 23724 44048 23730
rect 43996 23666 44048 23672
rect 44008 22778 44036 23666
rect 44192 23202 44220 24754
rect 44272 24064 44324 24070
rect 44272 24006 44324 24012
rect 44100 23174 44220 23202
rect 43996 22772 44048 22778
rect 43996 22714 44048 22720
rect 43444 22568 43496 22574
rect 43444 22510 43496 22516
rect 43444 22432 43496 22438
rect 43444 22374 43496 22380
rect 43812 22432 43864 22438
rect 43812 22374 43864 22380
rect 43168 21956 43220 21962
rect 43168 21898 43220 21904
rect 43180 21690 43208 21898
rect 42892 21684 42944 21690
rect 42892 21626 42944 21632
rect 42984 21684 43036 21690
rect 42984 21626 43036 21632
rect 43168 21684 43220 21690
rect 43168 21626 43220 21632
rect 42892 21344 42944 21350
rect 42892 21286 42944 21292
rect 42904 21146 42932 21286
rect 42892 21140 42944 21146
rect 42892 21082 42944 21088
rect 43456 20942 43484 22374
rect 43536 21888 43588 21894
rect 43536 21830 43588 21836
rect 43548 21690 43576 21830
rect 43536 21684 43588 21690
rect 43536 21626 43588 21632
rect 43824 21350 43852 22374
rect 43996 21888 44048 21894
rect 43996 21830 44048 21836
rect 44008 21554 44036 21830
rect 44100 21554 44128 23174
rect 44180 23112 44232 23118
rect 44180 23054 44232 23060
rect 44192 22098 44220 23054
rect 44284 22642 44312 24006
rect 44652 23594 44680 27950
rect 44744 27334 44772 29038
rect 44836 27470 44864 29582
rect 45112 29306 45140 29990
rect 45100 29300 45152 29306
rect 45100 29242 45152 29248
rect 45204 28694 45232 31282
rect 45664 30954 45692 31758
rect 46216 31414 46244 32234
rect 46204 31408 46256 31414
rect 46204 31350 46256 31356
rect 45836 31272 45888 31278
rect 45836 31214 45888 31220
rect 45744 31136 45796 31142
rect 45744 31078 45796 31084
rect 45572 30926 45692 30954
rect 45572 30734 45600 30926
rect 45756 30870 45784 31078
rect 45744 30864 45796 30870
rect 45744 30806 45796 30812
rect 45848 30802 45876 31214
rect 45928 31136 45980 31142
rect 45928 31078 45980 31084
rect 45940 30938 45968 31078
rect 45928 30932 45980 30938
rect 45928 30874 45980 30880
rect 45836 30796 45888 30802
rect 45836 30738 45888 30744
rect 45560 30728 45612 30734
rect 45560 30670 45612 30676
rect 45652 30728 45704 30734
rect 45652 30670 45704 30676
rect 45664 29714 45692 30670
rect 45744 30660 45796 30666
rect 45744 30602 45796 30608
rect 45756 30394 45784 30602
rect 45744 30388 45796 30394
rect 45744 30330 45796 30336
rect 45744 30184 45796 30190
rect 45744 30126 45796 30132
rect 45756 30054 45784 30126
rect 46020 30116 46072 30122
rect 46020 30058 46072 30064
rect 45744 30048 45796 30054
rect 45744 29990 45796 29996
rect 45652 29708 45704 29714
rect 45652 29650 45704 29656
rect 45664 29306 45692 29650
rect 45652 29300 45704 29306
rect 45652 29242 45704 29248
rect 45560 28960 45612 28966
rect 45560 28902 45612 28908
rect 45192 28688 45244 28694
rect 45192 28630 45244 28636
rect 45572 28558 45600 28902
rect 45664 28626 45692 29242
rect 45652 28620 45704 28626
rect 45652 28562 45704 28568
rect 45192 28552 45244 28558
rect 45192 28494 45244 28500
rect 45560 28552 45612 28558
rect 45560 28494 45612 28500
rect 45204 28218 45232 28494
rect 45192 28212 45244 28218
rect 45192 28154 45244 28160
rect 44916 27600 44968 27606
rect 44916 27542 44968 27548
rect 44824 27464 44876 27470
rect 44824 27406 44876 27412
rect 44732 27328 44784 27334
rect 44732 27270 44784 27276
rect 44744 25140 44772 27270
rect 44928 27062 44956 27542
rect 45652 27464 45704 27470
rect 45652 27406 45704 27412
rect 45284 27396 45336 27402
rect 45284 27338 45336 27344
rect 44916 27056 44968 27062
rect 44916 26998 44968 27004
rect 44824 26512 44876 26518
rect 44824 26454 44876 26460
rect 44836 25294 44864 26454
rect 45192 26376 45244 26382
rect 45192 26318 45244 26324
rect 45204 25838 45232 26318
rect 45296 26042 45324 27338
rect 45664 26450 45692 27406
rect 45756 27334 45784 29990
rect 46032 27606 46060 30058
rect 46112 29096 46164 29102
rect 46112 29038 46164 29044
rect 46124 28762 46152 29038
rect 46112 28756 46164 28762
rect 46112 28698 46164 28704
rect 46400 28150 46428 33458
rect 46492 33114 46520 33458
rect 46480 33108 46532 33114
rect 46480 33050 46532 33056
rect 46664 32496 46716 32502
rect 46664 32438 46716 32444
rect 46676 32366 46704 32438
rect 46664 32360 46716 32366
rect 46664 32302 46716 32308
rect 47032 32360 47084 32366
rect 47032 32302 47084 32308
rect 46676 30598 46704 32302
rect 47044 32026 47072 32302
rect 47032 32020 47084 32026
rect 47032 31962 47084 31968
rect 47124 32020 47176 32026
rect 47124 31962 47176 31968
rect 46756 31816 46808 31822
rect 46756 31758 46808 31764
rect 46768 31278 46796 31758
rect 47136 31754 47164 31962
rect 47320 31822 47348 40394
rect 50294 40284 50602 40293
rect 50294 40282 50300 40284
rect 50356 40282 50380 40284
rect 50436 40282 50460 40284
rect 50516 40282 50540 40284
rect 50596 40282 50602 40284
rect 50356 40230 50358 40282
rect 50538 40230 50540 40282
rect 50294 40228 50300 40230
rect 50356 40228 50380 40230
rect 50436 40228 50460 40230
rect 50516 40228 50540 40230
rect 50596 40228 50602 40230
rect 50294 40219 50602 40228
rect 50294 39196 50602 39205
rect 50294 39194 50300 39196
rect 50356 39194 50380 39196
rect 50436 39194 50460 39196
rect 50516 39194 50540 39196
rect 50596 39194 50602 39196
rect 50356 39142 50358 39194
rect 50538 39142 50540 39194
rect 50294 39140 50300 39142
rect 50356 39140 50380 39142
rect 50436 39140 50460 39142
rect 50516 39140 50540 39142
rect 50596 39140 50602 39142
rect 50294 39131 50602 39140
rect 50294 38108 50602 38117
rect 50294 38106 50300 38108
rect 50356 38106 50380 38108
rect 50436 38106 50460 38108
rect 50516 38106 50540 38108
rect 50596 38106 50602 38108
rect 50356 38054 50358 38106
rect 50538 38054 50540 38106
rect 50294 38052 50300 38054
rect 50356 38052 50380 38054
rect 50436 38052 50460 38054
rect 50516 38052 50540 38054
rect 50596 38052 50602 38054
rect 50294 38043 50602 38052
rect 50294 37020 50602 37029
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36955 50602 36964
rect 50294 35932 50602 35941
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35867 50602 35876
rect 55312 34944 55364 34950
rect 55312 34886 55364 34892
rect 50294 34844 50602 34853
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34779 50602 34788
rect 49700 34604 49752 34610
rect 49700 34546 49752 34552
rect 49712 33674 49740 34546
rect 50804 34536 50856 34542
rect 50804 34478 50856 34484
rect 51448 34536 51500 34542
rect 51448 34478 51500 34484
rect 50816 34202 50844 34478
rect 51172 34400 51224 34406
rect 51172 34342 51224 34348
rect 50804 34196 50856 34202
rect 50804 34138 50856 34144
rect 50160 33992 50212 33998
rect 50160 33934 50212 33940
rect 49528 33658 49740 33674
rect 50172 33658 50200 33934
rect 50294 33756 50602 33765
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33691 50602 33700
rect 51184 33674 51212 34342
rect 51264 33924 51316 33930
rect 51264 33866 51316 33872
rect 49516 33652 49740 33658
rect 49568 33646 49740 33652
rect 49516 33594 49568 33600
rect 49240 33584 49292 33590
rect 49240 33526 49292 33532
rect 47400 33516 47452 33522
rect 47400 33458 47452 33464
rect 47412 32434 47440 33458
rect 47860 33448 47912 33454
rect 47860 33390 47912 33396
rect 47872 33114 47900 33390
rect 47860 33108 47912 33114
rect 47860 33050 47912 33056
rect 49252 32910 49280 33526
rect 47676 32904 47728 32910
rect 47676 32846 47728 32852
rect 48320 32904 48372 32910
rect 48320 32846 48372 32852
rect 49240 32904 49292 32910
rect 49240 32846 49292 32852
rect 47688 32434 47716 32846
rect 47400 32428 47452 32434
rect 47400 32370 47452 32376
rect 47676 32428 47728 32434
rect 47676 32370 47728 32376
rect 47308 31816 47360 31822
rect 47308 31758 47360 31764
rect 46952 31726 47164 31754
rect 46952 31686 46980 31726
rect 46940 31680 46992 31686
rect 46940 31622 46992 31628
rect 47032 31680 47084 31686
rect 47032 31622 47084 31628
rect 46756 31272 46808 31278
rect 46756 31214 46808 31220
rect 46664 30592 46716 30598
rect 46664 30534 46716 30540
rect 46572 30388 46624 30394
rect 46572 30330 46624 30336
rect 46584 29646 46612 30330
rect 46572 29640 46624 29646
rect 46572 29582 46624 29588
rect 46572 29504 46624 29510
rect 46572 29446 46624 29452
rect 46848 29504 46900 29510
rect 46848 29446 46900 29452
rect 46584 28626 46612 29446
rect 46860 29306 46888 29446
rect 46848 29300 46900 29306
rect 46848 29242 46900 29248
rect 46572 28620 46624 28626
rect 46572 28562 46624 28568
rect 46584 28490 46612 28562
rect 46572 28484 46624 28490
rect 46572 28426 46624 28432
rect 46388 28144 46440 28150
rect 46388 28086 46440 28092
rect 46400 27674 46428 28086
rect 46388 27668 46440 27674
rect 46388 27610 46440 27616
rect 45836 27600 45888 27606
rect 45836 27542 45888 27548
rect 46020 27600 46072 27606
rect 46020 27542 46072 27548
rect 45744 27328 45796 27334
rect 45744 27270 45796 27276
rect 45756 26994 45784 27270
rect 45744 26988 45796 26994
rect 45744 26930 45796 26936
rect 45848 26858 45876 27542
rect 45928 27464 45980 27470
rect 45928 27406 45980 27412
rect 45940 27062 45968 27406
rect 45928 27056 45980 27062
rect 45928 26998 45980 27004
rect 46032 26994 46060 27542
rect 46480 27464 46532 27470
rect 46480 27406 46532 27412
rect 46110 27160 46166 27169
rect 46492 27130 46520 27406
rect 46110 27095 46112 27104
rect 46164 27095 46166 27104
rect 46480 27124 46532 27130
rect 46112 27066 46164 27072
rect 46480 27066 46532 27072
rect 46020 26988 46072 26994
rect 46572 26988 46624 26994
rect 46020 26930 46072 26936
rect 46400 26948 46572 26976
rect 46032 26858 46060 26930
rect 45836 26852 45888 26858
rect 45836 26794 45888 26800
rect 46020 26852 46072 26858
rect 46020 26794 46072 26800
rect 45652 26444 45704 26450
rect 45652 26386 45704 26392
rect 45376 26366 45428 26372
rect 45428 26314 45600 26330
rect 45376 26308 45600 26314
rect 45388 26302 45600 26308
rect 45284 26036 45336 26042
rect 45284 25978 45336 25984
rect 45572 25906 45600 26302
rect 45744 26240 45796 26246
rect 45744 26182 45796 26188
rect 45560 25900 45612 25906
rect 45560 25842 45612 25848
rect 45192 25832 45244 25838
rect 45192 25774 45244 25780
rect 44824 25288 44876 25294
rect 44824 25230 44876 25236
rect 45008 25152 45060 25158
rect 44744 25112 44864 25140
rect 44640 23588 44692 23594
rect 44640 23530 44692 23536
rect 44364 23520 44416 23526
rect 44364 23462 44416 23468
rect 44272 22636 44324 22642
rect 44272 22578 44324 22584
rect 44180 22092 44232 22098
rect 44180 22034 44232 22040
rect 44192 21690 44220 22034
rect 44284 22030 44312 22578
rect 44272 22024 44324 22030
rect 44272 21966 44324 21972
rect 44180 21684 44232 21690
rect 44180 21626 44232 21632
rect 44376 21554 44404 23462
rect 44836 22506 44864 25112
rect 45008 25094 45060 25100
rect 45020 24954 45048 25094
rect 45008 24948 45060 24954
rect 45008 24890 45060 24896
rect 45204 24818 45232 25774
rect 45284 25288 45336 25294
rect 45284 25230 45336 25236
rect 45192 24812 45244 24818
rect 45192 24754 45244 24760
rect 45008 24744 45060 24750
rect 45008 24686 45060 24692
rect 45020 24410 45048 24686
rect 45008 24404 45060 24410
rect 45008 24346 45060 24352
rect 45296 24206 45324 25230
rect 45572 25226 45600 25842
rect 45560 25220 45612 25226
rect 45560 25162 45612 25168
rect 45756 24954 45784 26182
rect 45744 24948 45796 24954
rect 45744 24890 45796 24896
rect 45376 24812 45428 24818
rect 45376 24754 45428 24760
rect 45388 24614 45416 24754
rect 45848 24682 45876 26794
rect 46400 26586 46428 26948
rect 46572 26930 46624 26936
rect 46388 26580 46440 26586
rect 46388 26522 46440 26528
rect 46400 26382 46428 26522
rect 46952 26382 46980 31622
rect 47044 31482 47072 31622
rect 47136 31482 47164 31726
rect 47216 31680 47268 31686
rect 47216 31622 47268 31628
rect 47032 31476 47084 31482
rect 47032 31418 47084 31424
rect 47124 31476 47176 31482
rect 47124 31418 47176 31424
rect 47124 31136 47176 31142
rect 47124 31078 47176 31084
rect 47032 30184 47084 30190
rect 47032 30126 47084 30132
rect 47044 29850 47072 30126
rect 47136 29850 47164 31078
rect 47228 30666 47256 31622
rect 47412 30802 47440 32370
rect 47688 31754 47716 32370
rect 48332 31958 48360 32846
rect 48964 32836 49016 32842
rect 48964 32778 49016 32784
rect 48596 32020 48648 32026
rect 48596 31962 48648 31968
rect 48320 31952 48372 31958
rect 48320 31894 48372 31900
rect 47676 31748 47728 31754
rect 47676 31690 47728 31696
rect 48320 31340 48372 31346
rect 48320 31282 48372 31288
rect 47400 30796 47452 30802
rect 47400 30738 47452 30744
rect 47216 30660 47268 30666
rect 47216 30602 47268 30608
rect 47308 30592 47360 30598
rect 47308 30534 47360 30540
rect 47320 30326 47348 30534
rect 47308 30320 47360 30326
rect 47308 30262 47360 30268
rect 47032 29844 47084 29850
rect 47032 29786 47084 29792
rect 47124 29844 47176 29850
rect 47124 29786 47176 29792
rect 47320 29646 47348 30262
rect 47412 29714 47440 30738
rect 47860 30048 47912 30054
rect 47860 29990 47912 29996
rect 47872 29714 47900 29990
rect 47400 29708 47452 29714
rect 47400 29650 47452 29656
rect 47860 29708 47912 29714
rect 47860 29650 47912 29656
rect 47308 29640 47360 29646
rect 47308 29582 47360 29588
rect 48228 29096 48280 29102
rect 48228 29038 48280 29044
rect 47124 28960 47176 28966
rect 47124 28902 47176 28908
rect 47136 28150 47164 28902
rect 48136 28756 48188 28762
rect 48136 28698 48188 28704
rect 48044 28484 48096 28490
rect 48044 28426 48096 28432
rect 47124 28144 47176 28150
rect 47124 28086 47176 28092
rect 47582 28112 47638 28121
rect 47216 28076 47268 28082
rect 47582 28047 47584 28056
rect 47216 28018 47268 28024
rect 47636 28047 47638 28056
rect 47860 28076 47912 28082
rect 47584 28018 47636 28024
rect 47860 28018 47912 28024
rect 47124 28008 47176 28014
rect 47124 27950 47176 27956
rect 47136 26450 47164 27950
rect 47228 27062 47256 28018
rect 47768 27940 47820 27946
rect 47768 27882 47820 27888
rect 47780 27470 47808 27882
rect 47768 27464 47820 27470
rect 47768 27406 47820 27412
rect 47216 27056 47268 27062
rect 47216 26998 47268 27004
rect 47676 26988 47728 26994
rect 47676 26930 47728 26936
rect 47308 26852 47360 26858
rect 47308 26794 47360 26800
rect 47124 26444 47176 26450
rect 47124 26386 47176 26392
rect 47320 26382 47348 26794
rect 47584 26784 47636 26790
rect 47584 26726 47636 26732
rect 46388 26376 46440 26382
rect 46388 26318 46440 26324
rect 46940 26376 46992 26382
rect 46940 26318 46992 26324
rect 47308 26376 47360 26382
rect 47308 26318 47360 26324
rect 46480 26308 46532 26314
rect 46480 26250 46532 26256
rect 46020 26036 46072 26042
rect 46020 25978 46072 25984
rect 45928 25968 45980 25974
rect 45928 25910 45980 25916
rect 45940 25294 45968 25910
rect 46032 25294 46060 25978
rect 46492 25838 46520 26250
rect 46848 26240 46900 26246
rect 46848 26182 46900 26188
rect 46480 25832 46532 25838
rect 46480 25774 46532 25780
rect 46296 25764 46348 25770
rect 46296 25706 46348 25712
rect 46308 25294 46336 25706
rect 46860 25362 46888 26182
rect 46940 26036 46992 26042
rect 46940 25978 46992 25984
rect 46952 25362 46980 25978
rect 47308 25492 47360 25498
rect 47308 25434 47360 25440
rect 46848 25356 46900 25362
rect 46848 25298 46900 25304
rect 46949 25356 47001 25362
rect 46949 25298 47001 25304
rect 45928 25288 45980 25294
rect 45928 25230 45980 25236
rect 46020 25288 46072 25294
rect 46020 25230 46072 25236
rect 46296 25288 46348 25294
rect 46296 25230 46348 25236
rect 47032 25220 47084 25226
rect 47032 25162 47084 25168
rect 46204 25152 46256 25158
rect 46204 25094 46256 25100
rect 46388 25152 46440 25158
rect 46388 25094 46440 25100
rect 46216 24886 46244 25094
rect 46204 24880 46256 24886
rect 46204 24822 46256 24828
rect 45652 24676 45704 24682
rect 45652 24618 45704 24624
rect 45836 24676 45888 24682
rect 45836 24618 45888 24624
rect 45376 24608 45428 24614
rect 45376 24550 45428 24556
rect 45468 24608 45520 24614
rect 45468 24550 45520 24556
rect 45480 24410 45508 24550
rect 45468 24404 45520 24410
rect 45468 24346 45520 24352
rect 45664 24206 45692 24618
rect 46216 24614 46244 24822
rect 46400 24818 46428 25094
rect 46768 24908 46980 24936
rect 46388 24812 46440 24818
rect 46388 24754 46440 24760
rect 46664 24812 46716 24818
rect 46768 24800 46796 24908
rect 46716 24772 46796 24800
rect 46664 24754 46716 24760
rect 46204 24608 46256 24614
rect 46204 24550 46256 24556
rect 45284 24200 45336 24206
rect 45284 24142 45336 24148
rect 45652 24200 45704 24206
rect 45652 24142 45704 24148
rect 45100 24132 45152 24138
rect 45100 24074 45152 24080
rect 45112 23526 45140 24074
rect 46572 23656 46624 23662
rect 46572 23598 46624 23604
rect 45100 23520 45152 23526
rect 45100 23462 45152 23468
rect 45928 23520 45980 23526
rect 45928 23462 45980 23468
rect 45284 23044 45336 23050
rect 45284 22986 45336 22992
rect 45296 22778 45324 22986
rect 45284 22772 45336 22778
rect 45284 22714 45336 22720
rect 45940 22574 45968 23462
rect 46584 22778 46612 23598
rect 46664 23248 46716 23254
rect 46664 23190 46716 23196
rect 46572 22772 46624 22778
rect 46572 22714 46624 22720
rect 45928 22568 45980 22574
rect 45928 22510 45980 22516
rect 44824 22500 44876 22506
rect 44824 22442 44876 22448
rect 44548 21956 44600 21962
rect 44548 21898 44600 21904
rect 44560 21622 44588 21898
rect 44732 21888 44784 21894
rect 44732 21830 44784 21836
rect 44744 21622 44772 21830
rect 44548 21616 44600 21622
rect 44548 21558 44600 21564
rect 44732 21616 44784 21622
rect 44732 21558 44784 21564
rect 43996 21548 44048 21554
rect 43996 21490 44048 21496
rect 44088 21548 44140 21554
rect 44088 21490 44140 21496
rect 44364 21548 44416 21554
rect 44364 21490 44416 21496
rect 43812 21344 43864 21350
rect 43812 21286 43864 21292
rect 44008 21010 44036 21490
rect 43996 21004 44048 21010
rect 43996 20946 44048 20952
rect 43444 20936 43496 20942
rect 43444 20878 43496 20884
rect 44100 20874 44128 21490
rect 44376 21146 44404 21490
rect 44732 21412 44784 21418
rect 44732 21354 44784 21360
rect 44640 21344 44692 21350
rect 44640 21286 44692 21292
rect 44364 21140 44416 21146
rect 44364 21082 44416 21088
rect 44652 20942 44680 21286
rect 44744 21146 44772 21354
rect 44732 21140 44784 21146
rect 44732 21082 44784 21088
rect 44640 20936 44692 20942
rect 44640 20878 44692 20884
rect 44088 20868 44140 20874
rect 44088 20810 44140 20816
rect 42616 19304 42668 19310
rect 42616 19246 42668 19252
rect 42628 2650 42656 19246
rect 44836 16046 44864 22442
rect 45652 22024 45704 22030
rect 45652 21966 45704 21972
rect 45468 21684 45520 21690
rect 45468 21626 45520 21632
rect 45480 21010 45508 21626
rect 45664 21146 45692 21966
rect 46204 21888 46256 21894
rect 46204 21830 46256 21836
rect 46216 21622 46244 21830
rect 46676 21690 46704 23190
rect 46768 22642 46796 24772
rect 46952 24732 46980 24908
rect 47044 24886 47072 25162
rect 47032 24880 47084 24886
rect 47032 24822 47084 24828
rect 47216 24812 47268 24818
rect 47216 24754 47268 24760
rect 46952 24704 47164 24732
rect 47136 24614 47164 24704
rect 47124 24608 47176 24614
rect 47124 24550 47176 24556
rect 47124 24404 47176 24410
rect 47124 24346 47176 24352
rect 46940 23044 46992 23050
rect 46940 22986 46992 22992
rect 46952 22778 46980 22986
rect 47032 22976 47084 22982
rect 47032 22918 47084 22924
rect 47044 22778 47072 22918
rect 46940 22772 46992 22778
rect 46940 22714 46992 22720
rect 47032 22772 47084 22778
rect 47032 22714 47084 22720
rect 46756 22636 46808 22642
rect 46756 22578 46808 22584
rect 47136 22030 47164 24346
rect 47228 24070 47256 24754
rect 47216 24064 47268 24070
rect 47216 24006 47268 24012
rect 47228 22506 47256 24006
rect 47320 23322 47348 25434
rect 47400 25152 47452 25158
rect 47400 25094 47452 25100
rect 47412 24818 47440 25094
rect 47400 24812 47452 24818
rect 47400 24754 47452 24760
rect 47492 24744 47544 24750
rect 47492 24686 47544 24692
rect 47504 24138 47532 24686
rect 47596 24410 47624 26726
rect 47688 26246 47716 26930
rect 47676 26240 47728 26246
rect 47676 26182 47728 26188
rect 47688 25838 47716 26182
rect 47676 25832 47728 25838
rect 47676 25774 47728 25780
rect 47676 24880 47728 24886
rect 47676 24822 47728 24828
rect 47584 24404 47636 24410
rect 47584 24346 47636 24352
rect 47688 24206 47716 24822
rect 47676 24200 47728 24206
rect 47676 24142 47728 24148
rect 47492 24132 47544 24138
rect 47492 24074 47544 24080
rect 47688 24070 47716 24142
rect 47676 24064 47728 24070
rect 47676 24006 47728 24012
rect 47780 23882 47808 27406
rect 47872 26586 47900 28018
rect 47952 27940 48004 27946
rect 47952 27882 48004 27888
rect 47964 27674 47992 27882
rect 47952 27668 48004 27674
rect 47952 27610 48004 27616
rect 47860 26580 47912 26586
rect 47860 26522 47912 26528
rect 47872 25770 47900 26522
rect 47964 25906 47992 27610
rect 48056 26382 48084 28426
rect 48148 27878 48176 28698
rect 48240 28422 48268 29038
rect 48332 28762 48360 31282
rect 48412 31136 48464 31142
rect 48412 31078 48464 31084
rect 48504 31136 48556 31142
rect 48504 31078 48556 31084
rect 48424 30258 48452 31078
rect 48516 30938 48544 31078
rect 48504 30932 48556 30938
rect 48504 30874 48556 30880
rect 48412 30252 48464 30258
rect 48412 30194 48464 30200
rect 48320 28756 48372 28762
rect 48320 28698 48372 28704
rect 48332 28626 48360 28698
rect 48320 28620 48372 28626
rect 48320 28562 48372 28568
rect 48228 28416 48280 28422
rect 48228 28358 48280 28364
rect 48240 28014 48268 28358
rect 48228 28008 48280 28014
rect 48228 27950 48280 27956
rect 48136 27872 48188 27878
rect 48136 27814 48188 27820
rect 48228 27872 48280 27878
rect 48228 27814 48280 27820
rect 48148 27470 48176 27814
rect 48136 27464 48188 27470
rect 48136 27406 48188 27412
rect 48240 27282 48268 27814
rect 48608 27470 48636 31962
rect 48976 31890 49004 32778
rect 49252 32434 49280 32846
rect 49240 32428 49292 32434
rect 49240 32370 49292 32376
rect 49056 32224 49108 32230
rect 49056 32166 49108 32172
rect 49516 32224 49568 32230
rect 49516 32166 49568 32172
rect 49068 31958 49096 32166
rect 49056 31952 49108 31958
rect 49056 31894 49108 31900
rect 48964 31884 49016 31890
rect 48964 31826 49016 31832
rect 48976 31754 49004 31826
rect 48884 31726 49004 31754
rect 48884 31278 48912 31726
rect 48964 31680 49016 31686
rect 48964 31622 49016 31628
rect 48872 31272 48924 31278
rect 48872 31214 48924 31220
rect 48688 31136 48740 31142
rect 48688 31078 48740 31084
rect 48780 31136 48832 31142
rect 48780 31078 48832 31084
rect 48700 29306 48728 31078
rect 48792 30938 48820 31078
rect 48780 30932 48832 30938
rect 48780 30874 48832 30880
rect 48976 30326 49004 31622
rect 48964 30320 49016 30326
rect 48964 30262 49016 30268
rect 48976 29714 49004 30262
rect 48964 29708 49016 29714
rect 48964 29650 49016 29656
rect 48688 29300 48740 29306
rect 48688 29242 48740 29248
rect 49068 28218 49096 31894
rect 49528 31822 49556 32166
rect 49516 31816 49568 31822
rect 49516 31758 49568 31764
rect 49712 31754 49740 33646
rect 50160 33652 50212 33658
rect 50160 33594 50212 33600
rect 50908 33646 51212 33674
rect 50908 33590 50936 33646
rect 51184 33590 51212 33646
rect 50896 33584 50948 33590
rect 50896 33526 50948 33532
rect 51172 33584 51224 33590
rect 51172 33526 51224 33532
rect 51276 33522 51304 33866
rect 49792 33516 49844 33522
rect 49792 33458 49844 33464
rect 51264 33516 51316 33522
rect 51264 33458 51316 33464
rect 49804 31822 49832 33458
rect 50804 33448 50856 33454
rect 50804 33390 50856 33396
rect 50436 33380 50488 33386
rect 50436 33322 50488 33328
rect 50448 32910 50476 33322
rect 50816 33046 50844 33390
rect 50896 33312 50948 33318
rect 50896 33254 50948 33260
rect 50988 33312 51040 33318
rect 50988 33254 51040 33260
rect 50804 33040 50856 33046
rect 50804 32982 50856 32988
rect 50436 32904 50488 32910
rect 50436 32846 50488 32852
rect 49884 32768 49936 32774
rect 49884 32710 49936 32716
rect 49896 32502 49924 32710
rect 50294 32668 50602 32677
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32603 50602 32612
rect 49884 32496 49936 32502
rect 49884 32438 49936 32444
rect 50908 31958 50936 33254
rect 51000 32910 51028 33254
rect 50988 32904 51040 32910
rect 50988 32846 51040 32852
rect 51264 32768 51316 32774
rect 51264 32710 51316 32716
rect 51080 32020 51132 32026
rect 51080 31962 51132 31968
rect 50896 31952 50948 31958
rect 50896 31894 50948 31900
rect 49792 31816 49844 31822
rect 49792 31758 49844 31764
rect 49620 31726 49740 31754
rect 49240 31680 49292 31686
rect 49240 31622 49292 31628
rect 49252 31482 49280 31622
rect 49240 31476 49292 31482
rect 49240 31418 49292 31424
rect 49516 31136 49568 31142
rect 49516 31078 49568 31084
rect 49240 29504 49292 29510
rect 49240 29446 49292 29452
rect 49424 29504 49476 29510
rect 49424 29446 49476 29452
rect 49252 29306 49280 29446
rect 49240 29300 49292 29306
rect 49240 29242 49292 29248
rect 49148 29164 49200 29170
rect 49148 29106 49200 29112
rect 49160 28762 49188 29106
rect 49436 28994 49464 29446
rect 49252 28966 49464 28994
rect 49148 28756 49200 28762
rect 49148 28698 49200 28704
rect 49160 28422 49188 28698
rect 49148 28416 49200 28422
rect 49148 28358 49200 28364
rect 49056 28212 49108 28218
rect 49056 28154 49108 28160
rect 49252 28082 49280 28966
rect 49240 28076 49292 28082
rect 49240 28018 49292 28024
rect 48320 27464 48372 27470
rect 48318 27432 48320 27441
rect 48596 27464 48648 27470
rect 48372 27432 48374 27441
rect 48596 27406 48648 27412
rect 49056 27464 49108 27470
rect 49056 27406 49108 27412
rect 48318 27367 48374 27376
rect 48148 27254 48268 27282
rect 48688 27328 48740 27334
rect 48688 27270 48740 27276
rect 48780 27328 48832 27334
rect 48780 27270 48832 27276
rect 48044 26376 48096 26382
rect 48148 26353 48176 27254
rect 48228 26988 48280 26994
rect 48228 26930 48280 26936
rect 48044 26318 48096 26324
rect 48134 26344 48190 26353
rect 48056 25906 48084 26318
rect 48134 26279 48190 26288
rect 47952 25900 48004 25906
rect 47952 25842 48004 25848
rect 48044 25900 48096 25906
rect 48044 25842 48096 25848
rect 47860 25764 47912 25770
rect 47860 25706 47912 25712
rect 47964 25498 47992 25842
rect 48148 25498 48176 26279
rect 48240 25974 48268 26930
rect 48504 26784 48556 26790
rect 48504 26726 48556 26732
rect 48516 26586 48544 26726
rect 48504 26580 48556 26586
rect 48504 26522 48556 26528
rect 48504 26444 48556 26450
rect 48504 26386 48556 26392
rect 48412 26308 48464 26314
rect 48412 26250 48464 26256
rect 48228 25968 48280 25974
rect 48228 25910 48280 25916
rect 48424 25906 48452 26250
rect 48412 25900 48464 25906
rect 48412 25842 48464 25848
rect 48424 25498 48452 25842
rect 47952 25492 48004 25498
rect 47952 25434 48004 25440
rect 48136 25492 48188 25498
rect 48136 25434 48188 25440
rect 48412 25492 48464 25498
rect 48412 25434 48464 25440
rect 48148 24274 48176 25434
rect 48424 24886 48452 25434
rect 48412 24880 48464 24886
rect 48412 24822 48464 24828
rect 48516 24818 48544 26386
rect 48596 25152 48648 25158
rect 48596 25094 48648 25100
rect 48228 24812 48280 24818
rect 48228 24754 48280 24760
rect 48504 24812 48556 24818
rect 48504 24754 48556 24760
rect 48240 24410 48268 24754
rect 48608 24750 48636 25094
rect 48596 24744 48648 24750
rect 48596 24686 48648 24692
rect 48412 24608 48464 24614
rect 48412 24550 48464 24556
rect 48228 24404 48280 24410
rect 48228 24346 48280 24352
rect 48136 24268 48188 24274
rect 48188 24228 48268 24256
rect 48136 24210 48188 24216
rect 48136 24064 48188 24070
rect 48136 24006 48188 24012
rect 47688 23854 47808 23882
rect 47308 23316 47360 23322
rect 47308 23258 47360 23264
rect 47216 22500 47268 22506
rect 47216 22442 47268 22448
rect 47124 22024 47176 22030
rect 47124 21966 47176 21972
rect 46664 21684 46716 21690
rect 46664 21626 46716 21632
rect 46204 21616 46256 21622
rect 46204 21558 46256 21564
rect 45652 21140 45704 21146
rect 45652 21082 45704 21088
rect 45468 21004 45520 21010
rect 45468 20946 45520 20952
rect 47032 20936 47084 20942
rect 47032 20878 47084 20884
rect 45744 20256 45796 20262
rect 45744 20198 45796 20204
rect 45756 19718 45784 20198
rect 47044 19922 47072 20878
rect 47124 20800 47176 20806
rect 47124 20742 47176 20748
rect 47032 19916 47084 19922
rect 47032 19858 47084 19864
rect 45744 19712 45796 19718
rect 45744 19654 45796 19660
rect 45652 18624 45704 18630
rect 45652 18566 45704 18572
rect 45664 18086 45692 18566
rect 45652 18080 45704 18086
rect 45652 18022 45704 18028
rect 44824 16040 44876 16046
rect 44824 15982 44876 15988
rect 45756 6914 45784 19654
rect 47044 18834 47072 19858
rect 47032 18828 47084 18834
rect 47032 18770 47084 18776
rect 46940 18692 46992 18698
rect 46940 18634 46992 18640
rect 46952 18426 46980 18634
rect 46940 18420 46992 18426
rect 46940 18362 46992 18368
rect 46940 16992 46992 16998
rect 46940 16934 46992 16940
rect 45928 16652 45980 16658
rect 45928 16594 45980 16600
rect 45940 16114 45968 16594
rect 46952 16590 46980 16934
rect 47044 16794 47072 18770
rect 47136 18306 47164 20742
rect 47216 19712 47268 19718
rect 47216 19654 47268 19660
rect 47228 19514 47256 19654
rect 47216 19508 47268 19514
rect 47216 19450 47268 19456
rect 47216 19236 47268 19242
rect 47216 19178 47268 19184
rect 47228 18426 47256 19178
rect 47400 19168 47452 19174
rect 47400 19110 47452 19116
rect 47412 18766 47440 19110
rect 47400 18760 47452 18766
rect 47400 18702 47452 18708
rect 47308 18624 47360 18630
rect 47308 18566 47360 18572
rect 47216 18420 47268 18426
rect 47216 18362 47268 18368
rect 47136 18278 47256 18306
rect 47320 18290 47348 18566
rect 47688 18426 47716 23854
rect 48044 23520 48096 23526
rect 48044 23462 48096 23468
rect 48056 23254 48084 23462
rect 48044 23248 48096 23254
rect 48044 23190 48096 23196
rect 47860 23112 47912 23118
rect 47860 23054 47912 23060
rect 47872 22778 47900 23054
rect 47952 22976 48004 22982
rect 47952 22918 48004 22924
rect 47964 22778 47992 22918
rect 48056 22778 48084 23190
rect 47860 22772 47912 22778
rect 47860 22714 47912 22720
rect 47952 22772 48004 22778
rect 47952 22714 48004 22720
rect 48044 22772 48096 22778
rect 48044 22714 48096 22720
rect 48044 22636 48096 22642
rect 48044 22578 48096 22584
rect 47952 22094 48004 22098
rect 48056 22094 48084 22578
rect 48148 22098 48176 24006
rect 48240 23254 48268 24228
rect 48424 24188 48452 24550
rect 48596 24200 48648 24206
rect 48424 24160 48596 24188
rect 48596 24142 48648 24148
rect 48596 23520 48648 23526
rect 48596 23462 48648 23468
rect 48608 23322 48636 23462
rect 48596 23316 48648 23322
rect 48596 23258 48648 23264
rect 48228 23248 48280 23254
rect 48228 23190 48280 23196
rect 47952 22092 48084 22094
rect 48004 22052 48084 22092
rect 47952 22034 48004 22040
rect 47768 21344 47820 21350
rect 47768 21286 47820 21292
rect 47780 21146 47808 21286
rect 47768 21140 47820 21146
rect 47768 21082 47820 21088
rect 47952 21004 48004 21010
rect 47952 20946 48004 20952
rect 47964 19514 47992 20946
rect 47952 19508 48004 19514
rect 47952 19450 48004 19456
rect 47676 18420 47728 18426
rect 47676 18362 47728 18368
rect 47124 16992 47176 16998
rect 47124 16934 47176 16940
rect 47032 16788 47084 16794
rect 47032 16730 47084 16736
rect 46940 16584 46992 16590
rect 46940 16526 46992 16532
rect 45928 16108 45980 16114
rect 45928 16050 45980 16056
rect 45940 15570 45968 16050
rect 45928 15564 45980 15570
rect 45928 15506 45980 15512
rect 45940 13394 45968 15506
rect 46572 15428 46624 15434
rect 46572 15370 46624 15376
rect 46584 15162 46612 15370
rect 46572 15156 46624 15162
rect 46572 15098 46624 15104
rect 47136 14890 47164 16934
rect 47124 14884 47176 14890
rect 47124 14826 47176 14832
rect 47136 14056 47164 14826
rect 47044 14028 47164 14056
rect 45928 13388 45980 13394
rect 45928 13330 45980 13336
rect 46296 13388 46348 13394
rect 46296 13330 46348 13336
rect 46308 12434 46336 13330
rect 46848 13252 46900 13258
rect 46848 13194 46900 13200
rect 46860 12986 46888 13194
rect 46848 12980 46900 12986
rect 46848 12922 46900 12928
rect 47044 12850 47072 14028
rect 47124 13932 47176 13938
rect 47124 13874 47176 13880
rect 47136 12850 47164 13874
rect 47032 12844 47084 12850
rect 47032 12786 47084 12792
rect 47124 12844 47176 12850
rect 47124 12786 47176 12792
rect 46308 12406 46428 12434
rect 46400 12306 46428 12406
rect 46388 12300 46440 12306
rect 46388 12242 46440 12248
rect 45664 6886 45784 6914
rect 42616 2644 42668 2650
rect 42616 2586 42668 2592
rect 45664 2514 45692 6886
rect 45652 2508 45704 2514
rect 45652 2450 45704 2456
rect 47228 2446 47256 18278
rect 47308 18284 47360 18290
rect 47308 18226 47360 18232
rect 47860 17672 47912 17678
rect 47860 17614 47912 17620
rect 47308 17536 47360 17542
rect 47308 17478 47360 17484
rect 47320 17338 47348 17478
rect 47872 17338 47900 17614
rect 47308 17332 47360 17338
rect 47308 17274 47360 17280
rect 47860 17332 47912 17338
rect 47860 17274 47912 17280
rect 48056 17270 48084 22052
rect 48136 22092 48188 22098
rect 48700 22094 48728 27270
rect 48792 26994 48820 27270
rect 48780 26988 48832 26994
rect 48780 26930 48832 26936
rect 48792 26790 48820 26930
rect 48780 26784 48832 26790
rect 48780 26726 48832 26732
rect 48792 26042 48820 26726
rect 48780 26036 48832 26042
rect 48780 25978 48832 25984
rect 48872 25288 48924 25294
rect 48872 25230 48924 25236
rect 48780 24948 48832 24954
rect 48780 24890 48832 24896
rect 48792 24274 48820 24890
rect 48884 24410 48912 25230
rect 48964 24744 49016 24750
rect 48964 24686 49016 24692
rect 48976 24410 49004 24686
rect 48872 24404 48924 24410
rect 48872 24346 48924 24352
rect 48964 24404 49016 24410
rect 48964 24346 49016 24352
rect 48780 24268 48832 24274
rect 48780 24210 48832 24216
rect 48964 24200 49016 24206
rect 48964 24142 49016 24148
rect 48976 23730 49004 24142
rect 48964 23724 49016 23730
rect 48964 23666 49016 23672
rect 48976 23254 49004 23666
rect 48964 23248 49016 23254
rect 48964 23190 49016 23196
rect 48872 22432 48924 22438
rect 48872 22374 48924 22380
rect 48136 22034 48188 22040
rect 48608 22066 48728 22094
rect 48320 20936 48372 20942
rect 48320 20878 48372 20884
rect 48228 20596 48280 20602
rect 48332 20584 48360 20878
rect 48412 20868 48464 20874
rect 48412 20810 48464 20816
rect 48280 20556 48360 20584
rect 48228 20538 48280 20544
rect 48424 20534 48452 20810
rect 48504 20800 48556 20806
rect 48504 20742 48556 20748
rect 48516 20602 48544 20742
rect 48504 20596 48556 20602
rect 48504 20538 48556 20544
rect 48412 20528 48464 20534
rect 48412 20470 48464 20476
rect 48608 20466 48636 22066
rect 48688 21956 48740 21962
rect 48688 21898 48740 21904
rect 48504 20460 48556 20466
rect 48504 20402 48556 20408
rect 48596 20460 48648 20466
rect 48596 20402 48648 20408
rect 48320 20256 48372 20262
rect 48320 20198 48372 20204
rect 48332 20058 48360 20198
rect 48516 20058 48544 20402
rect 48320 20052 48372 20058
rect 48320 19994 48372 20000
rect 48504 20052 48556 20058
rect 48504 19994 48556 20000
rect 48596 19848 48648 19854
rect 48596 19790 48648 19796
rect 48412 19712 48464 19718
rect 48412 19654 48464 19660
rect 48320 19168 48372 19174
rect 48320 19110 48372 19116
rect 48332 18766 48360 19110
rect 48424 18766 48452 19654
rect 48320 18760 48372 18766
rect 48320 18702 48372 18708
rect 48412 18760 48464 18766
rect 48412 18702 48464 18708
rect 48608 18426 48636 19790
rect 48596 18420 48648 18426
rect 48596 18362 48648 18368
rect 48320 17876 48372 17882
rect 48320 17818 48372 17824
rect 48044 17264 48096 17270
rect 48096 17212 48176 17218
rect 48044 17206 48176 17212
rect 48056 17190 48176 17206
rect 47676 17128 47728 17134
rect 47676 17070 47728 17076
rect 48044 17128 48096 17134
rect 48044 17070 48096 17076
rect 47688 16590 47716 17070
rect 48056 16794 48084 17070
rect 48044 16788 48096 16794
rect 48044 16730 48096 16736
rect 47676 16584 47728 16590
rect 47676 16526 47728 16532
rect 47688 16114 47716 16526
rect 47676 16108 47728 16114
rect 47676 16050 47728 16056
rect 48044 16108 48096 16114
rect 48044 16050 48096 16056
rect 47492 15360 47544 15366
rect 47492 15302 47544 15308
rect 47584 15360 47636 15366
rect 47584 15302 47636 15308
rect 47504 14958 47532 15302
rect 47596 15026 47624 15302
rect 47584 15020 47636 15026
rect 47584 14962 47636 14968
rect 47492 14952 47544 14958
rect 47492 14894 47544 14900
rect 47584 13932 47636 13938
rect 47584 13874 47636 13880
rect 47596 13530 47624 13874
rect 47584 13524 47636 13530
rect 47584 13466 47636 13472
rect 47688 12850 47716 16050
rect 47952 15904 48004 15910
rect 47952 15846 48004 15852
rect 47964 15706 47992 15846
rect 47952 15700 48004 15706
rect 47952 15642 48004 15648
rect 48056 15366 48084 16050
rect 48044 15360 48096 15366
rect 48044 15302 48096 15308
rect 48148 15026 48176 17190
rect 48332 16182 48360 17818
rect 48700 17338 48728 21898
rect 48780 21480 48832 21486
rect 48780 21422 48832 21428
rect 48792 20602 48820 21422
rect 48780 20596 48832 20602
rect 48780 20538 48832 20544
rect 48884 18290 48912 22374
rect 49068 21078 49096 27406
rect 49252 27334 49280 28018
rect 49424 28008 49476 28014
rect 49424 27950 49476 27956
rect 49240 27328 49292 27334
rect 49240 27270 49292 27276
rect 49148 25764 49200 25770
rect 49148 25706 49200 25712
rect 49160 25158 49188 25706
rect 49436 25702 49464 27950
rect 49424 25696 49476 25702
rect 49424 25638 49476 25644
rect 49424 25424 49476 25430
rect 49424 25366 49476 25372
rect 49148 25152 49200 25158
rect 49148 25094 49200 25100
rect 49160 21962 49188 25094
rect 49240 24880 49292 24886
rect 49240 24822 49292 24828
rect 49252 22710 49280 24822
rect 49332 23520 49384 23526
rect 49332 23462 49384 23468
rect 49240 22704 49292 22710
rect 49240 22646 49292 22652
rect 49344 22030 49372 23462
rect 49332 22024 49384 22030
rect 49332 21966 49384 21972
rect 49148 21956 49200 21962
rect 49148 21898 49200 21904
rect 49240 21888 49292 21894
rect 49240 21830 49292 21836
rect 49056 21072 49108 21078
rect 49056 21014 49108 21020
rect 49068 20398 49096 21014
rect 49148 20596 49200 20602
rect 49148 20538 49200 20544
rect 49056 20392 49108 20398
rect 49056 20334 49108 20340
rect 49160 19514 49188 20538
rect 49148 19508 49200 19514
rect 49148 19450 49200 19456
rect 49056 19304 49108 19310
rect 49056 19246 49108 19252
rect 48872 18284 48924 18290
rect 48872 18226 48924 18232
rect 48688 17332 48740 17338
rect 48688 17274 48740 17280
rect 48700 16794 48728 17274
rect 48780 17196 48832 17202
rect 48780 17138 48832 17144
rect 48792 17066 48820 17138
rect 48780 17060 48832 17066
rect 48780 17002 48832 17008
rect 48688 16788 48740 16794
rect 48688 16730 48740 16736
rect 48320 16176 48372 16182
rect 48320 16118 48372 16124
rect 48700 16114 48728 16730
rect 48412 16108 48464 16114
rect 48412 16050 48464 16056
rect 48688 16108 48740 16114
rect 48688 16050 48740 16056
rect 48320 15972 48372 15978
rect 48320 15914 48372 15920
rect 47952 15020 48004 15026
rect 47952 14962 48004 14968
rect 48136 15020 48188 15026
rect 48136 14962 48188 14968
rect 47964 13938 47992 14962
rect 48332 14074 48360 15914
rect 48424 15162 48452 16050
rect 48504 16040 48556 16046
rect 48504 15982 48556 15988
rect 48516 15434 48544 15982
rect 48504 15428 48556 15434
rect 48504 15370 48556 15376
rect 48412 15156 48464 15162
rect 48412 15098 48464 15104
rect 48516 15026 48544 15370
rect 49068 15162 49096 19246
rect 49148 18624 49200 18630
rect 49148 18566 49200 18572
rect 49160 18426 49188 18566
rect 49148 18420 49200 18426
rect 49148 18362 49200 18368
rect 49252 17678 49280 21830
rect 49436 21690 49464 25366
rect 49424 21684 49476 21690
rect 49344 21644 49424 21672
rect 49344 20602 49372 21644
rect 49424 21626 49476 21632
rect 49528 21554 49556 31078
rect 49620 30394 49648 31726
rect 50294 31580 50602 31589
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31515 50602 31524
rect 51092 31346 51120 31962
rect 51080 31340 51132 31346
rect 51080 31282 51132 31288
rect 51172 30660 51224 30666
rect 51172 30602 51224 30608
rect 50160 30592 50212 30598
rect 50160 30534 50212 30540
rect 49608 30388 49660 30394
rect 49608 30330 49660 30336
rect 50172 30326 50200 30534
rect 50294 30492 50602 30501
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30427 50602 30436
rect 50160 30320 50212 30326
rect 50160 30262 50212 30268
rect 50160 29776 50212 29782
rect 50160 29718 50212 29724
rect 49976 29640 50028 29646
rect 49976 29582 50028 29588
rect 49792 29028 49844 29034
rect 49792 28970 49844 28976
rect 49700 28484 49752 28490
rect 49700 28426 49752 28432
rect 49712 28218 49740 28426
rect 49700 28212 49752 28218
rect 49700 28154 49752 28160
rect 49700 27396 49752 27402
rect 49700 27338 49752 27344
rect 49606 27160 49662 27169
rect 49606 27095 49662 27104
rect 49620 23254 49648 27095
rect 49712 26994 49740 27338
rect 49700 26988 49752 26994
rect 49700 26930 49752 26936
rect 49804 26314 49832 28970
rect 49884 28688 49936 28694
rect 49884 28630 49936 28636
rect 49792 26308 49844 26314
rect 49792 26250 49844 26256
rect 49804 25702 49832 26250
rect 49792 25696 49844 25702
rect 49790 25664 49792 25673
rect 49844 25664 49846 25673
rect 49790 25599 49846 25608
rect 49792 23860 49844 23866
rect 49792 23802 49844 23808
rect 49804 23662 49832 23802
rect 49792 23656 49844 23662
rect 49792 23598 49844 23604
rect 49608 23248 49660 23254
rect 49608 23190 49660 23196
rect 49804 22778 49832 23598
rect 49792 22772 49844 22778
rect 49792 22714 49844 22720
rect 49896 21554 49924 28630
rect 49988 28422 50016 29582
rect 50172 28762 50200 29718
rect 50620 29708 50672 29714
rect 50620 29650 50672 29656
rect 50294 29404 50602 29413
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29339 50602 29348
rect 50160 28756 50212 28762
rect 50160 28698 50212 28704
rect 50252 28620 50304 28626
rect 50252 28562 50304 28568
rect 49976 28416 50028 28422
rect 49976 28358 50028 28364
rect 50068 28416 50120 28422
rect 50264 28404 50292 28562
rect 50632 28558 50660 29650
rect 51080 29640 51132 29646
rect 51080 29582 51132 29588
rect 50710 28656 50766 28665
rect 51092 28608 51120 29582
rect 50710 28591 50766 28600
rect 50620 28552 50672 28558
rect 50620 28494 50672 28500
rect 50724 28490 50752 28591
rect 51000 28580 51120 28608
rect 50712 28484 50764 28490
rect 50712 28426 50764 28432
rect 50068 28358 50120 28364
rect 50172 28376 50292 28404
rect 49988 27878 50016 28358
rect 49976 27872 50028 27878
rect 49976 27814 50028 27820
rect 50080 27713 50108 28358
rect 50172 28218 50200 28376
rect 50294 28316 50602 28325
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28251 50602 28260
rect 50160 28212 50212 28218
rect 50160 28154 50212 28160
rect 50158 28112 50214 28121
rect 50158 28047 50160 28056
rect 50212 28047 50214 28056
rect 50160 28018 50212 28024
rect 50066 27704 50122 27713
rect 50066 27639 50122 27648
rect 50620 27600 50672 27606
rect 50618 27568 50620 27577
rect 50672 27568 50674 27577
rect 50618 27503 50674 27512
rect 51000 27470 51028 28580
rect 51184 28082 51212 30602
rect 51172 28076 51224 28082
rect 51172 28018 51224 28024
rect 49976 27464 50028 27470
rect 49976 27406 50028 27412
rect 50988 27464 51040 27470
rect 50988 27406 51040 27412
rect 49988 27062 50016 27406
rect 50896 27328 50948 27334
rect 50896 27270 50948 27276
rect 50294 27228 50602 27237
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27163 50602 27172
rect 49976 27056 50028 27062
rect 49976 26998 50028 27004
rect 50908 26994 50936 27270
rect 50896 26988 50948 26994
rect 50896 26930 50948 26936
rect 50160 26920 50212 26926
rect 50160 26862 50212 26868
rect 50172 26586 50200 26862
rect 50804 26784 50856 26790
rect 50804 26726 50856 26732
rect 50160 26580 50212 26586
rect 50160 26522 50212 26528
rect 50294 26140 50602 26149
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26075 50602 26084
rect 50816 25974 50844 26726
rect 51080 26512 51132 26518
rect 51080 26454 51132 26460
rect 50804 25968 50856 25974
rect 50804 25910 50856 25916
rect 51092 25906 51120 26454
rect 51276 26042 51304 32710
rect 51460 31822 51488 34478
rect 52184 34400 52236 34406
rect 52184 34342 52236 34348
rect 51540 33856 51592 33862
rect 51540 33798 51592 33804
rect 51552 33522 51580 33798
rect 52196 33522 52224 34342
rect 52644 34196 52696 34202
rect 52644 34138 52696 34144
rect 52656 33658 52684 34138
rect 52644 33652 52696 33658
rect 52644 33594 52696 33600
rect 51540 33516 51592 33522
rect 51540 33458 51592 33464
rect 52184 33516 52236 33522
rect 52184 33458 52236 33464
rect 51552 32774 51580 33458
rect 52656 33318 52684 33594
rect 52644 33312 52696 33318
rect 52644 33254 52696 33260
rect 51540 32768 51592 32774
rect 51540 32710 51592 32716
rect 52552 31952 52604 31958
rect 52552 31894 52604 31900
rect 52460 31884 52512 31890
rect 52460 31826 52512 31832
rect 51448 31816 51500 31822
rect 51448 31758 51500 31764
rect 52092 31816 52144 31822
rect 52092 31758 52144 31764
rect 51816 31272 51868 31278
rect 51816 31214 51868 31220
rect 51356 31136 51408 31142
rect 51356 31078 51408 31084
rect 51724 31136 51776 31142
rect 51724 31078 51776 31084
rect 51368 29578 51396 31078
rect 51736 30802 51764 31078
rect 51828 30938 51856 31214
rect 51816 30932 51868 30938
rect 51816 30874 51868 30880
rect 51724 30796 51776 30802
rect 51724 30738 51776 30744
rect 51632 30592 51684 30598
rect 51632 30534 51684 30540
rect 51644 30258 51672 30534
rect 51736 30394 51764 30738
rect 51816 30660 51868 30666
rect 51816 30602 51868 30608
rect 51724 30388 51776 30394
rect 51724 30330 51776 30336
rect 51632 30252 51684 30258
rect 51632 30194 51684 30200
rect 51448 29640 51500 29646
rect 51448 29582 51500 29588
rect 51356 29572 51408 29578
rect 51356 29514 51408 29520
rect 51356 29232 51408 29238
rect 51354 29200 51356 29209
rect 51460 29220 51488 29582
rect 51540 29572 51592 29578
rect 51540 29514 51592 29520
rect 51552 29481 51580 29514
rect 51538 29472 51594 29481
rect 51538 29407 51594 29416
rect 51408 29200 51488 29220
rect 51410 29192 51488 29200
rect 51354 29135 51410 29144
rect 51540 29164 51592 29170
rect 51540 29106 51592 29112
rect 51552 28762 51580 29106
rect 51540 28756 51592 28762
rect 51540 28698 51592 28704
rect 51540 28416 51592 28422
rect 51644 28404 51672 30194
rect 51828 30190 51856 30602
rect 52104 30258 52132 31758
rect 52472 31482 52500 31826
rect 52460 31476 52512 31482
rect 52460 31418 52512 31424
rect 52564 31142 52592 31894
rect 52552 31136 52604 31142
rect 52552 31078 52604 31084
rect 52092 30252 52144 30258
rect 52092 30194 52144 30200
rect 51816 30184 51868 30190
rect 51816 30126 51868 30132
rect 51828 29850 51856 30126
rect 52104 30122 52132 30194
rect 52092 30116 52144 30122
rect 52092 30058 52144 30064
rect 51908 30048 51960 30054
rect 51908 29990 51960 29996
rect 52000 30048 52052 30054
rect 52184 30048 52236 30054
rect 52052 29996 52132 30002
rect 52000 29990 52132 29996
rect 52184 29990 52236 29996
rect 51816 29844 51868 29850
rect 51816 29786 51868 29792
rect 51828 29646 51856 29786
rect 51816 29640 51868 29646
rect 51736 29600 51816 29628
rect 51736 28558 51764 29600
rect 51816 29582 51868 29588
rect 51816 29164 51868 29170
rect 51816 29106 51868 29112
rect 51828 28762 51856 29106
rect 51816 28756 51868 28762
rect 51816 28698 51868 28704
rect 51724 28552 51776 28558
rect 51776 28512 51856 28540
rect 51724 28494 51776 28500
rect 51592 28376 51672 28404
rect 51724 28416 51776 28422
rect 51540 28358 51592 28364
rect 51724 28358 51776 28364
rect 51448 27396 51500 27402
rect 51448 27338 51500 27344
rect 51460 27130 51488 27338
rect 51552 27130 51580 28358
rect 51632 27872 51684 27878
rect 51632 27814 51684 27820
rect 51448 27124 51500 27130
rect 51448 27066 51500 27072
rect 51540 27124 51592 27130
rect 51540 27066 51592 27072
rect 51644 26926 51672 27814
rect 51632 26920 51684 26926
rect 51632 26862 51684 26868
rect 51736 26858 51764 28358
rect 51724 26852 51776 26858
rect 51724 26794 51776 26800
rect 51632 26784 51684 26790
rect 51632 26726 51684 26732
rect 51264 26036 51316 26042
rect 51264 25978 51316 25984
rect 51080 25900 51132 25906
rect 51080 25842 51132 25848
rect 51356 25900 51408 25906
rect 51356 25842 51408 25848
rect 50160 25832 50212 25838
rect 50160 25774 50212 25780
rect 50068 23656 50120 23662
rect 50068 23598 50120 23604
rect 49976 23316 50028 23322
rect 49976 23258 50028 23264
rect 49988 22094 50016 23258
rect 50080 23186 50108 23598
rect 50068 23180 50120 23186
rect 50068 23122 50120 23128
rect 50172 22098 50200 25774
rect 51368 25498 51396 25842
rect 51644 25498 51672 26726
rect 51828 26382 51856 28512
rect 51920 28150 51948 29990
rect 52012 29974 52132 29990
rect 52104 29850 52132 29974
rect 52092 29844 52144 29850
rect 52092 29786 52144 29792
rect 52000 29776 52052 29782
rect 52000 29718 52052 29724
rect 52012 29102 52040 29718
rect 52000 29096 52052 29102
rect 52000 29038 52052 29044
rect 52104 28994 52132 29786
rect 52196 29646 52224 29990
rect 52184 29640 52236 29646
rect 52184 29582 52236 29588
rect 52460 29640 52512 29646
rect 52460 29582 52512 29588
rect 52276 29504 52328 29510
rect 52276 29446 52328 29452
rect 52012 28966 52132 28994
rect 52012 28558 52040 28966
rect 52000 28552 52052 28558
rect 52000 28494 52052 28500
rect 52184 28552 52236 28558
rect 52184 28494 52236 28500
rect 51908 28144 51960 28150
rect 51908 28086 51960 28092
rect 51920 27470 51948 28086
rect 51908 27464 51960 27470
rect 51908 27406 51960 27412
rect 51920 26586 51948 27406
rect 52196 27062 52224 28494
rect 52184 27056 52236 27062
rect 52184 26998 52236 27004
rect 51908 26580 51960 26586
rect 51908 26522 51960 26528
rect 51816 26376 51868 26382
rect 51816 26318 51868 26324
rect 51356 25492 51408 25498
rect 51356 25434 51408 25440
rect 51632 25492 51684 25498
rect 51632 25434 51684 25440
rect 50294 25052 50602 25061
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24987 50602 24996
rect 51632 24812 51684 24818
rect 51632 24754 51684 24760
rect 51816 24812 51868 24818
rect 51816 24754 51868 24760
rect 52092 24812 52144 24818
rect 52092 24754 52144 24760
rect 51080 24608 51132 24614
rect 51080 24550 51132 24556
rect 51448 24608 51500 24614
rect 51448 24550 51500 24556
rect 50620 24200 50672 24206
rect 50620 24142 50672 24148
rect 50632 24070 50660 24142
rect 51092 24138 51120 24550
rect 51460 24206 51488 24550
rect 51644 24342 51672 24754
rect 51724 24608 51776 24614
rect 51724 24550 51776 24556
rect 51736 24410 51764 24550
rect 51828 24410 51856 24754
rect 52104 24410 52132 24754
rect 51724 24404 51776 24410
rect 51724 24346 51776 24352
rect 51816 24404 51868 24410
rect 51816 24346 51868 24352
rect 52092 24404 52144 24410
rect 52092 24346 52144 24352
rect 51632 24336 51684 24342
rect 51632 24278 51684 24284
rect 52288 24206 52316 29446
rect 52472 29306 52500 29582
rect 52460 29300 52512 29306
rect 52460 29242 52512 29248
rect 52552 29300 52604 29306
rect 52552 29242 52604 29248
rect 52564 29034 52592 29242
rect 52656 29170 52684 33254
rect 52736 32768 52788 32774
rect 52736 32710 52788 32716
rect 52748 32570 52776 32710
rect 52736 32564 52788 32570
rect 52736 32506 52788 32512
rect 55128 32564 55180 32570
rect 55128 32506 55180 32512
rect 53748 32496 53800 32502
rect 53748 32438 53800 32444
rect 53196 32428 53248 32434
rect 53196 32370 53248 32376
rect 53104 32224 53156 32230
rect 53104 32166 53156 32172
rect 53012 31748 53064 31754
rect 53012 31690 53064 31696
rect 53024 31482 53052 31690
rect 53012 31476 53064 31482
rect 53012 31418 53064 31424
rect 52920 31408 52972 31414
rect 52920 31350 52972 31356
rect 52932 30258 52960 31350
rect 53116 31278 53144 32166
rect 53104 31272 53156 31278
rect 53104 31214 53156 31220
rect 53208 31124 53236 32370
rect 53760 31414 53788 32438
rect 54392 32360 54444 32366
rect 54392 32302 54444 32308
rect 54404 32026 54432 32302
rect 55036 32224 55088 32230
rect 55036 32166 55088 32172
rect 54392 32020 54444 32026
rect 54392 31962 54444 31968
rect 55048 31754 55076 32166
rect 55140 31822 55168 32506
rect 55128 31816 55180 31822
rect 55128 31758 55180 31764
rect 54956 31726 55076 31754
rect 54852 31680 54904 31686
rect 54852 31622 54904 31628
rect 54864 31414 54892 31622
rect 53748 31408 53800 31414
rect 53748 31350 53800 31356
rect 54852 31408 54904 31414
rect 54852 31350 54904 31356
rect 54956 31278 54984 31726
rect 55140 31346 55168 31758
rect 55220 31748 55272 31754
rect 55220 31690 55272 31696
rect 55232 31482 55260 31690
rect 55220 31476 55272 31482
rect 55220 31418 55272 31424
rect 55128 31340 55180 31346
rect 55128 31282 55180 31288
rect 54944 31272 54996 31278
rect 54944 31214 54996 31220
rect 54852 31204 54904 31210
rect 54852 31146 54904 31152
rect 53116 31096 53236 31124
rect 54484 31136 54536 31142
rect 53116 30734 53144 31096
rect 54484 31078 54536 31084
rect 54496 30938 54524 31078
rect 54484 30932 54536 30938
rect 54484 30874 54536 30880
rect 53104 30728 53156 30734
rect 53104 30670 53156 30676
rect 53472 30592 53524 30598
rect 53472 30534 53524 30540
rect 54300 30592 54352 30598
rect 54300 30534 54352 30540
rect 53484 30394 53512 30534
rect 53472 30388 53524 30394
rect 53472 30330 53524 30336
rect 53564 30320 53616 30326
rect 53208 30268 53564 30274
rect 53208 30262 53616 30268
rect 53208 30258 53604 30262
rect 54312 30258 54340 30534
rect 54864 30326 54892 31146
rect 54852 30320 54904 30326
rect 54852 30262 54904 30268
rect 52920 30252 52972 30258
rect 52920 30194 52972 30200
rect 53196 30252 53604 30258
rect 53248 30246 53604 30252
rect 54300 30252 54352 30258
rect 53196 30194 53248 30200
rect 54300 30194 54352 30200
rect 54668 30252 54720 30258
rect 54668 30194 54720 30200
rect 53208 29850 53236 30194
rect 54576 30184 54628 30190
rect 54576 30126 54628 30132
rect 53380 30048 53432 30054
rect 53380 29990 53432 29996
rect 54392 30048 54444 30054
rect 54392 29990 54444 29996
rect 53392 29850 53420 29990
rect 53196 29844 53248 29850
rect 53196 29786 53248 29792
rect 53380 29844 53432 29850
rect 53380 29786 53432 29792
rect 54404 29714 54432 29990
rect 54392 29708 54444 29714
rect 54392 29650 54444 29656
rect 53564 29640 53616 29646
rect 53484 29600 53564 29628
rect 53012 29504 53064 29510
rect 52918 29472 52974 29481
rect 53012 29446 53064 29452
rect 52918 29407 52974 29416
rect 52644 29164 52696 29170
rect 52644 29106 52696 29112
rect 52552 29028 52604 29034
rect 52552 28970 52604 28976
rect 52932 28994 52960 29407
rect 53024 29306 53052 29446
rect 53012 29300 53064 29306
rect 53012 29242 53064 29248
rect 53484 29170 53512 29600
rect 53564 29582 53616 29588
rect 53840 29572 53892 29578
rect 53840 29514 53892 29520
rect 53564 29504 53616 29510
rect 53564 29446 53616 29452
rect 53104 29164 53156 29170
rect 53104 29106 53156 29112
rect 53472 29164 53524 29170
rect 53472 29106 53524 29112
rect 52932 28966 53052 28994
rect 52552 28552 52604 28558
rect 52552 28494 52604 28500
rect 52564 28082 52592 28494
rect 52368 28076 52420 28082
rect 52368 28018 52420 28024
rect 52552 28076 52604 28082
rect 52552 28018 52604 28024
rect 52380 27656 52408 28018
rect 52920 28008 52972 28014
rect 52920 27950 52972 27956
rect 52932 27674 52960 27950
rect 52920 27668 52972 27674
rect 52380 27628 52500 27656
rect 52472 25906 52500 27628
rect 52920 27610 52972 27616
rect 53024 27334 53052 28966
rect 53012 27328 53064 27334
rect 53012 27270 53064 27276
rect 52736 26376 52788 26382
rect 52736 26318 52788 26324
rect 52748 26042 52776 26318
rect 52828 26308 52880 26314
rect 52828 26250 52880 26256
rect 52736 26036 52788 26042
rect 52736 25978 52788 25984
rect 52460 25900 52512 25906
rect 52460 25842 52512 25848
rect 52736 25696 52788 25702
rect 52736 25638 52788 25644
rect 52748 25498 52776 25638
rect 52736 25492 52788 25498
rect 52736 25434 52788 25440
rect 52460 24880 52512 24886
rect 52460 24822 52512 24828
rect 52368 24608 52420 24614
rect 52368 24550 52420 24556
rect 51448 24200 51500 24206
rect 51448 24142 51500 24148
rect 52276 24200 52328 24206
rect 52276 24142 52328 24148
rect 51080 24132 51132 24138
rect 51080 24074 51132 24080
rect 50620 24064 50672 24070
rect 50620 24006 50672 24012
rect 50712 24064 50764 24070
rect 50712 24006 50764 24012
rect 51356 24064 51408 24070
rect 51356 24006 51408 24012
rect 51908 24064 51960 24070
rect 51908 24006 51960 24012
rect 50294 23964 50602 23973
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23899 50602 23908
rect 50632 23866 50660 24006
rect 50528 23860 50580 23866
rect 50528 23802 50580 23808
rect 50620 23860 50672 23866
rect 50620 23802 50672 23808
rect 50540 23730 50568 23802
rect 50528 23724 50580 23730
rect 50528 23666 50580 23672
rect 50344 23588 50396 23594
rect 50344 23530 50396 23536
rect 50356 23118 50384 23530
rect 50344 23112 50396 23118
rect 50344 23054 50396 23060
rect 50540 23050 50568 23666
rect 50724 23594 50752 24006
rect 50712 23588 50764 23594
rect 50712 23530 50764 23536
rect 50620 23520 50672 23526
rect 50620 23462 50672 23468
rect 50528 23044 50580 23050
rect 50528 22986 50580 22992
rect 50294 22876 50602 22885
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22811 50602 22820
rect 49988 22066 50108 22094
rect 49424 21548 49476 21554
rect 49424 21490 49476 21496
rect 49516 21548 49568 21554
rect 49516 21490 49568 21496
rect 49884 21548 49936 21554
rect 49884 21490 49936 21496
rect 49436 21146 49464 21490
rect 49608 21412 49660 21418
rect 49608 21354 49660 21360
rect 49620 21146 49648 21354
rect 49700 21344 49752 21350
rect 49700 21286 49752 21292
rect 49712 21146 49740 21286
rect 49424 21140 49476 21146
rect 49424 21082 49476 21088
rect 49608 21140 49660 21146
rect 49608 21082 49660 21088
rect 49700 21140 49752 21146
rect 49700 21082 49752 21088
rect 50080 21010 50108 22066
rect 50160 22092 50212 22098
rect 50160 22034 50212 22040
rect 50294 21788 50602 21797
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21723 50602 21732
rect 50160 21548 50212 21554
rect 50160 21490 50212 21496
rect 50528 21548 50580 21554
rect 50528 21490 50580 21496
rect 50068 21004 50120 21010
rect 50068 20946 50120 20952
rect 49976 20936 50028 20942
rect 49976 20878 50028 20884
rect 49332 20596 49384 20602
rect 49332 20538 49384 20544
rect 49700 20596 49752 20602
rect 49700 20538 49752 20544
rect 49424 20392 49476 20398
rect 49424 20334 49476 20340
rect 49436 19922 49464 20334
rect 49424 19916 49476 19922
rect 49424 19858 49476 19864
rect 49608 19848 49660 19854
rect 49344 19796 49608 19802
rect 49344 19790 49660 19796
rect 49344 19774 49648 19790
rect 49344 19514 49372 19774
rect 49516 19712 49568 19718
rect 49516 19654 49568 19660
rect 49332 19508 49384 19514
rect 49332 19450 49384 19456
rect 49528 19334 49556 19654
rect 49712 19378 49740 20538
rect 49792 19848 49844 19854
rect 49792 19790 49844 19796
rect 49436 19306 49556 19334
rect 49700 19372 49752 19378
rect 49700 19314 49752 19320
rect 49804 19310 49832 19790
rect 49884 19372 49936 19378
rect 49884 19314 49936 19320
rect 49436 18834 49464 19306
rect 49792 19304 49844 19310
rect 49792 19246 49844 19252
rect 49896 18970 49924 19314
rect 49884 18964 49936 18970
rect 49884 18906 49936 18912
rect 49424 18828 49476 18834
rect 49424 18770 49476 18776
rect 49516 18828 49568 18834
rect 49516 18770 49568 18776
rect 49332 18692 49384 18698
rect 49332 18634 49384 18640
rect 49344 18426 49372 18634
rect 49332 18420 49384 18426
rect 49332 18362 49384 18368
rect 49240 17672 49292 17678
rect 49240 17614 49292 17620
rect 49148 17536 49200 17542
rect 49148 17478 49200 17484
rect 49240 17536 49292 17542
rect 49240 17478 49292 17484
rect 49056 15156 49108 15162
rect 49056 15098 49108 15104
rect 48504 15020 48556 15026
rect 48504 14962 48556 14968
rect 48688 15020 48740 15026
rect 48688 14962 48740 14968
rect 48780 15020 48832 15026
rect 48780 14962 48832 14968
rect 48516 14618 48544 14962
rect 48700 14618 48728 14962
rect 48504 14612 48556 14618
rect 48504 14554 48556 14560
rect 48688 14612 48740 14618
rect 48688 14554 48740 14560
rect 48504 14272 48556 14278
rect 48504 14214 48556 14220
rect 48320 14068 48372 14074
rect 48320 14010 48372 14016
rect 47952 13932 48004 13938
rect 47952 13874 48004 13880
rect 48516 13870 48544 14214
rect 48504 13864 48556 13870
rect 48504 13806 48556 13812
rect 47952 13524 48004 13530
rect 47952 13466 48004 13472
rect 47768 13184 47820 13190
rect 47768 13126 47820 13132
rect 47780 12986 47808 13126
rect 47768 12980 47820 12986
rect 47768 12922 47820 12928
rect 47964 12850 47992 13466
rect 48320 13320 48372 13326
rect 48320 13262 48372 13268
rect 48332 12986 48360 13262
rect 48320 12980 48372 12986
rect 48320 12922 48372 12928
rect 47676 12844 47728 12850
rect 47676 12786 47728 12792
rect 47952 12844 48004 12850
rect 47952 12786 48004 12792
rect 48504 12640 48556 12646
rect 48504 12582 48556 12588
rect 48516 12238 48544 12582
rect 48504 12232 48556 12238
rect 48504 12174 48556 12180
rect 48792 10810 48820 14962
rect 49160 14618 49188 17478
rect 49252 17338 49280 17478
rect 49240 17332 49292 17338
rect 49240 17274 49292 17280
rect 49332 17196 49384 17202
rect 49332 17138 49384 17144
rect 49344 17082 49372 17138
rect 49252 17054 49372 17082
rect 49252 16998 49280 17054
rect 49240 16992 49292 16998
rect 49240 16934 49292 16940
rect 49332 16992 49384 16998
rect 49332 16934 49384 16940
rect 49240 16788 49292 16794
rect 49240 16730 49292 16736
rect 49252 16250 49280 16730
rect 49240 16244 49292 16250
rect 49240 16186 49292 16192
rect 49252 15638 49280 16186
rect 49240 15632 49292 15638
rect 49240 15574 49292 15580
rect 49344 15502 49372 16934
rect 49436 16794 49464 18770
rect 49424 16788 49476 16794
rect 49424 16730 49476 16736
rect 49424 15972 49476 15978
rect 49424 15914 49476 15920
rect 49436 15502 49464 15914
rect 49528 15910 49556 18770
rect 49792 18760 49844 18766
rect 49792 18702 49844 18708
rect 49606 18456 49662 18465
rect 49606 18391 49662 18400
rect 49620 18358 49648 18391
rect 49608 18352 49660 18358
rect 49608 18294 49660 18300
rect 49620 17882 49648 18294
rect 49804 18086 49832 18702
rect 49884 18624 49936 18630
rect 49884 18566 49936 18572
rect 49896 18426 49924 18566
rect 49884 18420 49936 18426
rect 49884 18362 49936 18368
rect 49792 18080 49844 18086
rect 49792 18022 49844 18028
rect 49608 17876 49660 17882
rect 49608 17818 49660 17824
rect 49608 17604 49660 17610
rect 49608 17546 49660 17552
rect 49620 16182 49648 17546
rect 49608 16176 49660 16182
rect 49608 16118 49660 16124
rect 49516 15904 49568 15910
rect 49516 15846 49568 15852
rect 49620 15586 49648 16118
rect 49528 15558 49648 15586
rect 49240 15496 49292 15502
rect 49240 15438 49292 15444
rect 49332 15496 49384 15502
rect 49332 15438 49384 15444
rect 49424 15496 49476 15502
rect 49424 15438 49476 15444
rect 49252 15162 49280 15438
rect 49528 15366 49556 15558
rect 49516 15360 49568 15366
rect 49516 15302 49568 15308
rect 49240 15156 49292 15162
rect 49240 15098 49292 15104
rect 49148 14612 49200 14618
rect 49148 14554 49200 14560
rect 49332 14408 49384 14414
rect 49332 14350 49384 14356
rect 49344 14074 49372 14350
rect 49332 14068 49384 14074
rect 49332 14010 49384 14016
rect 49240 13864 49292 13870
rect 49240 13806 49292 13812
rect 49332 13864 49384 13870
rect 49332 13806 49384 13812
rect 49148 13796 49200 13802
rect 49148 13738 49200 13744
rect 49160 13326 49188 13738
rect 49148 13320 49200 13326
rect 49148 13262 49200 13268
rect 48780 10804 48832 10810
rect 48780 10746 48832 10752
rect 49252 7206 49280 13806
rect 49344 13530 49372 13806
rect 49332 13524 49384 13530
rect 49332 13466 49384 13472
rect 49700 12776 49752 12782
rect 49700 12718 49752 12724
rect 49712 12442 49740 12718
rect 49700 12436 49752 12442
rect 49700 12378 49752 12384
rect 49608 12096 49660 12102
rect 49608 12038 49660 12044
rect 49620 11898 49648 12038
rect 49608 11892 49660 11898
rect 49608 11834 49660 11840
rect 49240 7200 49292 7206
rect 49240 7142 49292 7148
rect 49804 2650 49832 18022
rect 49988 16810 50016 20878
rect 50172 19530 50200 21490
rect 50540 21146 50568 21490
rect 50528 21140 50580 21146
rect 50528 21082 50580 21088
rect 50294 20700 50602 20709
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20635 50602 20644
rect 50632 20602 50660 23462
rect 51172 23248 51224 23254
rect 51224 23208 51304 23236
rect 51172 23190 51224 23196
rect 50804 22976 50856 22982
rect 50804 22918 50856 22924
rect 50816 22778 50844 22918
rect 50804 22772 50856 22778
rect 50804 22714 50856 22720
rect 50804 22568 50856 22574
rect 50804 22510 50856 22516
rect 50712 20868 50764 20874
rect 50712 20810 50764 20816
rect 50620 20596 50672 20602
rect 50620 20538 50672 20544
rect 50342 20496 50398 20505
rect 50342 20431 50398 20440
rect 50356 19854 50384 20431
rect 50344 19848 50396 19854
rect 50344 19790 50396 19796
rect 50436 19848 50488 19854
rect 50488 19796 50660 19802
rect 50436 19790 50660 19796
rect 50448 19774 50660 19790
rect 50294 19612 50602 19621
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19547 50602 19556
rect 50080 19502 50200 19530
rect 50632 19514 50660 19774
rect 50620 19508 50672 19514
rect 50080 17882 50108 19502
rect 50620 19450 50672 19456
rect 50160 19372 50212 19378
rect 50160 19314 50212 19320
rect 50068 17876 50120 17882
rect 50068 17818 50120 17824
rect 49896 16782 50016 16810
rect 49896 15706 49924 16782
rect 49976 16652 50028 16658
rect 49976 16594 50028 16600
rect 49988 16250 50016 16594
rect 49976 16244 50028 16250
rect 49976 16186 50028 16192
rect 49884 15700 49936 15706
rect 49884 15642 49936 15648
rect 50068 15496 50120 15502
rect 50068 15438 50120 15444
rect 49976 15428 50028 15434
rect 49976 15370 50028 15376
rect 49884 13932 49936 13938
rect 49884 13874 49936 13880
rect 49896 12238 49924 13874
rect 49988 13462 50016 15370
rect 50080 15162 50108 15438
rect 50172 15162 50200 19314
rect 50618 18864 50674 18873
rect 50618 18799 50674 18808
rect 50632 18766 50660 18799
rect 50620 18760 50672 18766
rect 50620 18702 50672 18708
rect 50294 18524 50602 18533
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18459 50602 18468
rect 50294 17436 50602 17445
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17371 50602 17380
rect 50294 16348 50602 16357
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16283 50602 16292
rect 50724 15706 50752 20810
rect 50816 18884 50844 22510
rect 51172 22024 51224 22030
rect 51172 21966 51224 21972
rect 51080 21616 51132 21622
rect 51080 21558 51132 21564
rect 50988 21548 51040 21554
rect 50988 21490 51040 21496
rect 51000 21146 51028 21490
rect 50988 21140 51040 21146
rect 50988 21082 51040 21088
rect 50988 20936 51040 20942
rect 50988 20878 51040 20884
rect 50896 19984 50948 19990
rect 50896 19926 50948 19932
rect 50908 19310 50936 19926
rect 51000 19378 51028 20878
rect 51092 20058 51120 21558
rect 51080 20052 51132 20058
rect 51080 19994 51132 20000
rect 51184 19718 51212 21966
rect 51276 20058 51304 23208
rect 51368 23118 51396 24006
rect 51920 23118 51948 24006
rect 52380 23118 52408 24550
rect 52472 23254 52500 24822
rect 52840 23798 52868 26250
rect 52920 24064 52972 24070
rect 52920 24006 52972 24012
rect 52828 23792 52880 23798
rect 52828 23734 52880 23740
rect 52932 23730 52960 24006
rect 52736 23724 52788 23730
rect 52736 23666 52788 23672
rect 52920 23724 52972 23730
rect 52920 23666 52972 23672
rect 52748 23322 52776 23666
rect 52736 23316 52788 23322
rect 52736 23258 52788 23264
rect 52460 23248 52512 23254
rect 52460 23190 52512 23196
rect 52472 23118 52500 23190
rect 51356 23112 51408 23118
rect 51356 23054 51408 23060
rect 51908 23112 51960 23118
rect 51908 23054 51960 23060
rect 52368 23112 52420 23118
rect 52368 23054 52420 23060
rect 52460 23112 52512 23118
rect 52460 23054 52512 23060
rect 51724 23044 51776 23050
rect 51724 22986 51776 22992
rect 51448 22976 51500 22982
rect 51448 22918 51500 22924
rect 51460 21418 51488 22918
rect 51736 22094 51764 22986
rect 52276 22976 52328 22982
rect 52276 22918 52328 22924
rect 51736 22066 51948 22094
rect 51448 21412 51500 21418
rect 51448 21354 51500 21360
rect 51448 20936 51500 20942
rect 51448 20878 51500 20884
rect 51460 20602 51488 20878
rect 51448 20596 51500 20602
rect 51448 20538 51500 20544
rect 51816 20256 51868 20262
rect 51816 20198 51868 20204
rect 51828 20058 51856 20198
rect 51264 20052 51316 20058
rect 51264 19994 51316 20000
rect 51816 20052 51868 20058
rect 51816 19994 51868 20000
rect 51172 19712 51224 19718
rect 51172 19654 51224 19660
rect 50988 19372 51040 19378
rect 50988 19314 51040 19320
rect 50896 19304 50948 19310
rect 50896 19246 50948 19252
rect 51172 19304 51224 19310
rect 51172 19246 51224 19252
rect 50988 18896 51040 18902
rect 50816 18856 50988 18884
rect 50988 18838 51040 18844
rect 51000 18086 51028 18838
rect 50988 18080 51040 18086
rect 50988 18022 51040 18028
rect 50896 16788 50948 16794
rect 51000 16776 51028 18022
rect 50948 16748 51028 16776
rect 50896 16730 50948 16736
rect 50712 15700 50764 15706
rect 50712 15642 50764 15648
rect 50804 15496 50856 15502
rect 50632 15444 50804 15450
rect 50632 15438 50856 15444
rect 50632 15422 50844 15438
rect 50294 15260 50602 15269
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15195 50602 15204
rect 50632 15162 50660 15422
rect 50068 15156 50120 15162
rect 50068 15098 50120 15104
rect 50160 15156 50212 15162
rect 50160 15098 50212 15104
rect 50620 15156 50672 15162
rect 50620 15098 50672 15104
rect 50436 15088 50488 15094
rect 50436 15030 50488 15036
rect 50068 15020 50120 15026
rect 50068 14962 50120 14968
rect 49976 13456 50028 13462
rect 49976 13398 50028 13404
rect 49976 13184 50028 13190
rect 49976 13126 50028 13132
rect 49988 12986 50016 13126
rect 49976 12980 50028 12986
rect 49976 12922 50028 12928
rect 50080 12850 50108 14962
rect 50448 14414 50476 15030
rect 50528 15020 50580 15026
rect 50632 15008 50660 15098
rect 50580 14980 50660 15008
rect 50528 14962 50580 14968
rect 50528 14816 50580 14822
rect 50528 14758 50580 14764
rect 50540 14618 50568 14758
rect 50632 14618 50660 14980
rect 50712 15020 50764 15026
rect 50712 14962 50764 14968
rect 50724 14618 50752 14962
rect 50528 14612 50580 14618
rect 50528 14554 50580 14560
rect 50620 14612 50672 14618
rect 50620 14554 50672 14560
rect 50712 14612 50764 14618
rect 50712 14554 50764 14560
rect 50436 14408 50488 14414
rect 50436 14350 50488 14356
rect 50294 14172 50602 14181
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14107 50602 14116
rect 50712 13184 50764 13190
rect 50712 13126 50764 13132
rect 50896 13184 50948 13190
rect 50896 13126 50948 13132
rect 50294 13084 50602 13093
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13019 50602 13028
rect 50620 12912 50672 12918
rect 50620 12854 50672 12860
rect 50068 12844 50120 12850
rect 50068 12786 50120 12792
rect 50632 12434 50660 12854
rect 50724 12850 50752 13126
rect 50908 12986 50936 13126
rect 50896 12980 50948 12986
rect 50896 12922 50948 12928
rect 50712 12844 50764 12850
rect 50712 12786 50764 12792
rect 50540 12406 50660 12434
rect 49884 12232 49936 12238
rect 49884 12174 49936 12180
rect 49896 11898 49924 12174
rect 50540 12170 50568 12406
rect 51000 12238 51028 16748
rect 51184 16590 51212 19246
rect 51276 18766 51304 19994
rect 51356 19848 51408 19854
rect 51356 19790 51408 19796
rect 51816 19848 51868 19854
rect 51816 19790 51868 19796
rect 51368 19514 51396 19790
rect 51632 19712 51684 19718
rect 51632 19654 51684 19660
rect 51356 19508 51408 19514
rect 51356 19450 51408 19456
rect 51644 19378 51672 19654
rect 51632 19372 51684 19378
rect 51632 19314 51684 19320
rect 51724 19372 51776 19378
rect 51724 19314 51776 19320
rect 51736 18970 51764 19314
rect 51724 18964 51776 18970
rect 51724 18906 51776 18912
rect 51264 18760 51316 18766
rect 51264 18702 51316 18708
rect 51632 18760 51684 18766
rect 51632 18702 51684 18708
rect 51724 18760 51776 18766
rect 51724 18702 51776 18708
rect 51540 18624 51592 18630
rect 51540 18566 51592 18572
rect 51552 18290 51580 18566
rect 51540 18284 51592 18290
rect 51540 18226 51592 18232
rect 51552 18154 51580 18226
rect 51540 18148 51592 18154
rect 51540 18090 51592 18096
rect 51356 18080 51408 18086
rect 51356 18022 51408 18028
rect 51368 17678 51396 18022
rect 51356 17672 51408 17678
rect 51356 17614 51408 17620
rect 51172 16584 51224 16590
rect 51172 16526 51224 16532
rect 51080 16108 51132 16114
rect 51080 16050 51132 16056
rect 51092 15994 51120 16050
rect 51184 15994 51212 16526
rect 51264 16448 51316 16454
rect 51264 16390 51316 16396
rect 51276 16114 51304 16390
rect 51264 16108 51316 16114
rect 51264 16050 51316 16056
rect 51092 15966 51212 15994
rect 51080 15428 51132 15434
rect 51080 15370 51132 15376
rect 51092 15162 51120 15370
rect 51080 15156 51132 15162
rect 51080 15098 51132 15104
rect 51184 12850 51212 15966
rect 51644 15706 51672 18702
rect 51736 18426 51764 18702
rect 51724 18420 51776 18426
rect 51724 18362 51776 18368
rect 51828 18290 51856 19790
rect 51920 19378 51948 22066
rect 52184 21956 52236 21962
rect 52184 21898 52236 21904
rect 52196 21690 52224 21898
rect 52184 21684 52236 21690
rect 52184 21626 52236 21632
rect 52288 20942 52316 22918
rect 52828 22772 52880 22778
rect 52828 22714 52880 22720
rect 52460 22432 52512 22438
rect 52460 22374 52512 22380
rect 52472 22030 52500 22374
rect 52460 22024 52512 22030
rect 52460 21966 52512 21972
rect 52368 21888 52420 21894
rect 52368 21830 52420 21836
rect 52736 21888 52788 21894
rect 52736 21830 52788 21836
rect 52276 20936 52328 20942
rect 52276 20878 52328 20884
rect 52380 20058 52408 21830
rect 52748 21690 52776 21830
rect 52736 21684 52788 21690
rect 52736 21626 52788 21632
rect 52840 20466 52868 22714
rect 53024 20534 53052 27270
rect 53116 25498 53144 29106
rect 53484 29073 53512 29106
rect 53470 29064 53526 29073
rect 53470 28999 53526 29008
rect 53196 28416 53248 28422
rect 53196 28358 53248 28364
rect 53288 28416 53340 28422
rect 53288 28358 53340 28364
rect 53208 27674 53236 28358
rect 53196 27668 53248 27674
rect 53196 27610 53248 27616
rect 53196 25832 53248 25838
rect 53196 25774 53248 25780
rect 53104 25492 53156 25498
rect 53104 25434 53156 25440
rect 53116 24954 53144 25434
rect 53104 24948 53156 24954
rect 53104 24890 53156 24896
rect 53116 22778 53144 24890
rect 53104 22772 53156 22778
rect 53104 22714 53156 22720
rect 53208 22438 53236 25774
rect 53300 24206 53328 28358
rect 53380 26784 53432 26790
rect 53380 26726 53432 26732
rect 53392 25294 53420 26726
rect 53472 26444 53524 26450
rect 53472 26386 53524 26392
rect 53484 26042 53512 26386
rect 53472 26036 53524 26042
rect 53472 25978 53524 25984
rect 53380 25288 53432 25294
rect 53380 25230 53432 25236
rect 53472 25152 53524 25158
rect 53472 25094 53524 25100
rect 53484 24954 53512 25094
rect 53472 24948 53524 24954
rect 53472 24890 53524 24896
rect 53576 24818 53604 29446
rect 53852 29306 53880 29514
rect 53840 29300 53892 29306
rect 53840 29242 53892 29248
rect 54588 29102 54616 30126
rect 54680 30054 54708 30194
rect 54668 30048 54720 30054
rect 54668 29990 54720 29996
rect 55140 29730 55168 31282
rect 55220 30252 55272 30258
rect 55220 30194 55272 30200
rect 55232 29850 55260 30194
rect 55220 29844 55272 29850
rect 55220 29786 55272 29792
rect 55048 29714 55168 29730
rect 55036 29708 55168 29714
rect 55088 29702 55168 29708
rect 55036 29650 55088 29656
rect 54576 29096 54628 29102
rect 54576 29038 54628 29044
rect 53656 28960 53708 28966
rect 53656 28902 53708 28908
rect 53668 28558 53696 28902
rect 53656 28552 53708 28558
rect 53656 28494 53708 28500
rect 53840 28212 53892 28218
rect 53840 28154 53892 28160
rect 53852 27470 53880 28154
rect 54024 28076 54076 28082
rect 54024 28018 54076 28024
rect 54036 27674 54064 28018
rect 54024 27668 54076 27674
rect 54024 27610 54076 27616
rect 53840 27464 53892 27470
rect 53840 27406 53892 27412
rect 53840 27328 53892 27334
rect 53840 27270 53892 27276
rect 53852 26874 53880 27270
rect 54588 27130 54616 29038
rect 55048 28994 55076 29650
rect 55128 29640 55180 29646
rect 55324 29594 55352 34886
rect 55496 34604 55548 34610
rect 55496 34546 55548 34552
rect 55508 33522 55536 34546
rect 55692 33658 55720 42570
rect 56796 41414 56824 43046
rect 57440 42770 57468 43182
rect 57060 42764 57112 42770
rect 57060 42706 57112 42712
rect 57428 42764 57480 42770
rect 57428 42706 57480 42712
rect 56876 42560 56928 42566
rect 56876 42502 56928 42508
rect 56612 41386 56824 41414
rect 56612 38654 56640 41386
rect 56244 38626 56640 38654
rect 56048 35216 56100 35222
rect 56048 35158 56100 35164
rect 55864 35080 55916 35086
rect 55864 35022 55916 35028
rect 55876 34610 55904 35022
rect 56060 34678 56088 35158
rect 56140 35080 56192 35086
rect 56140 35022 56192 35028
rect 56152 34746 56180 35022
rect 56140 34740 56192 34746
rect 56140 34682 56192 34688
rect 56244 34678 56272 38626
rect 56784 37664 56836 37670
rect 56784 37606 56836 37612
rect 56416 35488 56468 35494
rect 56416 35430 56468 35436
rect 56428 34950 56456 35430
rect 56416 34944 56468 34950
rect 56416 34886 56468 34892
rect 56048 34672 56100 34678
rect 56048 34614 56100 34620
rect 56232 34672 56284 34678
rect 56232 34614 56284 34620
rect 55864 34604 55916 34610
rect 55864 34546 55916 34552
rect 56324 34400 56376 34406
rect 56324 34342 56376 34348
rect 55680 33652 55732 33658
rect 55680 33594 55732 33600
rect 55496 33516 55548 33522
rect 55496 33458 55548 33464
rect 55508 33402 55536 33458
rect 55508 33374 55628 33402
rect 55496 33312 55548 33318
rect 55496 33254 55548 33260
rect 55508 32298 55536 33254
rect 55600 33114 55628 33374
rect 55588 33108 55640 33114
rect 55588 33050 55640 33056
rect 56336 32994 56364 34342
rect 56428 34202 56456 34886
rect 56692 34740 56744 34746
rect 56692 34682 56744 34688
rect 56704 34610 56732 34682
rect 56692 34604 56744 34610
rect 56692 34546 56744 34552
rect 56508 34468 56560 34474
rect 56508 34410 56560 34416
rect 56416 34196 56468 34202
rect 56416 34138 56468 34144
rect 56520 33130 56548 34410
rect 56600 33856 56652 33862
rect 56600 33798 56652 33804
rect 56612 33658 56640 33798
rect 56600 33652 56652 33658
rect 56600 33594 56652 33600
rect 56600 33516 56652 33522
rect 56600 33458 56652 33464
rect 56244 32966 56364 32994
rect 56428 33102 56548 33130
rect 56612 33114 56640 33458
rect 56600 33108 56652 33114
rect 55588 32360 55640 32366
rect 55588 32302 55640 32308
rect 55496 32292 55548 32298
rect 55496 32234 55548 32240
rect 55600 32026 55628 32302
rect 55588 32020 55640 32026
rect 55588 31962 55640 31968
rect 56140 31136 56192 31142
rect 56140 31078 56192 31084
rect 55864 30048 55916 30054
rect 55864 29990 55916 29996
rect 55128 29582 55180 29588
rect 55140 29306 55168 29582
rect 55232 29566 55352 29594
rect 55128 29300 55180 29306
rect 55128 29242 55180 29248
rect 54864 28966 55076 28994
rect 54864 27470 54892 28966
rect 55232 28694 55260 29566
rect 55312 29504 55364 29510
rect 55312 29446 55364 29452
rect 55404 29504 55456 29510
rect 55404 29446 55456 29452
rect 55324 29306 55352 29446
rect 55312 29300 55364 29306
rect 55312 29242 55364 29248
rect 55416 29102 55444 29446
rect 55876 29306 55904 29990
rect 56048 29572 56100 29578
rect 56048 29514 56100 29520
rect 56060 29306 56088 29514
rect 55864 29300 55916 29306
rect 55864 29242 55916 29248
rect 56048 29300 56100 29306
rect 56048 29242 56100 29248
rect 56152 29170 56180 31078
rect 56140 29164 56192 29170
rect 56140 29106 56192 29112
rect 55404 29096 55456 29102
rect 55404 29038 55456 29044
rect 55864 28960 55916 28966
rect 55864 28902 55916 28908
rect 55220 28688 55272 28694
rect 55220 28630 55272 28636
rect 55876 28558 55904 28902
rect 55864 28552 55916 28558
rect 55864 28494 55916 28500
rect 55680 28008 55732 28014
rect 55680 27950 55732 27956
rect 55036 27872 55088 27878
rect 55036 27814 55088 27820
rect 55048 27470 55076 27814
rect 55692 27674 55720 27950
rect 55876 27878 55904 28494
rect 55864 27872 55916 27878
rect 55864 27814 55916 27820
rect 55680 27668 55732 27674
rect 55680 27610 55732 27616
rect 55876 27470 55904 27814
rect 56152 27538 56180 29106
rect 56140 27532 56192 27538
rect 56140 27474 56192 27480
rect 54852 27464 54904 27470
rect 54852 27406 54904 27412
rect 55036 27464 55088 27470
rect 55036 27406 55088 27412
rect 55864 27464 55916 27470
rect 55864 27406 55916 27412
rect 54116 27124 54168 27130
rect 54116 27066 54168 27072
rect 54576 27124 54628 27130
rect 54576 27066 54628 27072
rect 53932 26988 53984 26994
rect 53932 26930 53984 26936
rect 53668 26858 53880 26874
rect 53656 26852 53880 26858
rect 53708 26846 53880 26852
rect 53656 26794 53708 26800
rect 53944 26772 53972 26930
rect 53760 26744 53972 26772
rect 53760 26586 53788 26744
rect 53748 26580 53800 26586
rect 53748 26522 53800 26528
rect 53840 26580 53892 26586
rect 53840 26522 53892 26528
rect 53656 26512 53708 26518
rect 53852 26466 53880 26522
rect 53708 26460 53880 26466
rect 53656 26454 53880 26460
rect 53668 26438 53880 26454
rect 53748 26376 53800 26382
rect 53748 26318 53800 26324
rect 53840 26376 53892 26382
rect 53840 26318 53892 26324
rect 53760 26246 53788 26318
rect 53748 26240 53800 26246
rect 53748 26182 53800 26188
rect 53852 25974 53880 26318
rect 54128 26246 54156 27066
rect 54484 26920 54536 26926
rect 54484 26862 54536 26868
rect 54496 26586 54524 26862
rect 54484 26580 54536 26586
rect 54484 26522 54536 26528
rect 54588 26382 54616 27066
rect 54864 26994 54892 27406
rect 56152 27334 56180 27474
rect 56244 27441 56272 32966
rect 56428 32910 56456 33102
rect 56600 33050 56652 33056
rect 56508 33040 56560 33046
rect 56508 32982 56560 32988
rect 56416 32904 56468 32910
rect 56416 32846 56468 32852
rect 56520 32314 56548 32982
rect 56796 32774 56824 37606
rect 56888 34610 56916 42502
rect 57072 42022 57100 42706
rect 57532 42702 57560 43658
rect 57808 43382 57836 47942
rect 58360 46458 58388 49030
rect 58176 46430 58388 46458
rect 57888 45960 57940 45966
rect 57888 45902 57940 45908
rect 57900 45529 57928 45902
rect 57886 45520 57942 45529
rect 57886 45455 57942 45464
rect 57980 44192 58032 44198
rect 57980 44134 58032 44140
rect 57992 43654 58020 44134
rect 58072 43988 58124 43994
rect 58072 43930 58124 43936
rect 57980 43648 58032 43654
rect 57980 43590 58032 43596
rect 57796 43376 57848 43382
rect 57796 43318 57848 43324
rect 57520 42696 57572 42702
rect 57520 42638 57572 42644
rect 57808 42634 57836 43318
rect 57796 42628 57848 42634
rect 57796 42570 57848 42576
rect 57992 42362 58020 43590
rect 58084 43450 58112 43930
rect 58176 43450 58204 46430
rect 58348 46368 58400 46374
rect 58348 46310 58400 46316
rect 58360 45914 58388 46310
rect 58360 45886 58480 45914
rect 58348 45824 58400 45830
rect 58348 45766 58400 45772
rect 58360 43858 58388 45766
rect 58348 43852 58400 43858
rect 58348 43794 58400 43800
rect 58256 43648 58308 43654
rect 58256 43590 58308 43596
rect 58072 43444 58124 43450
rect 58072 43386 58124 43392
rect 58164 43444 58216 43450
rect 58164 43386 58216 43392
rect 58084 42906 58112 43386
rect 58072 42900 58124 42906
rect 58072 42842 58124 42848
rect 58176 42770 58204 43386
rect 58164 42764 58216 42770
rect 58164 42706 58216 42712
rect 58072 42560 58124 42566
rect 58072 42502 58124 42508
rect 57980 42356 58032 42362
rect 57980 42298 58032 42304
rect 56968 42016 57020 42022
rect 56968 41958 57020 41964
rect 57060 42016 57112 42022
rect 57060 41958 57112 41964
rect 56980 35086 57008 41958
rect 57072 39506 57100 41958
rect 58084 41154 58112 42502
rect 58164 41472 58216 41478
rect 58164 41414 58216 41420
rect 58176 41274 58204 41414
rect 58164 41268 58216 41274
rect 58164 41210 58216 41216
rect 57980 41132 58032 41138
rect 58084 41126 58204 41154
rect 58268 41138 58296 43590
rect 58360 42702 58388 43794
rect 58452 43246 58480 45886
rect 58440 43240 58492 43246
rect 58440 43182 58492 43188
rect 58532 43104 58584 43110
rect 58532 43046 58584 43052
rect 58348 42696 58400 42702
rect 58348 42638 58400 42644
rect 58348 41472 58400 41478
rect 58348 41414 58400 41420
rect 57980 41074 58032 41080
rect 57992 40186 58020 41074
rect 58176 41070 58204 41126
rect 58256 41132 58308 41138
rect 58256 41074 58308 41080
rect 58164 41064 58216 41070
rect 58164 41006 58216 41012
rect 58072 40928 58124 40934
rect 58072 40870 58124 40876
rect 58084 40730 58112 40870
rect 58072 40724 58124 40730
rect 58072 40666 58124 40672
rect 57980 40180 58032 40186
rect 57980 40122 58032 40128
rect 57888 40112 57940 40118
rect 57888 40054 57940 40060
rect 57796 39908 57848 39914
rect 57796 39850 57848 39856
rect 57808 39817 57836 39850
rect 57794 39808 57850 39817
rect 57794 39743 57850 39752
rect 57060 39500 57112 39506
rect 57060 39442 57112 39448
rect 57900 39438 57928 40054
rect 58072 39636 58124 39642
rect 58072 39578 58124 39584
rect 57888 39432 57940 39438
rect 57888 39374 57940 39380
rect 57336 39296 57388 39302
rect 57336 39238 57388 39244
rect 57612 39296 57664 39302
rect 57612 39238 57664 39244
rect 57348 38758 57376 39238
rect 57336 38752 57388 38758
rect 57336 38694 57388 38700
rect 57244 38480 57296 38486
rect 57244 38422 57296 38428
rect 57256 35086 57284 38422
rect 57348 38214 57376 38694
rect 57336 38208 57388 38214
rect 57336 38150 57388 38156
rect 56968 35080 57020 35086
rect 56968 35022 57020 35028
rect 57060 35080 57112 35086
rect 57060 35022 57112 35028
rect 57244 35080 57296 35086
rect 57244 35022 57296 35028
rect 56876 34604 56928 34610
rect 56876 34546 56928 34552
rect 57072 33998 57100 35022
rect 57060 33992 57112 33998
rect 57060 33934 57112 33940
rect 57348 33658 57376 38150
rect 57520 36304 57572 36310
rect 57520 36246 57572 36252
rect 57532 34610 57560 36246
rect 57520 34604 57572 34610
rect 57520 34546 57572 34552
rect 57624 33998 57652 39238
rect 58084 39098 58112 39578
rect 58176 39438 58204 41006
rect 58256 40928 58308 40934
rect 58256 40870 58308 40876
rect 58268 40730 58296 40870
rect 58256 40724 58308 40730
rect 58256 40666 58308 40672
rect 58360 40118 58388 41414
rect 58440 41132 58492 41138
rect 58440 41074 58492 41080
rect 58348 40112 58400 40118
rect 58348 40054 58400 40060
rect 58360 39438 58388 40054
rect 58164 39432 58216 39438
rect 58164 39374 58216 39380
rect 58348 39432 58400 39438
rect 58348 39374 58400 39380
rect 58256 39296 58308 39302
rect 58256 39238 58308 39244
rect 58072 39092 58124 39098
rect 58072 39034 58124 39040
rect 57980 38956 58032 38962
rect 57980 38898 58032 38904
rect 57992 38282 58020 38898
rect 57980 38276 58032 38282
rect 57980 38218 58032 38224
rect 57704 36576 57756 36582
rect 57704 36518 57756 36524
rect 57980 36576 58032 36582
rect 57980 36518 58032 36524
rect 57716 35494 57744 36518
rect 57992 36378 58020 36518
rect 57980 36372 58032 36378
rect 57980 36314 58032 36320
rect 58084 35698 58112 39034
rect 58268 39001 58296 39238
rect 58254 38992 58310 39001
rect 58254 38927 58310 38936
rect 58256 38820 58308 38826
rect 58256 38762 58308 38768
rect 58164 38752 58216 38758
rect 58164 38694 58216 38700
rect 58176 37670 58204 38694
rect 58268 38418 58296 38762
rect 58256 38412 58308 38418
rect 58256 38354 58308 38360
rect 58348 38276 58400 38282
rect 58348 38218 58400 38224
rect 58360 38185 58388 38218
rect 58346 38176 58402 38185
rect 58346 38111 58402 38120
rect 58452 38010 58480 41074
rect 58544 40526 58572 43046
rect 58532 40520 58584 40526
rect 58532 40462 58584 40468
rect 58532 39296 58584 39302
rect 58532 39238 58584 39244
rect 58440 38004 58492 38010
rect 58440 37946 58492 37952
rect 58256 37868 58308 37874
rect 58256 37810 58308 37816
rect 58164 37664 58216 37670
rect 58164 37606 58216 37612
rect 58268 37466 58296 37810
rect 58256 37460 58308 37466
rect 58256 37402 58308 37408
rect 58268 36922 58296 37402
rect 58256 36916 58308 36922
rect 58256 36858 58308 36864
rect 58164 36576 58216 36582
rect 58164 36518 58216 36524
rect 58072 35692 58124 35698
rect 58072 35634 58124 35640
rect 57704 35488 57756 35494
rect 57704 35430 57756 35436
rect 57888 35488 57940 35494
rect 57888 35430 57940 35436
rect 57716 35154 57744 35430
rect 57704 35148 57756 35154
rect 57704 35090 57756 35096
rect 57796 34060 57848 34066
rect 57796 34002 57848 34008
rect 57612 33992 57664 33998
rect 57612 33934 57664 33940
rect 57520 33856 57572 33862
rect 57520 33798 57572 33804
rect 57336 33652 57388 33658
rect 57336 33594 57388 33600
rect 57348 33436 57376 33594
rect 57532 33454 57560 33798
rect 57808 33522 57836 34002
rect 57900 33998 57928 35430
rect 57980 34536 58032 34542
rect 57980 34478 58032 34484
rect 57992 34202 58020 34478
rect 57980 34196 58032 34202
rect 57980 34138 58032 34144
rect 57888 33992 57940 33998
rect 57888 33934 57940 33940
rect 57980 33924 58032 33930
rect 57980 33866 58032 33872
rect 57992 33810 58020 33866
rect 57900 33782 58020 33810
rect 57796 33516 57848 33522
rect 57796 33458 57848 33464
rect 57520 33448 57572 33454
rect 57348 33408 57520 33436
rect 57520 33390 57572 33396
rect 57704 33448 57756 33454
rect 57704 33390 57756 33396
rect 56968 33312 57020 33318
rect 56968 33254 57020 33260
rect 57336 33312 57388 33318
rect 57336 33254 57388 33260
rect 56980 32910 57008 33254
rect 57348 32910 57376 33254
rect 57716 33114 57744 33390
rect 57704 33108 57756 33114
rect 57704 33050 57756 33056
rect 57900 33046 57928 33782
rect 58176 33658 58204 36518
rect 58544 36378 58572 39238
rect 58532 36372 58584 36378
rect 58532 36314 58584 36320
rect 58440 36100 58492 36106
rect 58440 36042 58492 36048
rect 58348 36032 58400 36038
rect 58348 35974 58400 35980
rect 58360 35766 58388 35974
rect 58348 35760 58400 35766
rect 58348 35702 58400 35708
rect 58452 35698 58480 36042
rect 58440 35692 58492 35698
rect 58440 35634 58492 35640
rect 58348 34400 58400 34406
rect 58348 34342 58400 34348
rect 58360 34202 58388 34342
rect 58348 34196 58400 34202
rect 58348 34138 58400 34144
rect 58452 33930 58480 35634
rect 58440 33924 58492 33930
rect 58440 33866 58492 33872
rect 58164 33652 58216 33658
rect 58164 33594 58216 33600
rect 57888 33040 57940 33046
rect 57888 32982 57940 32988
rect 56968 32904 57020 32910
rect 56968 32846 57020 32852
rect 57336 32904 57388 32910
rect 57336 32846 57388 32852
rect 56784 32768 56836 32774
rect 56784 32710 56836 32716
rect 56336 32286 56548 32314
rect 56336 28665 56364 32286
rect 56508 31816 56560 31822
rect 56508 31758 56560 31764
rect 56520 29850 56548 31758
rect 58636 31754 58664 52634
rect 58900 52420 58952 52426
rect 58900 52362 58952 52368
rect 58912 52057 58940 52362
rect 58898 52048 58954 52057
rect 58898 51983 58954 51992
rect 58900 51332 58952 51338
rect 58900 51274 58952 51280
rect 58716 51264 58768 51270
rect 58912 51241 58940 51274
rect 58716 51206 58768 51212
rect 58898 51232 58954 51241
rect 56876 31748 56928 31754
rect 56876 31690 56928 31696
rect 58544 31726 58664 31754
rect 56692 31680 56744 31686
rect 56692 31622 56744 31628
rect 56704 31278 56732 31622
rect 56888 31482 56916 31690
rect 58164 31680 58216 31686
rect 58164 31622 58216 31628
rect 58348 31680 58400 31686
rect 58348 31622 58400 31628
rect 56876 31476 56928 31482
rect 56876 31418 56928 31424
rect 56968 31408 57020 31414
rect 56968 31350 57020 31356
rect 56692 31272 56744 31278
rect 56692 31214 56744 31220
rect 56980 30938 57008 31350
rect 58176 31346 58204 31622
rect 57336 31340 57388 31346
rect 57336 31282 57388 31288
rect 58164 31340 58216 31346
rect 58164 31282 58216 31288
rect 57348 30938 57376 31282
rect 56968 30932 57020 30938
rect 56968 30874 57020 30880
rect 57336 30932 57388 30938
rect 57336 30874 57388 30880
rect 58360 30734 58388 31622
rect 58348 30728 58400 30734
rect 58348 30670 58400 30676
rect 57244 30592 57296 30598
rect 57244 30534 57296 30540
rect 57612 30592 57664 30598
rect 57612 30534 57664 30540
rect 58072 30592 58124 30598
rect 58072 30534 58124 30540
rect 56508 29844 56560 29850
rect 56508 29786 56560 29792
rect 56416 29164 56468 29170
rect 56416 29106 56468 29112
rect 56322 28656 56378 28665
rect 56322 28591 56378 28600
rect 56428 28558 56456 29106
rect 56416 28552 56468 28558
rect 56416 28494 56468 28500
rect 56520 28150 56548 29786
rect 57256 29646 57284 30534
rect 57520 30252 57572 30258
rect 57520 30194 57572 30200
rect 57532 29850 57560 30194
rect 57520 29844 57572 29850
rect 57520 29786 57572 29792
rect 56968 29640 57020 29646
rect 56968 29582 57020 29588
rect 57244 29640 57296 29646
rect 57244 29582 57296 29588
rect 56980 29306 57008 29582
rect 57624 29578 57652 30534
rect 57796 30388 57848 30394
rect 57796 30330 57848 30336
rect 57808 29646 57836 30330
rect 58084 30258 58112 30534
rect 58544 30258 58572 31726
rect 58622 30832 58678 30841
rect 58622 30767 58624 30776
rect 58676 30767 58678 30776
rect 58624 30738 58676 30744
rect 58072 30252 58124 30258
rect 58072 30194 58124 30200
rect 58532 30252 58584 30258
rect 58532 30194 58584 30200
rect 58624 30116 58676 30122
rect 58624 30058 58676 30064
rect 58072 30048 58124 30054
rect 58636 30025 58664 30058
rect 58072 29990 58124 29996
rect 58622 30016 58678 30025
rect 57796 29640 57848 29646
rect 57796 29582 57848 29588
rect 57612 29572 57664 29578
rect 57612 29514 57664 29520
rect 57060 29504 57112 29510
rect 57060 29446 57112 29452
rect 57072 29306 57100 29446
rect 56968 29300 57020 29306
rect 56968 29242 57020 29248
rect 57060 29300 57112 29306
rect 57060 29242 57112 29248
rect 57244 29164 57296 29170
rect 57244 29106 57296 29112
rect 57428 29164 57480 29170
rect 57428 29106 57480 29112
rect 57150 29064 57206 29073
rect 56692 29028 56744 29034
rect 57256 29050 57284 29106
rect 57206 29022 57284 29050
rect 57150 28999 57206 29008
rect 56692 28970 56744 28976
rect 56600 28416 56652 28422
rect 56600 28358 56652 28364
rect 56508 28144 56560 28150
rect 56508 28086 56560 28092
rect 56416 28076 56468 28082
rect 56416 28018 56468 28024
rect 56428 27674 56456 28018
rect 56416 27668 56468 27674
rect 56416 27610 56468 27616
rect 56416 27464 56468 27470
rect 56230 27432 56286 27441
rect 56416 27406 56468 27412
rect 56230 27367 56286 27376
rect 54944 27328 54996 27334
rect 54944 27270 54996 27276
rect 56140 27328 56192 27334
rect 56140 27270 56192 27276
rect 56324 27328 56376 27334
rect 56324 27270 56376 27276
rect 54852 26988 54904 26994
rect 54852 26930 54904 26936
rect 54956 26586 54984 27270
rect 56336 26926 56364 27270
rect 56048 26920 56100 26926
rect 56048 26862 56100 26868
rect 56324 26920 56376 26926
rect 56324 26862 56376 26868
rect 55404 26784 55456 26790
rect 55404 26726 55456 26732
rect 54760 26580 54812 26586
rect 54760 26522 54812 26528
rect 54944 26580 54996 26586
rect 54944 26522 54996 26528
rect 54484 26376 54536 26382
rect 54484 26318 54536 26324
rect 54576 26376 54628 26382
rect 54576 26318 54628 26324
rect 54208 26308 54260 26314
rect 54208 26250 54260 26256
rect 54116 26240 54168 26246
rect 54116 26182 54168 26188
rect 53840 25968 53892 25974
rect 53840 25910 53892 25916
rect 53748 25492 53800 25498
rect 53748 25434 53800 25440
rect 53760 25294 53788 25434
rect 53748 25288 53800 25294
rect 53748 25230 53800 25236
rect 53760 24954 53788 25230
rect 53840 25220 53892 25226
rect 53840 25162 53892 25168
rect 53748 24948 53800 24954
rect 53748 24890 53800 24896
rect 53380 24812 53432 24818
rect 53380 24754 53432 24760
rect 53564 24812 53616 24818
rect 53564 24754 53616 24760
rect 53392 24206 53420 24754
rect 53288 24200 53340 24206
rect 53288 24142 53340 24148
rect 53380 24200 53432 24206
rect 53380 24142 53432 24148
rect 53852 23866 53880 25162
rect 54128 24834 54156 26182
rect 54220 26042 54248 26250
rect 54300 26240 54352 26246
rect 54300 26182 54352 26188
rect 54208 26036 54260 26042
rect 54208 25978 54260 25984
rect 54312 25294 54340 26182
rect 54496 25362 54524 26318
rect 54484 25356 54536 25362
rect 54484 25298 54536 25304
rect 54300 25288 54352 25294
rect 54300 25230 54352 25236
rect 54128 24806 54340 24834
rect 54208 24064 54260 24070
rect 54208 24006 54260 24012
rect 53840 23860 53892 23866
rect 53840 23802 53892 23808
rect 54220 23730 54248 24006
rect 54312 23730 54340 24806
rect 54772 24750 54800 26522
rect 55312 26512 55364 26518
rect 55312 26454 55364 26460
rect 55220 26376 55272 26382
rect 55220 26318 55272 26324
rect 54852 26240 54904 26246
rect 54852 26182 54904 26188
rect 55036 26240 55088 26246
rect 55036 26182 55088 26188
rect 54864 25430 54892 26182
rect 54852 25424 54904 25430
rect 54852 25366 54904 25372
rect 54944 25356 54996 25362
rect 54944 25298 54996 25304
rect 54760 24744 54812 24750
rect 54760 24686 54812 24692
rect 53932 23724 53984 23730
rect 53932 23666 53984 23672
rect 54208 23724 54260 23730
rect 54208 23666 54260 23672
rect 54300 23724 54352 23730
rect 54300 23666 54352 23672
rect 54392 23724 54444 23730
rect 54392 23666 54444 23672
rect 53472 23112 53524 23118
rect 53472 23054 53524 23060
rect 53484 22778 53512 23054
rect 53472 22772 53524 22778
rect 53472 22714 53524 22720
rect 53196 22432 53248 22438
rect 53196 22374 53248 22380
rect 53564 22024 53616 22030
rect 53564 21966 53616 21972
rect 53576 21554 53604 21966
rect 53944 21894 53972 23666
rect 54312 22166 54340 23666
rect 54404 22982 54432 23666
rect 54484 23520 54536 23526
rect 54484 23462 54536 23468
rect 54496 23118 54524 23462
rect 54484 23112 54536 23118
rect 54484 23054 54536 23060
rect 54392 22976 54444 22982
rect 54392 22918 54444 22924
rect 54772 22760 54800 24686
rect 54852 24608 54904 24614
rect 54852 24550 54904 24556
rect 54864 23866 54892 24550
rect 54852 23860 54904 23866
rect 54852 23802 54904 23808
rect 54956 23730 54984 25298
rect 55048 25226 55076 26182
rect 55036 25220 55088 25226
rect 55036 25162 55088 25168
rect 55048 24342 55076 25162
rect 55232 24834 55260 26318
rect 55324 26042 55352 26454
rect 55312 26036 55364 26042
rect 55312 25978 55364 25984
rect 55416 25906 55444 26726
rect 56060 26586 56088 26862
rect 56048 26580 56100 26586
rect 56048 26522 56100 26528
rect 55404 25900 55456 25906
rect 55404 25842 55456 25848
rect 56336 25838 56364 26862
rect 56428 26330 56456 27406
rect 56520 26450 56548 28086
rect 56612 27470 56640 28358
rect 56600 27464 56652 27470
rect 56600 27406 56652 27412
rect 56508 26444 56560 26450
rect 56508 26386 56560 26392
rect 56428 26302 56640 26330
rect 56324 25832 56376 25838
rect 56324 25774 56376 25780
rect 56508 25832 56560 25838
rect 56508 25774 56560 25780
rect 56232 25288 56284 25294
rect 56232 25230 56284 25236
rect 55312 25152 55364 25158
rect 55312 25094 55364 25100
rect 55140 24818 55260 24834
rect 55128 24812 55260 24818
rect 55180 24806 55260 24812
rect 55128 24754 55180 24760
rect 55324 24614 55352 25094
rect 56048 24676 56100 24682
rect 56048 24618 56100 24624
rect 55312 24608 55364 24614
rect 55312 24550 55364 24556
rect 55956 24608 56008 24614
rect 55956 24550 56008 24556
rect 55036 24336 55088 24342
rect 55036 24278 55088 24284
rect 55968 24274 55996 24550
rect 55956 24268 56008 24274
rect 55956 24210 56008 24216
rect 54944 23724 54996 23730
rect 54944 23666 54996 23672
rect 54680 22732 54800 22760
rect 54300 22160 54352 22166
rect 54300 22102 54352 22108
rect 54484 22094 54536 22098
rect 54680 22094 54708 22732
rect 54760 22636 54812 22642
rect 54760 22578 54812 22584
rect 54772 22234 54800 22578
rect 54760 22228 54812 22234
rect 54760 22170 54812 22176
rect 54484 22092 54708 22094
rect 54536 22066 54708 22092
rect 54484 22034 54536 22040
rect 54024 22024 54076 22030
rect 54024 21966 54076 21972
rect 54116 22024 54168 22030
rect 54116 21966 54168 21972
rect 53932 21888 53984 21894
rect 53932 21830 53984 21836
rect 53564 21548 53616 21554
rect 53564 21490 53616 21496
rect 53012 20528 53064 20534
rect 53012 20470 53064 20476
rect 52828 20460 52880 20466
rect 52828 20402 52880 20408
rect 52368 20052 52420 20058
rect 52368 19994 52420 20000
rect 51908 19372 51960 19378
rect 51908 19314 51960 19320
rect 52276 19168 52328 19174
rect 52276 19110 52328 19116
rect 51908 18964 51960 18970
rect 51908 18906 51960 18912
rect 51724 18284 51776 18290
rect 51724 18226 51776 18232
rect 51816 18284 51868 18290
rect 51816 18226 51868 18232
rect 51736 18170 51764 18226
rect 51920 18170 51948 18906
rect 52288 18834 52316 19110
rect 52276 18828 52328 18834
rect 52276 18770 52328 18776
rect 52276 18624 52328 18630
rect 52276 18566 52328 18572
rect 52288 18426 52316 18566
rect 52276 18420 52328 18426
rect 52276 18362 52328 18368
rect 51736 18142 51948 18170
rect 52736 17536 52788 17542
rect 52736 17478 52788 17484
rect 52748 16998 52776 17478
rect 52736 16992 52788 16998
rect 52736 16934 52788 16940
rect 52748 16658 52776 16934
rect 52840 16794 52868 20402
rect 52920 20256 52972 20262
rect 52920 20198 52972 20204
rect 52932 16794 52960 20198
rect 52828 16788 52880 16794
rect 52828 16730 52880 16736
rect 52920 16788 52972 16794
rect 52920 16730 52972 16736
rect 52736 16652 52788 16658
rect 52736 16594 52788 16600
rect 51816 16516 51868 16522
rect 51816 16458 51868 16464
rect 51828 15910 51856 16458
rect 52552 16448 52604 16454
rect 52552 16390 52604 16396
rect 52564 16046 52592 16390
rect 52552 16040 52604 16046
rect 52552 15982 52604 15988
rect 51816 15904 51868 15910
rect 51816 15846 51868 15852
rect 51632 15700 51684 15706
rect 51632 15642 51684 15648
rect 51828 15570 51856 15846
rect 52748 15638 52776 16594
rect 52920 16516 52972 16522
rect 52920 16458 52972 16464
rect 52828 16448 52880 16454
rect 52828 16390 52880 16396
rect 52840 16250 52868 16390
rect 52828 16244 52880 16250
rect 52828 16186 52880 16192
rect 52932 15706 52960 16458
rect 52920 15700 52972 15706
rect 52920 15642 52972 15648
rect 52736 15632 52788 15638
rect 52736 15574 52788 15580
rect 51816 15564 51868 15570
rect 51816 15506 51868 15512
rect 51632 15496 51684 15502
rect 51632 15438 51684 15444
rect 52828 15496 52880 15502
rect 52828 15438 52880 15444
rect 51644 15162 51672 15438
rect 52840 15162 52868 15438
rect 53024 15162 53052 20470
rect 54036 19854 54064 21966
rect 54128 21690 54156 21966
rect 54484 21956 54536 21962
rect 54484 21898 54536 21904
rect 54208 21888 54260 21894
rect 54208 21830 54260 21836
rect 54116 21684 54168 21690
rect 54116 21626 54168 21632
rect 54220 19854 54248 21830
rect 54496 21690 54524 21898
rect 54484 21684 54536 21690
rect 54484 21626 54536 21632
rect 54588 21146 54616 22066
rect 54956 22030 54984 23666
rect 55312 23112 55364 23118
rect 55312 23054 55364 23060
rect 55324 22778 55352 23054
rect 56060 22982 56088 24618
rect 56244 24342 56272 25230
rect 56232 24336 56284 24342
rect 56232 24278 56284 24284
rect 56520 24206 56548 25774
rect 56612 25226 56640 26302
rect 56600 25220 56652 25226
rect 56600 25162 56652 25168
rect 56704 24410 56732 28970
rect 57164 28762 57192 28999
rect 57440 28762 57468 29106
rect 57152 28756 57204 28762
rect 57152 28698 57204 28704
rect 57428 28756 57480 28762
rect 57428 28698 57480 28704
rect 57624 28558 57652 29514
rect 57808 28558 57836 29582
rect 58084 29306 58112 29990
rect 58622 29951 58678 29960
rect 58728 29782 58756 51206
rect 58898 51167 58954 51176
rect 58808 49768 58860 49774
rect 58808 49710 58860 49716
rect 58900 49768 58952 49774
rect 58900 49710 58952 49716
rect 58820 43178 58848 49710
rect 58912 49609 58940 49710
rect 58898 49600 58954 49609
rect 58898 49535 58954 49544
rect 58900 49088 58952 49094
rect 58900 49030 58952 49036
rect 58912 48793 58940 49030
rect 58898 48784 58954 48793
rect 58898 48719 58954 48728
rect 58900 48068 58952 48074
rect 58900 48010 58952 48016
rect 58912 47977 58940 48010
rect 58898 47968 58954 47977
rect 58898 47903 58954 47912
rect 58900 47660 58952 47666
rect 58900 47602 58952 47608
rect 58912 47161 58940 47602
rect 58898 47152 58954 47161
rect 58898 47087 58954 47096
rect 58900 46436 58952 46442
rect 58900 46378 58952 46384
rect 58912 46345 58940 46378
rect 58898 46336 58954 46345
rect 58898 46271 58954 46280
rect 59004 45554 59032 52838
rect 59084 47456 59136 47462
rect 59084 47398 59136 47404
rect 58912 45526 59032 45554
rect 58808 43172 58860 43178
rect 58808 43114 58860 43120
rect 58806 43072 58862 43081
rect 58806 43007 58862 43016
rect 58820 42906 58848 43007
rect 58808 42900 58860 42906
rect 58808 42842 58860 42848
rect 58808 41540 58860 41546
rect 58808 41482 58860 41488
rect 58820 41449 58848 41482
rect 58806 41440 58862 41449
rect 58806 41375 58862 41384
rect 58808 40996 58860 41002
rect 58808 40938 58860 40944
rect 58820 38486 58848 40938
rect 58808 38480 58860 38486
rect 58808 38422 58860 38428
rect 58912 37482 58940 45526
rect 58992 44804 59044 44810
rect 58992 44746 59044 44752
rect 59004 44713 59032 44746
rect 58990 44704 59046 44713
rect 58990 44639 59046 44648
rect 58992 44192 59044 44198
rect 58992 44134 59044 44140
rect 59004 43897 59032 44134
rect 58990 43888 59046 43897
rect 58990 43823 59046 43832
rect 59096 43314 59124 47398
rect 59084 43308 59136 43314
rect 59084 43250 59136 43256
rect 58992 42696 59044 42702
rect 58992 42638 59044 42644
rect 59004 42265 59032 42638
rect 59096 42362 59124 43250
rect 59176 43172 59228 43178
rect 59176 43114 59228 43120
rect 59084 42356 59136 42362
rect 59084 42298 59136 42304
rect 58990 42256 59046 42265
rect 58990 42191 59046 42200
rect 58992 41472 59044 41478
rect 58992 41414 59044 41420
rect 59004 40633 59032 41414
rect 58990 40624 59046 40633
rect 58990 40559 59046 40568
rect 59188 37942 59216 43114
rect 59176 37936 59228 37942
rect 59176 37878 59228 37884
rect 58820 37454 58940 37482
rect 58716 29776 58768 29782
rect 58716 29718 58768 29724
rect 58532 29504 58584 29510
rect 58532 29446 58584 29452
rect 58072 29300 58124 29306
rect 58072 29242 58124 29248
rect 58544 29209 58572 29446
rect 58530 29200 58586 29209
rect 58530 29135 58586 29144
rect 57612 28552 57664 28558
rect 57612 28494 57664 28500
rect 57704 28552 57756 28558
rect 57704 28494 57756 28500
rect 57796 28552 57848 28558
rect 57796 28494 57848 28500
rect 58348 28552 58400 28558
rect 58348 28494 58400 28500
rect 57716 28218 57744 28494
rect 57704 28212 57756 28218
rect 57704 28154 57756 28160
rect 56784 28144 56836 28150
rect 56782 28112 56784 28121
rect 56836 28112 56838 28121
rect 56782 28047 56838 28056
rect 56784 27600 56836 27606
rect 56784 27542 56836 27548
rect 56796 25906 56824 27542
rect 56876 27532 56928 27538
rect 56876 27474 56928 27480
rect 56784 25900 56836 25906
rect 56784 25842 56836 25848
rect 56692 24404 56744 24410
rect 56692 24346 56744 24352
rect 56508 24200 56560 24206
rect 56508 24142 56560 24148
rect 56520 23848 56548 24142
rect 56520 23820 56732 23848
rect 56508 23724 56560 23730
rect 56508 23666 56560 23672
rect 56232 23656 56284 23662
rect 56232 23598 56284 23604
rect 56048 22976 56100 22982
rect 56048 22918 56100 22924
rect 55312 22772 55364 22778
rect 55312 22714 55364 22720
rect 55312 22636 55364 22642
rect 55312 22578 55364 22584
rect 55324 22234 55352 22578
rect 55312 22228 55364 22234
rect 55312 22170 55364 22176
rect 55128 22160 55180 22166
rect 55128 22102 55180 22108
rect 54944 22024 54996 22030
rect 54944 21966 54996 21972
rect 54760 21548 54812 21554
rect 54760 21490 54812 21496
rect 54772 21146 54800 21490
rect 54576 21140 54628 21146
rect 54576 21082 54628 21088
rect 54760 21140 54812 21146
rect 54760 21082 54812 21088
rect 55140 20890 55168 22102
rect 56244 22094 56272 23598
rect 56520 23322 56548 23666
rect 56600 23520 56652 23526
rect 56600 23462 56652 23468
rect 56508 23316 56560 23322
rect 56508 23258 56560 23264
rect 56612 22094 56640 23462
rect 56704 22438 56732 23820
rect 56796 23322 56824 25842
rect 56888 25770 56916 27474
rect 57716 27470 57744 28154
rect 57704 27464 57756 27470
rect 57704 27406 57756 27412
rect 57152 26988 57204 26994
rect 57152 26930 57204 26936
rect 56968 26784 57020 26790
rect 56968 26726 57020 26732
rect 56980 25838 57008 26726
rect 57060 26308 57112 26314
rect 57060 26250 57112 26256
rect 57072 26042 57100 26250
rect 57060 26036 57112 26042
rect 57060 25978 57112 25984
rect 56968 25832 57020 25838
rect 56968 25774 57020 25780
rect 56876 25764 56928 25770
rect 56876 25706 56928 25712
rect 57164 25294 57192 26930
rect 57152 25288 57204 25294
rect 57152 25230 57204 25236
rect 57808 25158 57836 28494
rect 58360 27674 58388 28494
rect 58820 28218 58848 37454
rect 58898 37360 58954 37369
rect 58898 37295 58900 37304
rect 58952 37295 58954 37304
rect 58900 37266 58952 37272
rect 58900 36644 58952 36650
rect 58900 36586 58952 36592
rect 58912 36553 58940 36586
rect 58898 36544 58954 36553
rect 58898 36479 58954 36488
rect 58900 36032 58952 36038
rect 58900 35974 58952 35980
rect 58912 35737 58940 35974
rect 58898 35728 58954 35737
rect 58898 35663 58954 35672
rect 58900 35012 58952 35018
rect 58900 34954 58952 34960
rect 58912 34921 58940 34954
rect 58898 34912 58954 34921
rect 58898 34847 58954 34856
rect 58900 34536 58952 34542
rect 58900 34478 58952 34484
rect 58912 34105 58940 34478
rect 58898 34096 58954 34105
rect 58898 34031 58954 34040
rect 58900 33380 58952 33386
rect 58900 33322 58952 33328
rect 58912 33289 58940 33322
rect 58898 33280 58954 33289
rect 58898 33215 58954 33224
rect 58900 32836 58952 32842
rect 58900 32778 58952 32784
rect 58912 32473 58940 32778
rect 58898 32464 58954 32473
rect 58898 32399 58954 32408
rect 58900 31816 58952 31822
rect 58900 31758 58952 31764
rect 58912 31657 58940 31758
rect 58898 31648 58954 31657
rect 58898 31583 58954 31592
rect 58898 28384 58954 28393
rect 58898 28319 58954 28328
rect 58808 28212 58860 28218
rect 58808 28154 58860 28160
rect 58348 27668 58400 27674
rect 58348 27610 58400 27616
rect 58714 27568 58770 27577
rect 58714 27503 58770 27512
rect 58728 27402 58756 27503
rect 58912 27470 58940 28319
rect 58900 27464 58952 27470
rect 58900 27406 58952 27412
rect 58716 27396 58768 27402
rect 58716 27338 58768 27344
rect 58164 27328 58216 27334
rect 58164 27270 58216 27276
rect 58176 27130 58204 27270
rect 58164 27124 58216 27130
rect 58164 27066 58216 27072
rect 58898 26752 58954 26761
rect 58898 26687 58954 26696
rect 58912 26382 58940 26687
rect 58900 26376 58952 26382
rect 58900 26318 58952 26324
rect 58256 26240 58308 26246
rect 58256 26182 58308 26188
rect 58268 26042 58296 26182
rect 58256 26036 58308 26042
rect 58256 25978 58308 25984
rect 57980 25968 58032 25974
rect 57980 25910 58032 25916
rect 58622 25936 58678 25945
rect 57992 25362 58020 25910
rect 58622 25871 58624 25880
rect 58676 25871 58678 25880
rect 58624 25842 58676 25848
rect 58072 25696 58124 25702
rect 58072 25638 58124 25644
rect 58084 25362 58112 25638
rect 57980 25356 58032 25362
rect 57980 25298 58032 25304
rect 58072 25356 58124 25362
rect 58072 25298 58124 25304
rect 57428 25152 57480 25158
rect 57428 25094 57480 25100
rect 57612 25152 57664 25158
rect 57612 25094 57664 25100
rect 57796 25152 57848 25158
rect 57796 25094 57848 25100
rect 57440 24954 57468 25094
rect 57428 24948 57480 24954
rect 57428 24890 57480 24896
rect 57060 24608 57112 24614
rect 57060 24550 57112 24556
rect 57072 24410 57100 24550
rect 57060 24404 57112 24410
rect 57060 24346 57112 24352
rect 57428 24200 57480 24206
rect 57428 24142 57480 24148
rect 56784 23316 56836 23322
rect 56784 23258 56836 23264
rect 57336 23112 57388 23118
rect 57336 23054 57388 23060
rect 57348 22778 57376 23054
rect 57440 22778 57468 24142
rect 57624 23118 57652 25094
rect 57992 24750 58020 25298
rect 58624 25220 58676 25226
rect 58624 25162 58676 25168
rect 58072 25152 58124 25158
rect 58636 25129 58664 25162
rect 58072 25094 58124 25100
rect 58622 25120 58678 25129
rect 58084 24954 58112 25094
rect 58622 25055 58678 25064
rect 58072 24948 58124 24954
rect 58072 24890 58124 24896
rect 57980 24744 58032 24750
rect 57980 24686 58032 24692
rect 57888 24608 57940 24614
rect 57888 24550 57940 24556
rect 58716 24608 58768 24614
rect 58716 24550 58768 24556
rect 57900 24410 57928 24550
rect 57888 24404 57940 24410
rect 57888 24346 57940 24352
rect 58728 24313 58756 24550
rect 58714 24304 58770 24313
rect 58714 24239 58770 24248
rect 58164 24200 58216 24206
rect 58164 24142 58216 24148
rect 57980 24064 58032 24070
rect 57980 24006 58032 24012
rect 57992 23866 58020 24006
rect 57980 23860 58032 23866
rect 57980 23802 58032 23808
rect 57888 23520 57940 23526
rect 57888 23462 57940 23468
rect 57900 23254 57928 23462
rect 57888 23248 57940 23254
rect 57888 23190 57940 23196
rect 57520 23112 57572 23118
rect 57520 23054 57572 23060
rect 57612 23112 57664 23118
rect 57612 23054 57664 23060
rect 57980 23112 58032 23118
rect 57980 23054 58032 23060
rect 57532 22778 57560 23054
rect 57336 22772 57388 22778
rect 57336 22714 57388 22720
rect 57428 22772 57480 22778
rect 57428 22714 57480 22720
rect 57520 22772 57572 22778
rect 57520 22714 57572 22720
rect 57428 22636 57480 22642
rect 57428 22578 57480 22584
rect 56692 22432 56744 22438
rect 56692 22374 56744 22380
rect 56968 22432 57020 22438
rect 56968 22374 57020 22380
rect 56980 22094 57008 22374
rect 57440 22234 57468 22578
rect 57428 22228 57480 22234
rect 57428 22170 57480 22176
rect 57624 22166 57652 23054
rect 57612 22160 57664 22166
rect 57612 22102 57664 22108
rect 56244 22066 56456 22094
rect 56612 22066 56732 22094
rect 55956 22024 56008 22030
rect 55956 21966 56008 21972
rect 55220 21956 55272 21962
rect 55220 21898 55272 21904
rect 55232 21350 55260 21898
rect 55968 21690 55996 21966
rect 55956 21684 56008 21690
rect 55956 21626 56008 21632
rect 56428 21486 56456 22066
rect 56416 21480 56468 21486
rect 56416 21422 56468 21428
rect 55220 21344 55272 21350
rect 55220 21286 55272 21292
rect 55404 21344 55456 21350
rect 55404 21286 55456 21292
rect 55048 20862 55168 20890
rect 54300 20256 54352 20262
rect 54300 20198 54352 20204
rect 54312 19854 54340 20198
rect 54024 19848 54076 19854
rect 53760 19808 54024 19836
rect 53656 19780 53708 19786
rect 53656 19722 53708 19728
rect 53472 19712 53524 19718
rect 53472 19654 53524 19660
rect 53380 17604 53432 17610
rect 53380 17546 53432 17552
rect 53196 16584 53248 16590
rect 53196 16526 53248 16532
rect 53288 16584 53340 16590
rect 53288 16526 53340 16532
rect 53104 15904 53156 15910
rect 53104 15846 53156 15852
rect 53116 15638 53144 15846
rect 53104 15632 53156 15638
rect 53104 15574 53156 15580
rect 53208 15162 53236 16526
rect 53300 16250 53328 16526
rect 53288 16244 53340 16250
rect 53288 16186 53340 16192
rect 53392 16182 53420 17546
rect 53484 16794 53512 19654
rect 53668 19514 53696 19722
rect 53656 19508 53708 19514
rect 53656 19450 53708 19456
rect 53656 19372 53708 19378
rect 53656 19314 53708 19320
rect 53668 18426 53696 19314
rect 53656 18420 53708 18426
rect 53656 18362 53708 18368
rect 53564 18284 53616 18290
rect 53564 18226 53616 18232
rect 53656 18284 53708 18290
rect 53760 18272 53788 19808
rect 54024 19790 54076 19796
rect 54208 19848 54260 19854
rect 54208 19790 54260 19796
rect 54300 19848 54352 19854
rect 54300 19790 54352 19796
rect 54220 19378 54248 19790
rect 55048 19786 55076 20862
rect 55128 20800 55180 20806
rect 55128 20742 55180 20748
rect 55036 19780 55088 19786
rect 55036 19722 55088 19728
rect 54208 19372 54260 19378
rect 54208 19314 54260 19320
rect 53840 19304 53892 19310
rect 53840 19246 53892 19252
rect 53852 18902 53880 19246
rect 55048 19174 55076 19722
rect 55140 19310 55168 20742
rect 55232 20058 55260 21286
rect 55416 21010 55444 21286
rect 55404 21004 55456 21010
rect 55404 20946 55456 20952
rect 56428 20942 56456 21422
rect 56600 21344 56652 21350
rect 56600 21286 56652 21292
rect 56612 21146 56640 21286
rect 56600 21140 56652 21146
rect 56600 21082 56652 21088
rect 55864 20936 55916 20942
rect 55864 20878 55916 20884
rect 55956 20936 56008 20942
rect 55956 20878 56008 20884
rect 56416 20936 56468 20942
rect 56416 20878 56468 20884
rect 55876 20602 55904 20878
rect 55968 20602 55996 20878
rect 55864 20596 55916 20602
rect 55864 20538 55916 20544
rect 55956 20596 56008 20602
rect 55956 20538 56008 20544
rect 56324 20460 56376 20466
rect 56324 20402 56376 20408
rect 55220 20052 55272 20058
rect 55220 19994 55272 20000
rect 55312 19848 55364 19854
rect 55312 19790 55364 19796
rect 55220 19780 55272 19786
rect 55220 19722 55272 19728
rect 55232 19514 55260 19722
rect 55220 19508 55272 19514
rect 55220 19450 55272 19456
rect 55128 19304 55180 19310
rect 55128 19246 55180 19252
rect 54852 19168 54904 19174
rect 54852 19110 54904 19116
rect 55036 19168 55088 19174
rect 55036 19110 55088 19116
rect 53840 18896 53892 18902
rect 53840 18838 53892 18844
rect 54760 18760 54812 18766
rect 54760 18702 54812 18708
rect 53932 18624 53984 18630
rect 53932 18566 53984 18572
rect 53944 18426 53972 18566
rect 54772 18426 54800 18702
rect 53932 18420 53984 18426
rect 53932 18362 53984 18368
rect 54760 18420 54812 18426
rect 54760 18362 54812 18368
rect 53840 18352 53892 18358
rect 53892 18300 54064 18306
rect 53840 18294 54064 18300
rect 53852 18278 54064 18294
rect 53708 18244 53788 18272
rect 53656 18226 53708 18232
rect 53576 18154 53604 18226
rect 53564 18148 53616 18154
rect 53564 18090 53616 18096
rect 53576 17882 53604 18090
rect 53564 17876 53616 17882
rect 53564 17818 53616 17824
rect 53472 16788 53524 16794
rect 53472 16730 53524 16736
rect 53564 16720 53616 16726
rect 53484 16668 53564 16674
rect 53484 16662 53616 16668
rect 53484 16646 53604 16662
rect 53380 16176 53432 16182
rect 53380 16118 53432 16124
rect 53392 15978 53420 16118
rect 53380 15972 53432 15978
rect 53380 15914 53432 15920
rect 51632 15156 51684 15162
rect 51632 15098 51684 15104
rect 52828 15156 52880 15162
rect 52828 15098 52880 15104
rect 53012 15156 53064 15162
rect 53012 15098 53064 15104
rect 53196 15156 53248 15162
rect 53196 15098 53248 15104
rect 53392 15094 53420 15914
rect 53484 15706 53512 16646
rect 53564 16584 53616 16590
rect 53564 16526 53616 16532
rect 53576 16250 53604 16526
rect 53668 16454 53696 18226
rect 53840 18216 53892 18222
rect 53840 18158 53892 18164
rect 53748 18080 53800 18086
rect 53748 18022 53800 18028
rect 53760 17678 53788 18022
rect 53852 17882 53880 18158
rect 53840 17876 53892 17882
rect 53840 17818 53892 17824
rect 53748 17672 53800 17678
rect 53748 17614 53800 17620
rect 53932 17672 53984 17678
rect 53932 17614 53984 17620
rect 53656 16448 53708 16454
rect 53656 16390 53708 16396
rect 53564 16244 53616 16250
rect 53564 16186 53616 16192
rect 53668 16182 53696 16390
rect 53656 16176 53708 16182
rect 53656 16118 53708 16124
rect 53472 15700 53524 15706
rect 53472 15642 53524 15648
rect 53484 15502 53512 15642
rect 53472 15496 53524 15502
rect 53472 15438 53524 15444
rect 53564 15496 53616 15502
rect 53564 15438 53616 15444
rect 53576 15162 53604 15438
rect 53668 15162 53696 16118
rect 53944 15706 53972 17614
rect 54036 15978 54064 18278
rect 54864 17882 54892 19110
rect 55220 18080 55272 18086
rect 55220 18022 55272 18028
rect 55232 17882 55260 18022
rect 54852 17876 54904 17882
rect 54852 17818 54904 17824
rect 55220 17876 55272 17882
rect 55220 17818 55272 17824
rect 54116 16448 54168 16454
rect 54116 16390 54168 16396
rect 54128 16250 54156 16390
rect 54116 16244 54168 16250
rect 54116 16186 54168 16192
rect 54024 15972 54076 15978
rect 54076 15932 54156 15960
rect 54024 15914 54076 15920
rect 53932 15700 53984 15706
rect 53932 15642 53984 15648
rect 54024 15428 54076 15434
rect 54024 15370 54076 15376
rect 54036 15162 54064 15370
rect 53564 15156 53616 15162
rect 53564 15098 53616 15104
rect 53656 15156 53708 15162
rect 53656 15098 53708 15104
rect 54024 15156 54076 15162
rect 54024 15098 54076 15104
rect 53380 15088 53432 15094
rect 53380 15030 53432 15036
rect 51448 15020 51500 15026
rect 51448 14962 51500 14968
rect 52736 15020 52788 15026
rect 52736 14962 52788 14968
rect 52920 15020 52972 15026
rect 52920 14962 52972 14968
rect 51460 14074 51488 14962
rect 52748 14618 52776 14962
rect 52736 14612 52788 14618
rect 52736 14554 52788 14560
rect 52276 14408 52328 14414
rect 52276 14350 52328 14356
rect 52092 14272 52144 14278
rect 52092 14214 52144 14220
rect 51448 14068 51500 14074
rect 51448 14010 51500 14016
rect 51264 13932 51316 13938
rect 51448 13932 51500 13938
rect 51316 13892 51448 13920
rect 51264 13874 51316 13880
rect 51448 13874 51500 13880
rect 51540 13932 51592 13938
rect 51540 13874 51592 13880
rect 51816 13932 51868 13938
rect 51816 13874 51868 13880
rect 51552 13530 51580 13874
rect 51540 13524 51592 13530
rect 51540 13466 51592 13472
rect 51448 13320 51500 13326
rect 51448 13262 51500 13268
rect 51460 12986 51488 13262
rect 51828 12986 51856 13874
rect 52104 13326 52132 14214
rect 52092 13320 52144 13326
rect 52092 13262 52144 13268
rect 52184 13320 52236 13326
rect 52184 13262 52236 13268
rect 51448 12980 51500 12986
rect 51448 12922 51500 12928
rect 51816 12980 51868 12986
rect 51816 12922 51868 12928
rect 51632 12912 51684 12918
rect 51632 12854 51684 12860
rect 51172 12844 51224 12850
rect 51172 12786 51224 12792
rect 51540 12776 51592 12782
rect 51078 12744 51134 12753
rect 51540 12718 51592 12724
rect 51078 12679 51080 12688
rect 51132 12679 51134 12688
rect 51080 12650 51132 12656
rect 51552 12442 51580 12718
rect 51540 12436 51592 12442
rect 51540 12378 51592 12384
rect 50988 12232 51040 12238
rect 50988 12174 51040 12180
rect 50528 12164 50580 12170
rect 50528 12106 50580 12112
rect 51644 12102 51672 12854
rect 52092 12436 52144 12442
rect 52196 12434 52224 13262
rect 52288 12986 52316 14350
rect 52932 14074 52960 14962
rect 53392 14414 53420 15030
rect 53380 14408 53432 14414
rect 53380 14350 53432 14356
rect 52920 14068 52972 14074
rect 52920 14010 52972 14016
rect 53012 14068 53064 14074
rect 53012 14010 53064 14016
rect 52920 13864 52972 13870
rect 53024 13852 53052 14010
rect 53104 13932 53156 13938
rect 53104 13874 53156 13880
rect 52972 13824 53052 13852
rect 52920 13806 52972 13812
rect 52644 13184 52696 13190
rect 52644 13126 52696 13132
rect 52920 13184 52972 13190
rect 53116 13172 53144 13874
rect 53392 13326 53420 14350
rect 53668 14074 53696 15098
rect 54128 15094 54156 15932
rect 54864 15570 54892 17818
rect 55128 17740 55180 17746
rect 55128 17682 55180 17688
rect 55140 17338 55168 17682
rect 55324 17678 55352 19790
rect 56336 19718 56364 20402
rect 56428 19854 56456 20878
rect 56704 20482 56732 22066
rect 56980 22066 57100 22094
rect 56876 22024 56928 22030
rect 56980 21978 57008 22066
rect 56928 21972 57008 21978
rect 56876 21966 57008 21972
rect 56784 21956 56836 21962
rect 56888 21950 57008 21966
rect 57072 21962 57100 22066
rect 57428 22092 57480 22098
rect 57428 22034 57480 22040
rect 57152 22024 57204 22030
rect 57152 21966 57204 21972
rect 57060 21956 57112 21962
rect 56784 21898 56836 21904
rect 57060 21898 57112 21904
rect 56796 21690 56824 21898
rect 56784 21684 56836 21690
rect 56784 21626 56836 21632
rect 57164 20534 57192 21966
rect 57440 21146 57468 22034
rect 57888 21956 57940 21962
rect 57888 21898 57940 21904
rect 57900 21690 57928 21898
rect 57992 21894 58020 23054
rect 58176 22778 58204 24142
rect 58898 23488 58954 23497
rect 58898 23423 58954 23432
rect 58256 23112 58308 23118
rect 58256 23054 58308 23060
rect 58268 22778 58296 23054
rect 58912 22778 58940 23423
rect 58164 22772 58216 22778
rect 58164 22714 58216 22720
rect 58256 22772 58308 22778
rect 58256 22714 58308 22720
rect 58900 22772 58952 22778
rect 58900 22714 58952 22720
rect 58806 22672 58862 22681
rect 58806 22607 58808 22616
rect 58860 22607 58862 22616
rect 58808 22578 58860 22584
rect 58900 21956 58952 21962
rect 58900 21898 58952 21904
rect 57980 21888 58032 21894
rect 57980 21830 58032 21836
rect 58072 21888 58124 21894
rect 58072 21830 58124 21836
rect 58256 21888 58308 21894
rect 58256 21830 58308 21836
rect 58348 21888 58400 21894
rect 58348 21830 58400 21836
rect 58716 21888 58768 21894
rect 58912 21865 58940 21898
rect 58716 21830 58768 21836
rect 58898 21856 58954 21865
rect 57888 21684 57940 21690
rect 57888 21626 57940 21632
rect 57888 21480 57940 21486
rect 57888 21422 57940 21428
rect 57900 21146 57928 21422
rect 57428 21140 57480 21146
rect 57428 21082 57480 21088
rect 57888 21140 57940 21146
rect 57888 21082 57940 21088
rect 57992 20942 58020 21830
rect 58084 21690 58112 21830
rect 58072 21684 58124 21690
rect 58072 21626 58124 21632
rect 57980 20936 58032 20942
rect 57980 20878 58032 20884
rect 57152 20528 57204 20534
rect 56704 20454 56824 20482
rect 57152 20470 57204 20476
rect 56692 20392 56744 20398
rect 56692 20334 56744 20340
rect 56704 20058 56732 20334
rect 56692 20052 56744 20058
rect 56692 19994 56744 20000
rect 56416 19848 56468 19854
rect 56416 19790 56468 19796
rect 55680 19712 55732 19718
rect 55680 19654 55732 19660
rect 56324 19712 56376 19718
rect 56324 19654 56376 19660
rect 55692 19378 55720 19654
rect 56138 19408 56194 19417
rect 55680 19372 55732 19378
rect 56138 19343 56140 19352
rect 55680 19314 55732 19320
rect 56192 19343 56194 19352
rect 56140 19314 56192 19320
rect 56336 18766 56364 19654
rect 56600 19440 56652 19446
rect 56600 19382 56652 19388
rect 55404 18760 55456 18766
rect 55404 18702 55456 18708
rect 56324 18760 56376 18766
rect 56324 18702 56376 18708
rect 55312 17672 55364 17678
rect 55312 17614 55364 17620
rect 55128 17332 55180 17338
rect 55128 17274 55180 17280
rect 55324 15910 55352 17614
rect 55416 17270 55444 18702
rect 56612 18426 56640 19382
rect 56796 18902 56824 20454
rect 57796 20256 57848 20262
rect 57796 20198 57848 20204
rect 57060 19780 57112 19786
rect 57060 19722 57112 19728
rect 57072 19514 57100 19722
rect 57336 19712 57388 19718
rect 57336 19654 57388 19660
rect 57060 19508 57112 19514
rect 57060 19450 57112 19456
rect 57348 19378 57376 19654
rect 57612 19508 57664 19514
rect 57612 19450 57664 19456
rect 57624 19417 57652 19450
rect 57610 19408 57666 19417
rect 57336 19372 57388 19378
rect 57808 19378 57836 20198
rect 58268 19854 58296 21830
rect 58360 20942 58388 21830
rect 58728 21049 58756 21830
rect 58898 21791 58954 21800
rect 58714 21040 58770 21049
rect 58714 20975 58770 20984
rect 58348 20936 58400 20942
rect 58348 20878 58400 20884
rect 58532 20256 58584 20262
rect 58530 20224 58532 20233
rect 58584 20224 58586 20233
rect 58530 20159 58586 20168
rect 58256 19848 58308 19854
rect 58256 19790 58308 19796
rect 58348 19508 58400 19514
rect 58348 19450 58400 19456
rect 57610 19343 57666 19352
rect 57796 19372 57848 19378
rect 57336 19314 57388 19320
rect 57796 19314 57848 19320
rect 57060 19304 57112 19310
rect 57428 19304 57480 19310
rect 57112 19252 57428 19258
rect 57060 19246 57480 19252
rect 57072 19230 57468 19246
rect 57612 19236 57664 19242
rect 57612 19178 57664 19184
rect 57336 19168 57388 19174
rect 57336 19110 57388 19116
rect 56784 18896 56836 18902
rect 56784 18838 56836 18844
rect 57348 18834 57376 19110
rect 57624 18970 57652 19178
rect 57612 18964 57664 18970
rect 57612 18906 57664 18912
rect 57336 18828 57388 18834
rect 57336 18770 57388 18776
rect 56600 18420 56652 18426
rect 56600 18362 56652 18368
rect 56968 18284 57020 18290
rect 56968 18226 57020 18232
rect 56508 17536 56560 17542
rect 56508 17478 56560 17484
rect 55404 17264 55456 17270
rect 55404 17206 55456 17212
rect 56520 17202 56548 17478
rect 56980 17338 57008 18226
rect 56968 17332 57020 17338
rect 56968 17274 57020 17280
rect 57348 17202 57376 18770
rect 57808 18766 57836 19314
rect 58360 18970 58388 19450
rect 58898 19408 58954 19417
rect 58898 19343 58954 19352
rect 58348 18964 58400 18970
rect 58348 18906 58400 18912
rect 58164 18896 58216 18902
rect 58164 18838 58216 18844
rect 58254 18864 58310 18873
rect 57796 18760 57848 18766
rect 58072 18760 58124 18766
rect 57796 18702 57848 18708
rect 57900 18720 58072 18748
rect 57900 18630 57928 18720
rect 58072 18702 58124 18708
rect 57888 18624 57940 18630
rect 57888 18566 57940 18572
rect 57980 18624 58032 18630
rect 57980 18566 58032 18572
rect 58072 18624 58124 18630
rect 58072 18566 58124 18572
rect 57796 18216 57848 18222
rect 57796 18158 57848 18164
rect 57612 18148 57664 18154
rect 57612 18090 57664 18096
rect 57624 17678 57652 18090
rect 57808 17785 57836 18158
rect 57900 17882 57928 18566
rect 57992 18426 58020 18566
rect 58084 18426 58112 18566
rect 57980 18420 58032 18426
rect 57980 18362 58032 18368
rect 58072 18420 58124 18426
rect 58072 18362 58124 18368
rect 57888 17876 57940 17882
rect 57888 17818 57940 17824
rect 57980 17876 58032 17882
rect 57980 17818 58032 17824
rect 57794 17776 57850 17785
rect 57794 17711 57850 17720
rect 57612 17672 57664 17678
rect 57900 17626 57928 17818
rect 57992 17660 58020 17818
rect 58072 17672 58124 17678
rect 57992 17632 58072 17660
rect 57612 17614 57664 17620
rect 57624 17202 57652 17614
rect 57704 17604 57756 17610
rect 57704 17546 57756 17552
rect 57808 17598 57928 17626
rect 58072 17614 58124 17620
rect 57716 17338 57744 17546
rect 57704 17332 57756 17338
rect 57704 17274 57756 17280
rect 56508 17196 56560 17202
rect 56508 17138 56560 17144
rect 57336 17196 57388 17202
rect 57336 17138 57388 17144
rect 57612 17196 57664 17202
rect 57612 17138 57664 17144
rect 56876 16720 56928 16726
rect 56876 16662 56928 16668
rect 55588 16584 55640 16590
rect 55588 16526 55640 16532
rect 56600 16584 56652 16590
rect 56600 16526 56652 16532
rect 55496 16448 55548 16454
rect 55496 16390 55548 16396
rect 55404 16108 55456 16114
rect 55404 16050 55456 16056
rect 55312 15904 55364 15910
rect 55312 15846 55364 15852
rect 54852 15564 54904 15570
rect 54852 15506 54904 15512
rect 54116 15088 54168 15094
rect 54116 15030 54168 15036
rect 53932 15020 53984 15026
rect 53932 14962 53984 14968
rect 53840 14952 53892 14958
rect 53840 14894 53892 14900
rect 53852 14074 53880 14894
rect 53944 14414 53972 14962
rect 54024 14884 54076 14890
rect 54024 14826 54076 14832
rect 53932 14408 53984 14414
rect 53932 14350 53984 14356
rect 54036 14278 54064 14826
rect 54024 14272 54076 14278
rect 54024 14214 54076 14220
rect 53656 14068 53708 14074
rect 53656 14010 53708 14016
rect 53840 14068 53892 14074
rect 54128 14056 54156 15030
rect 54760 14272 54812 14278
rect 54760 14214 54812 14220
rect 53840 14010 53892 14016
rect 53944 14028 54156 14056
rect 53944 13938 53972 14028
rect 53932 13932 53984 13938
rect 53932 13874 53984 13880
rect 54024 13932 54076 13938
rect 54024 13874 54076 13880
rect 53840 13728 53892 13734
rect 53840 13670 53892 13676
rect 53852 13530 53880 13670
rect 54036 13530 54064 13874
rect 54772 13802 54800 14214
rect 54760 13796 54812 13802
rect 54760 13738 54812 13744
rect 53840 13524 53892 13530
rect 53840 13466 53892 13472
rect 54024 13524 54076 13530
rect 54024 13466 54076 13472
rect 53380 13320 53432 13326
rect 53380 13262 53432 13268
rect 53564 13320 53616 13326
rect 53564 13262 53616 13268
rect 53932 13320 53984 13326
rect 53932 13262 53984 13268
rect 52972 13144 53144 13172
rect 52920 13126 52972 13132
rect 52276 12980 52328 12986
rect 52328 12940 52408 12968
rect 52276 12922 52328 12928
rect 52144 12406 52224 12434
rect 52092 12378 52144 12384
rect 52092 12232 52144 12238
rect 52092 12174 52144 12180
rect 52104 12102 52132 12174
rect 51632 12096 51684 12102
rect 51632 12038 51684 12044
rect 52092 12096 52144 12102
rect 52092 12038 52144 12044
rect 50294 11996 50602 12005
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11931 50602 11940
rect 49884 11892 49936 11898
rect 49884 11834 49936 11840
rect 52380 11694 52408 12940
rect 52656 12782 52684 13126
rect 52644 12776 52696 12782
rect 52644 12718 52696 12724
rect 52736 12776 52788 12782
rect 52736 12718 52788 12724
rect 52748 12306 52776 12718
rect 52736 12300 52788 12306
rect 52736 12242 52788 12248
rect 52932 12238 52960 13126
rect 53576 12986 53604 13262
rect 53564 12980 53616 12986
rect 53564 12922 53616 12928
rect 53944 12850 53972 13262
rect 54208 13252 54260 13258
rect 54208 13194 54260 13200
rect 54220 12986 54248 13194
rect 54208 12980 54260 12986
rect 54208 12922 54260 12928
rect 54772 12850 54800 13738
rect 54864 13734 54892 15506
rect 55324 14414 55352 15846
rect 55416 15706 55444 16050
rect 55404 15700 55456 15706
rect 55404 15642 55456 15648
rect 55508 15570 55536 16390
rect 55600 16250 55628 16526
rect 56612 16250 56640 16526
rect 56888 16522 56916 16662
rect 56876 16516 56928 16522
rect 56876 16458 56928 16464
rect 56784 16448 56836 16454
rect 56784 16390 56836 16396
rect 55588 16244 55640 16250
rect 55588 16186 55640 16192
rect 56600 16244 56652 16250
rect 56600 16186 56652 16192
rect 56796 16182 56824 16390
rect 56888 16182 56916 16458
rect 57348 16250 57376 17138
rect 57808 16794 57836 17598
rect 57900 17462 58020 17490
rect 57796 16788 57848 16794
rect 57796 16730 57848 16736
rect 57336 16244 57388 16250
rect 57336 16186 57388 16192
rect 56784 16176 56836 16182
rect 56784 16118 56836 16124
rect 56876 16176 56928 16182
rect 56876 16118 56928 16124
rect 56600 15904 56652 15910
rect 56600 15846 56652 15852
rect 56612 15706 56640 15846
rect 56600 15700 56652 15706
rect 56600 15642 56652 15648
rect 56796 15638 56824 16118
rect 56888 15638 56916 16118
rect 57808 16114 57836 16730
rect 57796 16108 57848 16114
rect 57796 16050 57848 16056
rect 57152 16040 57204 16046
rect 57152 15982 57204 15988
rect 57704 16040 57756 16046
rect 57704 15982 57756 15988
rect 57164 15706 57192 15982
rect 57716 15706 57744 15982
rect 57152 15700 57204 15706
rect 57152 15642 57204 15648
rect 57704 15700 57756 15706
rect 57704 15642 57756 15648
rect 57808 15638 57836 16050
rect 57900 15978 57928 17462
rect 57992 17338 58020 17462
rect 57980 17332 58032 17338
rect 57980 17274 58032 17280
rect 58176 17066 58204 18838
rect 58254 18799 58310 18808
rect 58268 17882 58296 18799
rect 58912 18766 58940 19343
rect 58348 18760 58400 18766
rect 58348 18702 58400 18708
rect 58900 18760 58952 18766
rect 58900 18702 58952 18708
rect 58360 18426 58388 18702
rect 58898 18592 58954 18601
rect 58898 18527 58954 18536
rect 58912 18426 58940 18527
rect 58348 18420 58400 18426
rect 58348 18362 58400 18368
rect 58900 18420 58952 18426
rect 58900 18362 58952 18368
rect 58348 18080 58400 18086
rect 58348 18022 58400 18028
rect 58256 17876 58308 17882
rect 58256 17818 58308 17824
rect 58256 17672 58308 17678
rect 58256 17614 58308 17620
rect 58268 17338 58296 17614
rect 58256 17332 58308 17338
rect 58256 17274 58308 17280
rect 58360 17202 58388 18022
rect 58348 17196 58400 17202
rect 58348 17138 58400 17144
rect 58164 17060 58216 17066
rect 58164 17002 58216 17008
rect 58900 17060 58952 17066
rect 58900 17002 58952 17008
rect 57980 16992 58032 16998
rect 58912 16969 58940 17002
rect 57980 16934 58032 16940
rect 58898 16960 58954 16969
rect 57992 16794 58020 16934
rect 58898 16895 58954 16904
rect 57980 16788 58032 16794
rect 57980 16730 58032 16736
rect 58164 16584 58216 16590
rect 58164 16526 58216 16532
rect 57980 16448 58032 16454
rect 57980 16390 58032 16396
rect 57888 15972 57940 15978
rect 57888 15914 57940 15920
rect 57992 15706 58020 16390
rect 58176 15706 58204 16526
rect 58900 16448 58952 16454
rect 58900 16390 58952 16396
rect 58532 16176 58584 16182
rect 58912 16153 58940 16390
rect 58532 16118 58584 16124
rect 58898 16144 58954 16153
rect 58348 16108 58400 16114
rect 58348 16050 58400 16056
rect 57980 15700 58032 15706
rect 57980 15642 58032 15648
rect 58164 15700 58216 15706
rect 58164 15642 58216 15648
rect 56508 15632 56560 15638
rect 56784 15632 56836 15638
rect 56560 15580 56640 15586
rect 56508 15574 56640 15580
rect 56784 15574 56836 15580
rect 56876 15632 56928 15638
rect 57796 15632 57848 15638
rect 56876 15574 56928 15580
rect 57624 15580 57796 15586
rect 57624 15574 57848 15580
rect 55496 15564 55548 15570
rect 56520 15558 56640 15574
rect 55496 15506 55548 15512
rect 56324 15360 56376 15366
rect 56324 15302 56376 15308
rect 55588 15020 55640 15026
rect 55588 14962 55640 14968
rect 55496 14816 55548 14822
rect 55496 14758 55548 14764
rect 55312 14408 55364 14414
rect 55312 14350 55364 14356
rect 55220 14340 55272 14346
rect 55220 14282 55272 14288
rect 55036 14272 55088 14278
rect 55036 14214 55088 14220
rect 55048 14074 55076 14214
rect 55232 14074 55260 14282
rect 55036 14068 55088 14074
rect 55036 14010 55088 14016
rect 55220 14068 55272 14074
rect 55220 14010 55272 14016
rect 54852 13728 54904 13734
rect 54852 13670 54904 13676
rect 54864 13530 54892 13670
rect 54852 13524 54904 13530
rect 54852 13466 54904 13472
rect 53840 12844 53892 12850
rect 53840 12786 53892 12792
rect 53932 12844 53984 12850
rect 53932 12786 53984 12792
rect 54760 12844 54812 12850
rect 54760 12786 54812 12792
rect 53852 12238 53880 12786
rect 54482 12744 54538 12753
rect 54864 12714 54892 13466
rect 55324 12918 55352 14350
rect 55508 14074 55536 14758
rect 55600 14074 55628 14962
rect 56140 14952 56192 14958
rect 56140 14894 56192 14900
rect 56152 14074 56180 14894
rect 55496 14068 55548 14074
rect 55496 14010 55548 14016
rect 55588 14068 55640 14074
rect 55588 14010 55640 14016
rect 56140 14068 56192 14074
rect 56140 14010 56192 14016
rect 56336 13870 56364 15302
rect 56612 13954 56640 15558
rect 57624 15558 57836 15574
rect 56968 15360 57020 15366
rect 56968 15302 57020 15308
rect 57520 15360 57572 15366
rect 57624 15348 57652 15558
rect 57704 15496 57756 15502
rect 57704 15438 57756 15444
rect 58072 15496 58124 15502
rect 58072 15438 58124 15444
rect 57716 15366 57744 15438
rect 57572 15320 57652 15348
rect 57704 15360 57756 15366
rect 57520 15302 57572 15308
rect 57704 15302 57756 15308
rect 56980 15162 57008 15302
rect 57716 15162 57744 15302
rect 56968 15156 57020 15162
rect 56968 15098 57020 15104
rect 57704 15156 57756 15162
rect 57704 15098 57756 15104
rect 57152 14952 57204 14958
rect 57152 14894 57204 14900
rect 57164 14618 57192 14894
rect 57888 14816 57940 14822
rect 57888 14758 57940 14764
rect 57152 14612 57204 14618
rect 57152 14554 57204 14560
rect 56692 14544 56744 14550
rect 56692 14486 56744 14492
rect 56704 14074 56732 14486
rect 56784 14340 56836 14346
rect 56784 14282 56836 14288
rect 56796 14074 56824 14282
rect 56692 14068 56744 14074
rect 56692 14010 56744 14016
rect 56784 14068 56836 14074
rect 56784 14010 56836 14016
rect 56612 13926 56732 13954
rect 56324 13864 56376 13870
rect 56324 13806 56376 13812
rect 56048 13456 56100 13462
rect 56048 13398 56100 13404
rect 55956 13320 56008 13326
rect 55956 13262 56008 13268
rect 55312 12912 55364 12918
rect 55312 12854 55364 12860
rect 54482 12679 54538 12688
rect 54852 12708 54904 12714
rect 54496 12646 54524 12679
rect 54852 12650 54904 12656
rect 54392 12640 54444 12646
rect 54392 12582 54444 12588
rect 54484 12640 54536 12646
rect 54484 12582 54536 12588
rect 54404 12238 54432 12582
rect 55968 12442 55996 13262
rect 55956 12436 56008 12442
rect 55956 12378 56008 12384
rect 56060 12374 56088 13398
rect 56140 12776 56192 12782
rect 56140 12718 56192 12724
rect 56152 12442 56180 12718
rect 56140 12436 56192 12442
rect 56140 12378 56192 12384
rect 56048 12368 56100 12374
rect 56048 12310 56100 12316
rect 56336 12238 56364 13806
rect 56600 13728 56652 13734
rect 56600 13670 56652 13676
rect 56612 13530 56640 13670
rect 56600 13524 56652 13530
rect 56600 13466 56652 13472
rect 56600 13388 56652 13394
rect 56600 13330 56652 13336
rect 56508 13184 56560 13190
rect 56508 13126 56560 13132
rect 56520 12918 56548 13126
rect 56508 12912 56560 12918
rect 56508 12854 56560 12860
rect 56612 12442 56640 13330
rect 56704 13190 56732 13926
rect 57900 13870 57928 14758
rect 58084 14550 58112 15438
rect 58072 14544 58124 14550
rect 58072 14486 58124 14492
rect 58084 14074 58112 14486
rect 58164 14272 58216 14278
rect 58164 14214 58216 14220
rect 58176 14074 58204 14214
rect 58072 14068 58124 14074
rect 58072 14010 58124 14016
rect 58164 14068 58216 14074
rect 58164 14010 58216 14016
rect 57888 13864 57940 13870
rect 57888 13806 57940 13812
rect 57980 13796 58032 13802
rect 57980 13738 58032 13744
rect 56692 13184 56744 13190
rect 56692 13126 56744 13132
rect 56600 12436 56652 12442
rect 57992 12434 58020 13738
rect 58360 13530 58388 16050
rect 58440 15428 58492 15434
rect 58440 15370 58492 15376
rect 58452 15026 58480 15370
rect 58440 15020 58492 15026
rect 58440 14962 58492 14968
rect 58348 13524 58400 13530
rect 58348 13466 58400 13472
rect 58544 12986 58572 16118
rect 58898 16079 58954 16088
rect 58898 15328 58954 15337
rect 58898 15263 58954 15272
rect 58912 14618 58940 15263
rect 58900 14612 58952 14618
rect 58900 14554 58952 14560
rect 58898 14512 58954 14521
rect 58898 14447 58954 14456
rect 58912 14074 58940 14447
rect 58900 14068 58952 14074
rect 58900 14010 58952 14016
rect 58898 13696 58954 13705
rect 58898 13631 58954 13640
rect 58912 13326 58940 13631
rect 58900 13320 58952 13326
rect 58900 13262 58952 13268
rect 58716 13184 58768 13190
rect 58716 13126 58768 13132
rect 58532 12980 58584 12986
rect 58176 12940 58532 12968
rect 58072 12844 58124 12850
rect 58072 12786 58124 12792
rect 56600 12378 56652 12384
rect 57900 12406 58020 12434
rect 52920 12232 52972 12238
rect 52920 12174 52972 12180
rect 53840 12232 53892 12238
rect 53840 12174 53892 12180
rect 54392 12232 54444 12238
rect 54392 12174 54444 12180
rect 56324 12232 56376 12238
rect 56324 12174 56376 12180
rect 57900 11914 57928 12406
rect 57980 12164 58032 12170
rect 57980 12106 58032 12112
rect 57992 12073 58020 12106
rect 57978 12064 58034 12073
rect 57978 11999 58034 12008
rect 57900 11886 58020 11914
rect 52368 11688 52420 11694
rect 52368 11630 52420 11636
rect 50294 10908 50602 10917
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10843 50602 10852
rect 57992 10266 58020 11886
rect 57980 10260 58032 10266
rect 57980 10202 58032 10208
rect 50294 9820 50602 9829
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9755 50602 9764
rect 50294 8732 50602 8741
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8667 50602 8676
rect 58084 8634 58112 12786
rect 58176 12434 58204 12940
rect 58532 12922 58584 12928
rect 58728 12889 58756 13126
rect 58714 12880 58770 12889
rect 58714 12815 58770 12824
rect 58348 12708 58400 12714
rect 58348 12650 58400 12656
rect 58176 12406 58296 12434
rect 58268 12238 58296 12406
rect 58256 12232 58308 12238
rect 58256 12174 58308 12180
rect 58360 9178 58388 12650
rect 58624 11552 58676 11558
rect 58624 11494 58676 11500
rect 58636 11257 58664 11494
rect 58622 11248 58678 11257
rect 58622 11183 58678 11192
rect 58900 10532 58952 10538
rect 58900 10474 58952 10480
rect 58912 10441 58940 10474
rect 58898 10432 58954 10441
rect 58898 10367 58954 10376
rect 58900 9716 58952 9722
rect 58900 9658 58952 9664
rect 58912 9625 58940 9658
rect 58898 9616 58954 9625
rect 58898 9551 58954 9560
rect 58348 9172 58400 9178
rect 58348 9114 58400 9120
rect 58900 8900 58952 8906
rect 58900 8842 58952 8848
rect 58912 8809 58940 8842
rect 58898 8800 58954 8809
rect 58898 8735 58954 8744
rect 58072 8628 58124 8634
rect 58072 8570 58124 8576
rect 58900 8356 58952 8362
rect 58900 8298 58952 8304
rect 58912 7993 58940 8298
rect 58898 7984 58954 7993
rect 58898 7919 58954 7928
rect 50294 7644 50602 7653
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7579 50602 7588
rect 58900 7268 58952 7274
rect 58900 7210 58952 7216
rect 58912 7177 58940 7210
rect 58898 7168 58954 7177
rect 58898 7103 58954 7112
rect 50294 6556 50602 6565
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6491 50602 6500
rect 50294 5468 50602 5477
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5403 50602 5412
rect 50294 4380 50602 4389
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4315 50602 4324
rect 50294 3292 50602 3301
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3227 50602 3236
rect 49792 2644 49844 2650
rect 49792 2586 49844 2592
rect 47596 2514 47716 2530
rect 47596 2508 47728 2514
rect 47596 2502 47676 2508
rect 42432 2440 42484 2446
rect 42432 2382 42484 2388
rect 47216 2440 47268 2446
rect 47216 2382 47268 2388
rect 42248 2032 42300 2038
rect 42248 1974 42300 1980
rect 42444 1306 42472 2382
rect 42352 1278 42472 1306
rect 42352 800 42380 1278
rect 47320 870 47440 898
rect 47320 800 47348 870
rect 2594 0 2650 800
rect 7562 0 7618 800
rect 12530 0 12586 800
rect 17498 0 17554 800
rect 22466 0 22522 800
rect 27434 0 27490 800
rect 32402 0 32458 800
rect 37370 0 37426 800
rect 42338 0 42394 800
rect 47306 0 47362 800
rect 47412 762 47440 870
rect 47596 762 47624 2502
rect 47676 2450 47728 2456
rect 52460 2440 52512 2446
rect 52460 2382 52512 2388
rect 50294 2204 50602 2213
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2139 50602 2148
rect 52472 1442 52500 2382
rect 57244 2372 57296 2378
rect 57244 2314 57296 2320
rect 52288 1414 52500 1442
rect 52288 800 52316 1414
rect 57256 800 57284 2314
rect 47412 734 47624 762
rect 52274 0 52330 800
rect 57242 0 57298 800
<< via2 >>
rect 938 56888 994 56944
rect 938 55256 994 55312
rect 1582 53760 1638 53816
rect 1582 52436 1584 52456
rect 1584 52436 1636 52456
rect 1636 52436 1638 52456
rect 1582 52400 1638 52436
rect 938 50360 994 50416
rect 938 48728 994 48784
rect 938 47096 994 47152
rect 1582 45464 1638 45520
rect 1582 44104 1638 44160
rect 938 42200 994 42256
rect 1214 40568 1270 40624
rect 938 38956 994 38992
rect 938 38936 940 38956
rect 940 38936 992 38956
rect 992 38936 994 38956
rect 1582 37304 1638 37360
rect 938 35692 994 35728
rect 938 35672 940 35692
rect 940 35672 992 35692
rect 992 35672 994 35692
rect 938 34060 994 34096
rect 938 34040 940 34060
rect 940 34040 992 34060
rect 992 34040 994 34060
rect 938 32408 994 32464
rect 938 30776 994 30832
rect 938 29144 994 29200
rect 4220 57146 4276 57148
rect 4300 57146 4356 57148
rect 4380 57146 4436 57148
rect 4460 57146 4516 57148
rect 4220 57094 4266 57146
rect 4266 57094 4276 57146
rect 4300 57094 4330 57146
rect 4330 57094 4342 57146
rect 4342 57094 4356 57146
rect 4380 57094 4394 57146
rect 4394 57094 4406 57146
rect 4406 57094 4436 57146
rect 4460 57094 4470 57146
rect 4470 57094 4516 57146
rect 4220 57092 4276 57094
rect 4300 57092 4356 57094
rect 4380 57092 4436 57094
rect 4460 57092 4516 57094
rect 4220 56058 4276 56060
rect 4300 56058 4356 56060
rect 4380 56058 4436 56060
rect 4460 56058 4516 56060
rect 4220 56006 4266 56058
rect 4266 56006 4276 56058
rect 4300 56006 4330 56058
rect 4330 56006 4342 56058
rect 4342 56006 4356 56058
rect 4380 56006 4394 56058
rect 4394 56006 4406 56058
rect 4406 56006 4436 56058
rect 4460 56006 4470 56058
rect 4470 56006 4516 56058
rect 4220 56004 4276 56006
rect 4300 56004 4356 56006
rect 4380 56004 4436 56006
rect 4460 56004 4516 56006
rect 4220 54970 4276 54972
rect 4300 54970 4356 54972
rect 4380 54970 4436 54972
rect 4460 54970 4516 54972
rect 4220 54918 4266 54970
rect 4266 54918 4276 54970
rect 4300 54918 4330 54970
rect 4330 54918 4342 54970
rect 4342 54918 4356 54970
rect 4380 54918 4394 54970
rect 4394 54918 4406 54970
rect 4406 54918 4436 54970
rect 4460 54918 4470 54970
rect 4470 54918 4516 54970
rect 4220 54916 4276 54918
rect 4300 54916 4356 54918
rect 4380 54916 4436 54918
rect 4460 54916 4516 54918
rect 4220 53882 4276 53884
rect 4300 53882 4356 53884
rect 4380 53882 4436 53884
rect 4460 53882 4516 53884
rect 4220 53830 4266 53882
rect 4266 53830 4276 53882
rect 4300 53830 4330 53882
rect 4330 53830 4342 53882
rect 4342 53830 4356 53882
rect 4380 53830 4394 53882
rect 4394 53830 4406 53882
rect 4406 53830 4436 53882
rect 4460 53830 4470 53882
rect 4470 53830 4516 53882
rect 4220 53828 4276 53830
rect 4300 53828 4356 53830
rect 4380 53828 4436 53830
rect 4460 53828 4516 53830
rect 4220 52794 4276 52796
rect 4300 52794 4356 52796
rect 4380 52794 4436 52796
rect 4460 52794 4516 52796
rect 4220 52742 4266 52794
rect 4266 52742 4276 52794
rect 4300 52742 4330 52794
rect 4330 52742 4342 52794
rect 4342 52742 4356 52794
rect 4380 52742 4394 52794
rect 4394 52742 4406 52794
rect 4406 52742 4436 52794
rect 4460 52742 4470 52794
rect 4470 52742 4516 52794
rect 4220 52740 4276 52742
rect 4300 52740 4356 52742
rect 4380 52740 4436 52742
rect 4460 52740 4516 52742
rect 4220 51706 4276 51708
rect 4300 51706 4356 51708
rect 4380 51706 4436 51708
rect 4460 51706 4516 51708
rect 4220 51654 4266 51706
rect 4266 51654 4276 51706
rect 4300 51654 4330 51706
rect 4330 51654 4342 51706
rect 4342 51654 4356 51706
rect 4380 51654 4394 51706
rect 4394 51654 4406 51706
rect 4406 51654 4436 51706
rect 4460 51654 4470 51706
rect 4470 51654 4516 51706
rect 4220 51652 4276 51654
rect 4300 51652 4356 51654
rect 4380 51652 4436 51654
rect 4460 51652 4516 51654
rect 4220 50618 4276 50620
rect 4300 50618 4356 50620
rect 4380 50618 4436 50620
rect 4460 50618 4516 50620
rect 4220 50566 4266 50618
rect 4266 50566 4276 50618
rect 4300 50566 4330 50618
rect 4330 50566 4342 50618
rect 4342 50566 4356 50618
rect 4380 50566 4394 50618
rect 4394 50566 4406 50618
rect 4406 50566 4436 50618
rect 4460 50566 4470 50618
rect 4470 50566 4516 50618
rect 4220 50564 4276 50566
rect 4300 50564 4356 50566
rect 4380 50564 4436 50566
rect 4460 50564 4516 50566
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 3422 35128 3478 35184
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 1582 27512 1638 27568
rect 1582 26152 1638 26208
rect 938 24248 994 24304
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 938 22616 994 22672
rect 938 20984 994 21040
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 7286 35164 7288 35184
rect 7288 35164 7340 35184
rect 7340 35164 7342 35184
rect 7286 35128 7342 35164
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 5630 25880 5686 25936
rect 938 19352 994 19408
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 1582 17856 1638 17912
rect 938 16108 994 16144
rect 938 16088 940 16108
rect 940 16088 992 16108
rect 992 16088 994 16108
rect 938 14456 994 14512
rect 938 12824 994 12880
rect 938 11192 994 11248
rect 1582 9560 1638 9616
rect 1582 8200 1638 8256
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 9034 25900 9090 25936
rect 9034 25880 9036 25900
rect 9036 25880 9088 25900
rect 9088 25880 9090 25900
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 938 6296 994 6352
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 938 4664 994 4720
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 938 3032 994 3088
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 57690 19636 57692
rect 19660 57690 19716 57692
rect 19740 57690 19796 57692
rect 19820 57690 19876 57692
rect 19580 57638 19626 57690
rect 19626 57638 19636 57690
rect 19660 57638 19690 57690
rect 19690 57638 19702 57690
rect 19702 57638 19716 57690
rect 19740 57638 19754 57690
rect 19754 57638 19766 57690
rect 19766 57638 19796 57690
rect 19820 57638 19830 57690
rect 19830 57638 19876 57690
rect 19580 57636 19636 57638
rect 19660 57636 19716 57638
rect 19740 57636 19796 57638
rect 19820 57636 19876 57638
rect 50300 57690 50356 57692
rect 50380 57690 50436 57692
rect 50460 57690 50516 57692
rect 50540 57690 50596 57692
rect 50300 57638 50346 57690
rect 50346 57638 50356 57690
rect 50380 57638 50410 57690
rect 50410 57638 50422 57690
rect 50422 57638 50436 57690
rect 50460 57638 50474 57690
rect 50474 57638 50486 57690
rect 50486 57638 50516 57690
rect 50540 57638 50550 57690
rect 50550 57638 50596 57690
rect 50300 57636 50356 57638
rect 50380 57636 50436 57638
rect 50460 57636 50516 57638
rect 50540 57636 50596 57638
rect 34940 57146 34996 57148
rect 35020 57146 35076 57148
rect 35100 57146 35156 57148
rect 35180 57146 35236 57148
rect 34940 57094 34986 57146
rect 34986 57094 34996 57146
rect 35020 57094 35050 57146
rect 35050 57094 35062 57146
rect 35062 57094 35076 57146
rect 35100 57094 35114 57146
rect 35114 57094 35126 57146
rect 35126 57094 35156 57146
rect 35180 57094 35190 57146
rect 35190 57094 35236 57146
rect 34940 57092 34996 57094
rect 35020 57092 35076 57094
rect 35100 57092 35156 57094
rect 35180 57092 35236 57094
rect 19580 56602 19636 56604
rect 19660 56602 19716 56604
rect 19740 56602 19796 56604
rect 19820 56602 19876 56604
rect 19580 56550 19626 56602
rect 19626 56550 19636 56602
rect 19660 56550 19690 56602
rect 19690 56550 19702 56602
rect 19702 56550 19716 56602
rect 19740 56550 19754 56602
rect 19754 56550 19766 56602
rect 19766 56550 19796 56602
rect 19820 56550 19830 56602
rect 19830 56550 19876 56602
rect 19580 56548 19636 56550
rect 19660 56548 19716 56550
rect 19740 56548 19796 56550
rect 19820 56548 19876 56550
rect 34940 56058 34996 56060
rect 35020 56058 35076 56060
rect 35100 56058 35156 56060
rect 35180 56058 35236 56060
rect 34940 56006 34986 56058
rect 34986 56006 34996 56058
rect 35020 56006 35050 56058
rect 35050 56006 35062 56058
rect 35062 56006 35076 56058
rect 35100 56006 35114 56058
rect 35114 56006 35126 56058
rect 35126 56006 35156 56058
rect 35180 56006 35190 56058
rect 35190 56006 35236 56058
rect 34940 56004 34996 56006
rect 35020 56004 35076 56006
rect 35100 56004 35156 56006
rect 35180 56004 35236 56006
rect 19580 55514 19636 55516
rect 19660 55514 19716 55516
rect 19740 55514 19796 55516
rect 19820 55514 19876 55516
rect 19580 55462 19626 55514
rect 19626 55462 19636 55514
rect 19660 55462 19690 55514
rect 19690 55462 19702 55514
rect 19702 55462 19716 55514
rect 19740 55462 19754 55514
rect 19754 55462 19766 55514
rect 19766 55462 19796 55514
rect 19820 55462 19830 55514
rect 19830 55462 19876 55514
rect 19580 55460 19636 55462
rect 19660 55460 19716 55462
rect 19740 55460 19796 55462
rect 19820 55460 19876 55462
rect 34940 54970 34996 54972
rect 35020 54970 35076 54972
rect 35100 54970 35156 54972
rect 35180 54970 35236 54972
rect 34940 54918 34986 54970
rect 34986 54918 34996 54970
rect 35020 54918 35050 54970
rect 35050 54918 35062 54970
rect 35062 54918 35076 54970
rect 35100 54918 35114 54970
rect 35114 54918 35126 54970
rect 35126 54918 35156 54970
rect 35180 54918 35190 54970
rect 35190 54918 35236 54970
rect 34940 54916 34996 54918
rect 35020 54916 35076 54918
rect 35100 54916 35156 54918
rect 35180 54916 35236 54918
rect 19580 54426 19636 54428
rect 19660 54426 19716 54428
rect 19740 54426 19796 54428
rect 19820 54426 19876 54428
rect 19580 54374 19626 54426
rect 19626 54374 19636 54426
rect 19660 54374 19690 54426
rect 19690 54374 19702 54426
rect 19702 54374 19716 54426
rect 19740 54374 19754 54426
rect 19754 54374 19766 54426
rect 19766 54374 19796 54426
rect 19820 54374 19830 54426
rect 19830 54374 19876 54426
rect 19580 54372 19636 54374
rect 19660 54372 19716 54374
rect 19740 54372 19796 54374
rect 19820 54372 19876 54374
rect 34940 53882 34996 53884
rect 35020 53882 35076 53884
rect 35100 53882 35156 53884
rect 35180 53882 35236 53884
rect 34940 53830 34986 53882
rect 34986 53830 34996 53882
rect 35020 53830 35050 53882
rect 35050 53830 35062 53882
rect 35062 53830 35076 53882
rect 35100 53830 35114 53882
rect 35114 53830 35126 53882
rect 35126 53830 35156 53882
rect 35180 53830 35190 53882
rect 35190 53830 35236 53882
rect 34940 53828 34996 53830
rect 35020 53828 35076 53830
rect 35100 53828 35156 53830
rect 35180 53828 35236 53830
rect 19580 53338 19636 53340
rect 19660 53338 19716 53340
rect 19740 53338 19796 53340
rect 19820 53338 19876 53340
rect 19580 53286 19626 53338
rect 19626 53286 19636 53338
rect 19660 53286 19690 53338
rect 19690 53286 19702 53338
rect 19702 53286 19716 53338
rect 19740 53286 19754 53338
rect 19754 53286 19766 53338
rect 19766 53286 19796 53338
rect 19820 53286 19830 53338
rect 19830 53286 19876 53338
rect 19580 53284 19636 53286
rect 19660 53284 19716 53286
rect 19740 53284 19796 53286
rect 19820 53284 19876 53286
rect 34940 52794 34996 52796
rect 35020 52794 35076 52796
rect 35100 52794 35156 52796
rect 35180 52794 35236 52796
rect 34940 52742 34986 52794
rect 34986 52742 34996 52794
rect 35020 52742 35050 52794
rect 35050 52742 35062 52794
rect 35062 52742 35076 52794
rect 35100 52742 35114 52794
rect 35114 52742 35126 52794
rect 35126 52742 35156 52794
rect 35180 52742 35190 52794
rect 35190 52742 35236 52794
rect 34940 52740 34996 52742
rect 35020 52740 35076 52742
rect 35100 52740 35156 52742
rect 35180 52740 35236 52742
rect 19580 52250 19636 52252
rect 19660 52250 19716 52252
rect 19740 52250 19796 52252
rect 19820 52250 19876 52252
rect 19580 52198 19626 52250
rect 19626 52198 19636 52250
rect 19660 52198 19690 52250
rect 19690 52198 19702 52250
rect 19702 52198 19716 52250
rect 19740 52198 19754 52250
rect 19754 52198 19766 52250
rect 19766 52198 19796 52250
rect 19820 52198 19830 52250
rect 19830 52198 19876 52250
rect 19580 52196 19636 52198
rect 19660 52196 19716 52198
rect 19740 52196 19796 52198
rect 19820 52196 19876 52198
rect 34940 51706 34996 51708
rect 35020 51706 35076 51708
rect 35100 51706 35156 51708
rect 35180 51706 35236 51708
rect 34940 51654 34986 51706
rect 34986 51654 34996 51706
rect 35020 51654 35050 51706
rect 35050 51654 35062 51706
rect 35062 51654 35076 51706
rect 35100 51654 35114 51706
rect 35114 51654 35126 51706
rect 35126 51654 35156 51706
rect 35180 51654 35190 51706
rect 35190 51654 35236 51706
rect 34940 51652 34996 51654
rect 35020 51652 35076 51654
rect 35100 51652 35156 51654
rect 35180 51652 35236 51654
rect 19580 51162 19636 51164
rect 19660 51162 19716 51164
rect 19740 51162 19796 51164
rect 19820 51162 19876 51164
rect 19580 51110 19626 51162
rect 19626 51110 19636 51162
rect 19660 51110 19690 51162
rect 19690 51110 19702 51162
rect 19702 51110 19716 51162
rect 19740 51110 19754 51162
rect 19754 51110 19766 51162
rect 19766 51110 19796 51162
rect 19820 51110 19830 51162
rect 19830 51110 19876 51162
rect 19580 51108 19636 51110
rect 19660 51108 19716 51110
rect 19740 51108 19796 51110
rect 19820 51108 19876 51110
rect 34940 50618 34996 50620
rect 35020 50618 35076 50620
rect 35100 50618 35156 50620
rect 35180 50618 35236 50620
rect 34940 50566 34986 50618
rect 34986 50566 34996 50618
rect 35020 50566 35050 50618
rect 35050 50566 35062 50618
rect 35062 50566 35076 50618
rect 35100 50566 35114 50618
rect 35114 50566 35126 50618
rect 35126 50566 35156 50618
rect 35180 50566 35190 50618
rect 35190 50566 35236 50618
rect 34940 50564 34996 50566
rect 35020 50564 35076 50566
rect 35100 50564 35156 50566
rect 35180 50564 35236 50566
rect 19580 50074 19636 50076
rect 19660 50074 19716 50076
rect 19740 50074 19796 50076
rect 19820 50074 19876 50076
rect 19580 50022 19626 50074
rect 19626 50022 19636 50074
rect 19660 50022 19690 50074
rect 19690 50022 19702 50074
rect 19702 50022 19716 50074
rect 19740 50022 19754 50074
rect 19754 50022 19766 50074
rect 19766 50022 19796 50074
rect 19820 50022 19830 50074
rect 19830 50022 19876 50074
rect 19580 50020 19636 50022
rect 19660 50020 19716 50022
rect 19740 50020 19796 50022
rect 19820 50020 19876 50022
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 44086 33108 44142 33144
rect 44086 33088 44088 33108
rect 44088 33088 44140 33108
rect 44140 33088 44142 33108
rect 41326 28076 41382 28112
rect 41326 28056 41328 28076
rect 41328 28056 41380 28076
rect 41380 28056 41382 28076
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 50300 56602 50356 56604
rect 50380 56602 50436 56604
rect 50460 56602 50516 56604
rect 50540 56602 50596 56604
rect 50300 56550 50346 56602
rect 50346 56550 50356 56602
rect 50380 56550 50410 56602
rect 50410 56550 50422 56602
rect 50422 56550 50436 56602
rect 50460 56550 50474 56602
rect 50474 56550 50486 56602
rect 50486 56550 50516 56602
rect 50540 56550 50550 56602
rect 50550 56550 50596 56602
rect 50300 56548 50356 56550
rect 50380 56548 50436 56550
rect 50460 56548 50516 56550
rect 50540 56548 50596 56550
rect 50300 55514 50356 55516
rect 50380 55514 50436 55516
rect 50460 55514 50516 55516
rect 50540 55514 50596 55516
rect 50300 55462 50346 55514
rect 50346 55462 50356 55514
rect 50380 55462 50410 55514
rect 50410 55462 50422 55514
rect 50422 55462 50436 55514
rect 50460 55462 50474 55514
rect 50474 55462 50486 55514
rect 50486 55462 50516 55514
rect 50540 55462 50550 55514
rect 50550 55462 50596 55514
rect 50300 55460 50356 55462
rect 50380 55460 50436 55462
rect 50460 55460 50516 55462
rect 50540 55460 50596 55462
rect 50300 54426 50356 54428
rect 50380 54426 50436 54428
rect 50460 54426 50516 54428
rect 50540 54426 50596 54428
rect 50300 54374 50346 54426
rect 50346 54374 50356 54426
rect 50380 54374 50410 54426
rect 50410 54374 50422 54426
rect 50422 54374 50436 54426
rect 50460 54374 50474 54426
rect 50474 54374 50486 54426
rect 50486 54374 50516 54426
rect 50540 54374 50550 54426
rect 50550 54374 50596 54426
rect 50300 54372 50356 54374
rect 50380 54372 50436 54374
rect 50460 54372 50516 54374
rect 50540 54372 50596 54374
rect 50300 53338 50356 53340
rect 50380 53338 50436 53340
rect 50460 53338 50516 53340
rect 50540 53338 50596 53340
rect 50300 53286 50346 53338
rect 50346 53286 50356 53338
rect 50380 53286 50410 53338
rect 50410 53286 50422 53338
rect 50422 53286 50436 53338
rect 50460 53286 50474 53338
rect 50474 53286 50486 53338
rect 50486 53286 50516 53338
rect 50540 53286 50550 53338
rect 50550 53286 50596 53338
rect 50300 53284 50356 53286
rect 50380 53284 50436 53286
rect 50460 53284 50516 53286
rect 50540 53284 50596 53286
rect 58898 52808 58954 52864
rect 50300 52250 50356 52252
rect 50380 52250 50436 52252
rect 50460 52250 50516 52252
rect 50540 52250 50596 52252
rect 50300 52198 50346 52250
rect 50346 52198 50356 52250
rect 50380 52198 50410 52250
rect 50410 52198 50422 52250
rect 50422 52198 50436 52250
rect 50460 52198 50474 52250
rect 50474 52198 50486 52250
rect 50486 52198 50516 52250
rect 50540 52198 50550 52250
rect 50550 52198 50596 52250
rect 50300 52196 50356 52198
rect 50380 52196 50436 52198
rect 50460 52196 50516 52198
rect 50540 52196 50596 52198
rect 50300 51162 50356 51164
rect 50380 51162 50436 51164
rect 50460 51162 50516 51164
rect 50540 51162 50596 51164
rect 50300 51110 50346 51162
rect 50346 51110 50356 51162
rect 50380 51110 50410 51162
rect 50410 51110 50422 51162
rect 50422 51110 50436 51162
rect 50460 51110 50474 51162
rect 50474 51110 50486 51162
rect 50486 51110 50516 51162
rect 50540 51110 50550 51162
rect 50550 51110 50596 51162
rect 50300 51108 50356 51110
rect 50380 51108 50436 51110
rect 50460 51108 50516 51110
rect 50540 51108 50596 51110
rect 50300 50074 50356 50076
rect 50380 50074 50436 50076
rect 50460 50074 50516 50076
rect 50540 50074 50596 50076
rect 50300 50022 50346 50074
rect 50346 50022 50356 50074
rect 50380 50022 50410 50074
rect 50410 50022 50422 50074
rect 50422 50022 50436 50074
rect 50460 50022 50474 50074
rect 50474 50022 50486 50074
rect 50486 50022 50516 50074
rect 50540 50022 50550 50074
rect 50550 50022 50596 50074
rect 50300 50020 50356 50022
rect 50380 50020 50436 50022
rect 50460 50020 50516 50022
rect 50540 50020 50596 50022
rect 50300 48986 50356 48988
rect 50380 48986 50436 48988
rect 50460 48986 50516 48988
rect 50540 48986 50596 48988
rect 50300 48934 50346 48986
rect 50346 48934 50356 48986
rect 50380 48934 50410 48986
rect 50410 48934 50422 48986
rect 50422 48934 50436 48986
rect 50460 48934 50474 48986
rect 50474 48934 50486 48986
rect 50486 48934 50516 48986
rect 50540 48934 50550 48986
rect 50550 48934 50596 48986
rect 50300 48932 50356 48934
rect 50380 48932 50436 48934
rect 50460 48932 50516 48934
rect 50540 48932 50596 48934
rect 50300 47898 50356 47900
rect 50380 47898 50436 47900
rect 50460 47898 50516 47900
rect 50540 47898 50596 47900
rect 50300 47846 50346 47898
rect 50346 47846 50356 47898
rect 50380 47846 50410 47898
rect 50410 47846 50422 47898
rect 50422 47846 50436 47898
rect 50460 47846 50474 47898
rect 50474 47846 50486 47898
rect 50486 47846 50516 47898
rect 50540 47846 50550 47898
rect 50550 47846 50596 47898
rect 50300 47844 50356 47846
rect 50380 47844 50436 47846
rect 50460 47844 50516 47846
rect 50540 47844 50596 47846
rect 50300 46810 50356 46812
rect 50380 46810 50436 46812
rect 50460 46810 50516 46812
rect 50540 46810 50596 46812
rect 50300 46758 50346 46810
rect 50346 46758 50356 46810
rect 50380 46758 50410 46810
rect 50410 46758 50422 46810
rect 50422 46758 50436 46810
rect 50460 46758 50474 46810
rect 50474 46758 50486 46810
rect 50486 46758 50516 46810
rect 50540 46758 50550 46810
rect 50550 46758 50596 46810
rect 50300 46756 50356 46758
rect 50380 46756 50436 46758
rect 50460 46756 50516 46758
rect 50540 46756 50596 46758
rect 50300 45722 50356 45724
rect 50380 45722 50436 45724
rect 50460 45722 50516 45724
rect 50540 45722 50596 45724
rect 50300 45670 50346 45722
rect 50346 45670 50356 45722
rect 50380 45670 50410 45722
rect 50410 45670 50422 45722
rect 50422 45670 50436 45722
rect 50460 45670 50474 45722
rect 50474 45670 50486 45722
rect 50486 45670 50516 45722
rect 50540 45670 50550 45722
rect 50550 45670 50596 45722
rect 50300 45668 50356 45670
rect 50380 45668 50436 45670
rect 50460 45668 50516 45670
rect 50540 45668 50596 45670
rect 50300 44634 50356 44636
rect 50380 44634 50436 44636
rect 50460 44634 50516 44636
rect 50540 44634 50596 44636
rect 50300 44582 50346 44634
rect 50346 44582 50356 44634
rect 50380 44582 50410 44634
rect 50410 44582 50422 44634
rect 50422 44582 50436 44634
rect 50460 44582 50474 44634
rect 50474 44582 50486 44634
rect 50486 44582 50516 44634
rect 50540 44582 50550 44634
rect 50550 44582 50596 44634
rect 50300 44580 50356 44582
rect 50380 44580 50436 44582
rect 50460 44580 50516 44582
rect 50540 44580 50596 44582
rect 50300 43546 50356 43548
rect 50380 43546 50436 43548
rect 50460 43546 50516 43548
rect 50540 43546 50596 43548
rect 50300 43494 50346 43546
rect 50346 43494 50356 43546
rect 50380 43494 50410 43546
rect 50410 43494 50422 43546
rect 50422 43494 50436 43546
rect 50460 43494 50474 43546
rect 50474 43494 50486 43546
rect 50486 43494 50516 43546
rect 50540 43494 50550 43546
rect 50550 43494 50596 43546
rect 50300 43492 50356 43494
rect 50380 43492 50436 43494
rect 50460 43492 50516 43494
rect 50540 43492 50596 43494
rect 50300 42458 50356 42460
rect 50380 42458 50436 42460
rect 50460 42458 50516 42460
rect 50540 42458 50596 42460
rect 50300 42406 50346 42458
rect 50346 42406 50356 42458
rect 50380 42406 50410 42458
rect 50410 42406 50422 42458
rect 50422 42406 50436 42458
rect 50460 42406 50474 42458
rect 50474 42406 50486 42458
rect 50486 42406 50516 42458
rect 50540 42406 50550 42458
rect 50550 42406 50596 42458
rect 50300 42404 50356 42406
rect 50380 42404 50436 42406
rect 50460 42404 50516 42406
rect 50540 42404 50596 42406
rect 50300 41370 50356 41372
rect 50380 41370 50436 41372
rect 50460 41370 50516 41372
rect 50540 41370 50596 41372
rect 50300 41318 50346 41370
rect 50346 41318 50356 41370
rect 50380 41318 50410 41370
rect 50410 41318 50422 41370
rect 50422 41318 50436 41370
rect 50460 41318 50474 41370
rect 50474 41318 50486 41370
rect 50486 41318 50516 41370
rect 50540 41318 50550 41370
rect 50550 41318 50596 41370
rect 50300 41316 50356 41318
rect 50380 41316 50436 41318
rect 50460 41316 50516 41318
rect 50540 41316 50596 41318
rect 46110 33108 46166 33144
rect 46110 33088 46112 33108
rect 46112 33088 46164 33108
rect 46164 33088 46166 33108
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 44454 26324 44456 26344
rect 44456 26324 44508 26344
rect 44508 26324 44510 26344
rect 44454 26288 44510 26324
rect 50300 40282 50356 40284
rect 50380 40282 50436 40284
rect 50460 40282 50516 40284
rect 50540 40282 50596 40284
rect 50300 40230 50346 40282
rect 50346 40230 50356 40282
rect 50380 40230 50410 40282
rect 50410 40230 50422 40282
rect 50422 40230 50436 40282
rect 50460 40230 50474 40282
rect 50474 40230 50486 40282
rect 50486 40230 50516 40282
rect 50540 40230 50550 40282
rect 50550 40230 50596 40282
rect 50300 40228 50356 40230
rect 50380 40228 50436 40230
rect 50460 40228 50516 40230
rect 50540 40228 50596 40230
rect 50300 39194 50356 39196
rect 50380 39194 50436 39196
rect 50460 39194 50516 39196
rect 50540 39194 50596 39196
rect 50300 39142 50346 39194
rect 50346 39142 50356 39194
rect 50380 39142 50410 39194
rect 50410 39142 50422 39194
rect 50422 39142 50436 39194
rect 50460 39142 50474 39194
rect 50474 39142 50486 39194
rect 50486 39142 50516 39194
rect 50540 39142 50550 39194
rect 50550 39142 50596 39194
rect 50300 39140 50356 39142
rect 50380 39140 50436 39142
rect 50460 39140 50516 39142
rect 50540 39140 50596 39142
rect 50300 38106 50356 38108
rect 50380 38106 50436 38108
rect 50460 38106 50516 38108
rect 50540 38106 50596 38108
rect 50300 38054 50346 38106
rect 50346 38054 50356 38106
rect 50380 38054 50410 38106
rect 50410 38054 50422 38106
rect 50422 38054 50436 38106
rect 50460 38054 50474 38106
rect 50474 38054 50486 38106
rect 50486 38054 50516 38106
rect 50540 38054 50550 38106
rect 50550 38054 50596 38106
rect 50300 38052 50356 38054
rect 50380 38052 50436 38054
rect 50460 38052 50516 38054
rect 50540 38052 50596 38054
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 46110 27124 46166 27160
rect 46110 27104 46112 27124
rect 46112 27104 46164 27124
rect 46164 27104 46166 27124
rect 47582 28076 47638 28112
rect 47582 28056 47584 28076
rect 47584 28056 47636 28076
rect 47636 28056 47638 28076
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 48318 27412 48320 27432
rect 48320 27412 48372 27432
rect 48372 27412 48374 27432
rect 48318 27376 48374 27412
rect 48134 26288 48190 26344
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 49606 27104 49662 27160
rect 49790 25644 49792 25664
rect 49792 25644 49844 25664
rect 49844 25644 49846 25664
rect 49790 25608 49846 25644
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50710 28600 50766 28656
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50158 28076 50214 28112
rect 50158 28056 50160 28076
rect 50160 28056 50212 28076
rect 50212 28056 50214 28076
rect 50066 27648 50122 27704
rect 50618 27548 50620 27568
rect 50620 27548 50672 27568
rect 50672 27548 50674 27568
rect 50618 27512 50674 27548
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 51538 29416 51594 29472
rect 51354 29180 51356 29200
rect 51356 29180 51408 29200
rect 51408 29180 51410 29200
rect 51354 29144 51410 29180
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 52918 29416 52974 29472
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 49606 18400 49662 18456
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50342 20440 50398 20496
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50618 18808 50674 18864
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 53470 29008 53526 29064
rect 57886 45464 57942 45520
rect 57794 39752 57850 39808
rect 58254 38936 58310 38992
rect 58346 38120 58402 38176
rect 58898 51992 58954 52048
rect 56322 28600 56378 28656
rect 58622 30796 58678 30832
rect 58622 30776 58624 30796
rect 58624 30776 58676 30796
rect 58676 30776 58678 30796
rect 57150 29008 57206 29064
rect 56230 27376 56286 27432
rect 58622 29960 58678 30016
rect 58898 51176 58954 51232
rect 58898 49544 58954 49600
rect 58898 48728 58954 48784
rect 58898 47912 58954 47968
rect 58898 47096 58954 47152
rect 58898 46280 58954 46336
rect 58806 43016 58862 43072
rect 58806 41384 58862 41440
rect 58990 44648 59046 44704
rect 58990 43832 59046 43888
rect 58990 42200 59046 42256
rect 58990 40568 59046 40624
rect 58530 29144 58586 29200
rect 56782 28092 56784 28112
rect 56784 28092 56836 28112
rect 56836 28092 56838 28112
rect 56782 28056 56838 28092
rect 58898 37324 58954 37360
rect 58898 37304 58900 37324
rect 58900 37304 58952 37324
rect 58952 37304 58954 37324
rect 58898 36488 58954 36544
rect 58898 35672 58954 35728
rect 58898 34856 58954 34912
rect 58898 34040 58954 34096
rect 58898 33224 58954 33280
rect 58898 32408 58954 32464
rect 58898 31592 58954 31648
rect 58898 28328 58954 28384
rect 58714 27512 58770 27568
rect 58898 26696 58954 26752
rect 58622 25900 58678 25936
rect 58622 25880 58624 25900
rect 58624 25880 58676 25900
rect 58676 25880 58678 25900
rect 58622 25064 58678 25120
rect 58714 24248 58770 24304
rect 51078 12708 51134 12744
rect 51078 12688 51080 12708
rect 51080 12688 51132 12708
rect 51132 12688 51134 12708
rect 58898 23432 58954 23488
rect 58806 22636 58862 22672
rect 58806 22616 58808 22636
rect 58808 22616 58860 22636
rect 58860 22616 58862 22636
rect 56138 19372 56194 19408
rect 56138 19352 56140 19372
rect 56140 19352 56192 19372
rect 56192 19352 56194 19372
rect 57610 19352 57666 19408
rect 58898 21800 58954 21856
rect 58714 20984 58770 21040
rect 58530 20204 58532 20224
rect 58532 20204 58584 20224
rect 58584 20204 58586 20224
rect 58530 20168 58586 20204
rect 58898 19352 58954 19408
rect 57794 17720 57850 17776
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 58254 18808 58310 18864
rect 58898 18536 58954 18592
rect 58898 16904 58954 16960
rect 54482 12688 54538 12744
rect 58898 16088 58954 16144
rect 58898 15272 58954 15328
rect 58898 14456 58954 14512
rect 58898 13640 58954 13696
rect 57978 12008 58034 12064
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 58714 12824 58770 12880
rect 58622 11192 58678 11248
rect 58898 10376 58954 10432
rect 58898 9560 58954 9616
rect 58898 8744 58954 8800
rect 58898 7928 58954 7984
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 58898 7112 58954 7168
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
<< metal3 >>
rect 19570 57696 19886 57697
rect 19570 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19886 57696
rect 19570 57631 19886 57632
rect 50290 57696 50606 57697
rect 50290 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50606 57696
rect 50290 57631 50606 57632
rect 4210 57152 4526 57153
rect 4210 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4526 57152
rect 4210 57087 4526 57088
rect 34930 57152 35246 57153
rect 34930 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35246 57152
rect 34930 57087 35246 57088
rect 0 56946 800 56976
rect 933 56946 999 56949
rect 0 56944 999 56946
rect 0 56888 938 56944
rect 994 56888 999 56944
rect 0 56886 999 56888
rect 0 56856 800 56886
rect 933 56883 999 56886
rect 19570 56608 19886 56609
rect 19570 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19886 56608
rect 19570 56543 19886 56544
rect 50290 56608 50606 56609
rect 50290 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50606 56608
rect 50290 56543 50606 56544
rect 4210 56064 4526 56065
rect 4210 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4526 56064
rect 4210 55999 4526 56000
rect 34930 56064 35246 56065
rect 34930 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35246 56064
rect 34930 55999 35246 56000
rect 19570 55520 19886 55521
rect 19570 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19886 55520
rect 19570 55455 19886 55456
rect 50290 55520 50606 55521
rect 50290 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50606 55520
rect 50290 55455 50606 55456
rect 0 55314 800 55344
rect 933 55314 999 55317
rect 0 55312 999 55314
rect 0 55256 938 55312
rect 994 55256 999 55312
rect 0 55254 999 55256
rect 0 55224 800 55254
rect 933 55251 999 55254
rect 4210 54976 4526 54977
rect 4210 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4526 54976
rect 4210 54911 4526 54912
rect 34930 54976 35246 54977
rect 34930 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35246 54976
rect 34930 54911 35246 54912
rect 19570 54432 19886 54433
rect 19570 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19886 54432
rect 19570 54367 19886 54368
rect 50290 54432 50606 54433
rect 50290 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50606 54432
rect 50290 54367 50606 54368
rect 4210 53888 4526 53889
rect 4210 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4526 53888
rect 4210 53823 4526 53824
rect 34930 53888 35246 53889
rect 34930 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35246 53888
rect 34930 53823 35246 53824
rect 1577 53816 1643 53821
rect 1577 53760 1582 53816
rect 1638 53760 1643 53816
rect 1577 53755 1643 53760
rect 0 53682 800 53712
rect 1580 53682 1640 53755
rect 0 53622 1640 53682
rect 0 53592 800 53622
rect 19570 53344 19886 53345
rect 19570 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19886 53344
rect 19570 53279 19886 53280
rect 50290 53344 50606 53345
rect 50290 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50606 53344
rect 50290 53279 50606 53280
rect 58893 52866 58959 52869
rect 59200 52866 60000 52896
rect 58893 52864 60000 52866
rect 58893 52808 58898 52864
rect 58954 52808 60000 52864
rect 58893 52806 60000 52808
rect 58893 52803 58959 52806
rect 4210 52800 4526 52801
rect 4210 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4526 52800
rect 4210 52735 4526 52736
rect 34930 52800 35246 52801
rect 34930 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35246 52800
rect 59200 52776 60000 52806
rect 34930 52735 35246 52736
rect 1577 52456 1643 52461
rect 1577 52400 1582 52456
rect 1638 52400 1643 52456
rect 1577 52395 1643 52400
rect 0 52050 800 52080
rect 1580 52050 1640 52395
rect 19570 52256 19886 52257
rect 19570 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19886 52256
rect 19570 52191 19886 52192
rect 50290 52256 50606 52257
rect 50290 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50606 52256
rect 50290 52191 50606 52192
rect 0 51990 1640 52050
rect 58893 52050 58959 52053
rect 59200 52050 60000 52080
rect 58893 52048 60000 52050
rect 58893 51992 58898 52048
rect 58954 51992 60000 52048
rect 58893 51990 60000 51992
rect 0 51960 800 51990
rect 58893 51987 58959 51990
rect 59200 51960 60000 51990
rect 4210 51712 4526 51713
rect 4210 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4526 51712
rect 4210 51647 4526 51648
rect 34930 51712 35246 51713
rect 34930 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35246 51712
rect 34930 51647 35246 51648
rect 58893 51234 58959 51237
rect 59200 51234 60000 51264
rect 58893 51232 60000 51234
rect 58893 51176 58898 51232
rect 58954 51176 60000 51232
rect 58893 51174 60000 51176
rect 58893 51171 58959 51174
rect 19570 51168 19886 51169
rect 19570 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19886 51168
rect 19570 51103 19886 51104
rect 50290 51168 50606 51169
rect 50290 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50606 51168
rect 59200 51144 60000 51174
rect 50290 51103 50606 51104
rect 4210 50624 4526 50625
rect 4210 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4526 50624
rect 4210 50559 4526 50560
rect 34930 50624 35246 50625
rect 34930 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35246 50624
rect 34930 50559 35246 50560
rect 0 50418 800 50448
rect 933 50418 999 50421
rect 0 50416 999 50418
rect 0 50360 938 50416
rect 994 50360 999 50416
rect 0 50358 999 50360
rect 0 50328 800 50358
rect 933 50355 999 50358
rect 59200 50328 60000 50448
rect 19570 50080 19886 50081
rect 19570 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19886 50080
rect 19570 50015 19886 50016
rect 50290 50080 50606 50081
rect 50290 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50606 50080
rect 50290 50015 50606 50016
rect 58893 49602 58959 49605
rect 59200 49602 60000 49632
rect 58893 49600 60000 49602
rect 58893 49544 58898 49600
rect 58954 49544 60000 49600
rect 58893 49542 60000 49544
rect 58893 49539 58959 49542
rect 4210 49536 4526 49537
rect 4210 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4526 49536
rect 4210 49471 4526 49472
rect 34930 49536 35246 49537
rect 34930 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35246 49536
rect 59200 49512 60000 49542
rect 34930 49471 35246 49472
rect 19570 48992 19886 48993
rect 19570 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19886 48992
rect 19570 48927 19886 48928
rect 50290 48992 50606 48993
rect 50290 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50606 48992
rect 50290 48927 50606 48928
rect 0 48786 800 48816
rect 933 48786 999 48789
rect 0 48784 999 48786
rect 0 48728 938 48784
rect 994 48728 999 48784
rect 0 48726 999 48728
rect 0 48696 800 48726
rect 933 48723 999 48726
rect 58893 48786 58959 48789
rect 59200 48786 60000 48816
rect 58893 48784 60000 48786
rect 58893 48728 58898 48784
rect 58954 48728 60000 48784
rect 58893 48726 60000 48728
rect 58893 48723 58959 48726
rect 59200 48696 60000 48726
rect 4210 48448 4526 48449
rect 4210 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4526 48448
rect 4210 48383 4526 48384
rect 34930 48448 35246 48449
rect 34930 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35246 48448
rect 34930 48383 35246 48384
rect 58893 47970 58959 47973
rect 59200 47970 60000 48000
rect 58893 47968 60000 47970
rect 58893 47912 58898 47968
rect 58954 47912 60000 47968
rect 58893 47910 60000 47912
rect 58893 47907 58959 47910
rect 19570 47904 19886 47905
rect 19570 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19886 47904
rect 19570 47839 19886 47840
rect 50290 47904 50606 47905
rect 50290 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50606 47904
rect 59200 47880 60000 47910
rect 50290 47839 50606 47840
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 0 47154 800 47184
rect 933 47154 999 47157
rect 0 47152 999 47154
rect 0 47096 938 47152
rect 994 47096 999 47152
rect 0 47094 999 47096
rect 0 47064 800 47094
rect 933 47091 999 47094
rect 58893 47154 58959 47157
rect 59200 47154 60000 47184
rect 58893 47152 60000 47154
rect 58893 47096 58898 47152
rect 58954 47096 60000 47152
rect 58893 47094 60000 47096
rect 58893 47091 58959 47094
rect 59200 47064 60000 47094
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 50290 46816 50606 46817
rect 50290 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50606 46816
rect 50290 46751 50606 46752
rect 58893 46338 58959 46341
rect 59200 46338 60000 46368
rect 58893 46336 60000 46338
rect 58893 46280 58898 46336
rect 58954 46280 60000 46336
rect 58893 46278 60000 46280
rect 58893 46275 58959 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 59200 46248 60000 46278
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 50290 45728 50606 45729
rect 50290 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50606 45728
rect 50290 45663 50606 45664
rect 0 45522 800 45552
rect 1577 45522 1643 45525
rect 0 45520 1643 45522
rect 0 45464 1582 45520
rect 1638 45464 1643 45520
rect 0 45462 1643 45464
rect 0 45432 800 45462
rect 1577 45459 1643 45462
rect 57881 45522 57947 45525
rect 59200 45522 60000 45552
rect 57881 45520 60000 45522
rect 57881 45464 57886 45520
rect 57942 45464 60000 45520
rect 57881 45462 60000 45464
rect 57881 45459 57947 45462
rect 59200 45432 60000 45462
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 58985 44706 59051 44709
rect 59200 44706 60000 44736
rect 58985 44704 60000 44706
rect 58985 44648 58990 44704
rect 59046 44648 60000 44704
rect 58985 44646 60000 44648
rect 58985 44643 59051 44646
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 50290 44640 50606 44641
rect 50290 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50606 44640
rect 59200 44616 60000 44646
rect 50290 44575 50606 44576
rect 1577 44162 1643 44165
rect 798 44160 1643 44162
rect 798 44104 1582 44160
rect 1638 44104 1643 44160
rect 798 44102 1643 44104
rect 798 43920 858 44102
rect 1577 44099 1643 44102
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 0 43830 858 43920
rect 58985 43890 59051 43893
rect 59200 43890 60000 43920
rect 58985 43888 60000 43890
rect 58985 43832 58990 43888
rect 59046 43832 60000 43888
rect 58985 43830 60000 43832
rect 0 43800 800 43830
rect 58985 43827 59051 43830
rect 59200 43800 60000 43830
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 19570 43487 19886 43488
rect 50290 43552 50606 43553
rect 50290 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50606 43552
rect 50290 43487 50606 43488
rect 58801 43074 58867 43077
rect 59200 43074 60000 43104
rect 58801 43072 60000 43074
rect 58801 43016 58806 43072
rect 58862 43016 60000 43072
rect 58801 43014 60000 43016
rect 58801 43011 58867 43014
rect 4210 43008 4526 43009
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 59200 42984 60000 43014
rect 34930 42943 35246 42944
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 50290 42464 50606 42465
rect 50290 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50606 42464
rect 50290 42399 50606 42400
rect 0 42258 800 42288
rect 933 42258 999 42261
rect 0 42256 999 42258
rect 0 42200 938 42256
rect 994 42200 999 42256
rect 0 42198 999 42200
rect 0 42168 800 42198
rect 933 42195 999 42198
rect 58985 42258 59051 42261
rect 59200 42258 60000 42288
rect 58985 42256 60000 42258
rect 58985 42200 58990 42256
rect 59046 42200 60000 42256
rect 58985 42198 60000 42200
rect 58985 42195 59051 42198
rect 59200 42168 60000 42198
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 58801 41442 58867 41445
rect 59200 41442 60000 41472
rect 58801 41440 60000 41442
rect 58801 41384 58806 41440
rect 58862 41384 60000 41440
rect 58801 41382 60000 41384
rect 58801 41379 58867 41382
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 50290 41376 50606 41377
rect 50290 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50606 41376
rect 59200 41352 60000 41382
rect 50290 41311 50606 41312
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 34930 40767 35246 40768
rect 0 40626 800 40656
rect 1209 40626 1275 40629
rect 0 40624 1275 40626
rect 0 40568 1214 40624
rect 1270 40568 1275 40624
rect 0 40566 1275 40568
rect 0 40536 800 40566
rect 1209 40563 1275 40566
rect 58985 40626 59051 40629
rect 59200 40626 60000 40656
rect 58985 40624 60000 40626
rect 58985 40568 58990 40624
rect 59046 40568 60000 40624
rect 58985 40566 60000 40568
rect 58985 40563 59051 40566
rect 59200 40536 60000 40566
rect 19570 40288 19886 40289
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 50290 40288 50606 40289
rect 50290 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50606 40288
rect 50290 40223 50606 40224
rect 57789 39810 57855 39813
rect 59200 39810 60000 39840
rect 57789 39808 60000 39810
rect 57789 39752 57794 39808
rect 57850 39752 60000 39808
rect 57789 39750 60000 39752
rect 57789 39747 57855 39750
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 59200 39720 60000 39750
rect 34930 39679 35246 39680
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 50290 39200 50606 39201
rect 50290 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50606 39200
rect 50290 39135 50606 39136
rect 0 38994 800 39024
rect 933 38994 999 38997
rect 0 38992 999 38994
rect 0 38936 938 38992
rect 994 38936 999 38992
rect 0 38934 999 38936
rect 0 38904 800 38934
rect 933 38931 999 38934
rect 58249 38994 58315 38997
rect 59200 38994 60000 39024
rect 58249 38992 60000 38994
rect 58249 38936 58254 38992
rect 58310 38936 60000 38992
rect 58249 38934 60000 38936
rect 58249 38931 58315 38934
rect 59200 38904 60000 38934
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 58341 38178 58407 38181
rect 59200 38178 60000 38208
rect 58341 38176 60000 38178
rect 58341 38120 58346 38176
rect 58402 38120 60000 38176
rect 58341 38118 60000 38120
rect 58341 38115 58407 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 19570 38047 19886 38048
rect 50290 38112 50606 38113
rect 50290 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50606 38112
rect 59200 38088 60000 38118
rect 50290 38047 50606 38048
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 0 37362 800 37392
rect 1577 37362 1643 37365
rect 0 37360 1643 37362
rect 0 37304 1582 37360
rect 1638 37304 1643 37360
rect 0 37302 1643 37304
rect 0 37272 800 37302
rect 1577 37299 1643 37302
rect 58893 37362 58959 37365
rect 59200 37362 60000 37392
rect 58893 37360 60000 37362
rect 58893 37304 58898 37360
rect 58954 37304 60000 37360
rect 58893 37302 60000 37304
rect 58893 37299 58959 37302
rect 59200 37272 60000 37302
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 50290 37024 50606 37025
rect 50290 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50606 37024
rect 50290 36959 50606 36960
rect 58893 36546 58959 36549
rect 59200 36546 60000 36576
rect 58893 36544 60000 36546
rect 58893 36488 58898 36544
rect 58954 36488 60000 36544
rect 58893 36486 60000 36488
rect 58893 36483 58959 36486
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 59200 36456 60000 36486
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 50290 35936 50606 35937
rect 50290 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50606 35936
rect 50290 35871 50606 35872
rect 0 35730 800 35760
rect 933 35730 999 35733
rect 0 35728 999 35730
rect 0 35672 938 35728
rect 994 35672 999 35728
rect 0 35670 999 35672
rect 0 35640 800 35670
rect 933 35667 999 35670
rect 58893 35730 58959 35733
rect 59200 35730 60000 35760
rect 58893 35728 60000 35730
rect 58893 35672 58898 35728
rect 58954 35672 60000 35728
rect 58893 35670 60000 35672
rect 58893 35667 58959 35670
rect 59200 35640 60000 35670
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 3417 35186 3483 35189
rect 7281 35186 7347 35189
rect 3417 35184 7347 35186
rect 3417 35128 3422 35184
rect 3478 35128 7286 35184
rect 7342 35128 7347 35184
rect 3417 35126 7347 35128
rect 3417 35123 3483 35126
rect 7281 35123 7347 35126
rect 58893 34914 58959 34917
rect 59200 34914 60000 34944
rect 58893 34912 60000 34914
rect 58893 34856 58898 34912
rect 58954 34856 60000 34912
rect 58893 34854 60000 34856
rect 58893 34851 58959 34854
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 50290 34848 50606 34849
rect 50290 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50606 34848
rect 59200 34824 60000 34854
rect 50290 34783 50606 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 0 34098 800 34128
rect 933 34098 999 34101
rect 0 34096 999 34098
rect 0 34040 938 34096
rect 994 34040 999 34096
rect 0 34038 999 34040
rect 0 34008 800 34038
rect 933 34035 999 34038
rect 58893 34098 58959 34101
rect 59200 34098 60000 34128
rect 58893 34096 60000 34098
rect 58893 34040 58898 34096
rect 58954 34040 60000 34096
rect 58893 34038 60000 34040
rect 58893 34035 58959 34038
rect 59200 34008 60000 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 50290 33760 50606 33761
rect 50290 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50606 33760
rect 50290 33695 50606 33696
rect 58893 33282 58959 33285
rect 59200 33282 60000 33312
rect 58893 33280 60000 33282
rect 58893 33224 58898 33280
rect 58954 33224 60000 33280
rect 58893 33222 60000 33224
rect 58893 33219 58959 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 59200 33192 60000 33222
rect 34930 33151 35246 33152
rect 44081 33146 44147 33149
rect 46105 33146 46171 33149
rect 44081 33144 46171 33146
rect 44081 33088 44086 33144
rect 44142 33088 46110 33144
rect 46166 33088 46171 33144
rect 44081 33086 46171 33088
rect 44081 33083 44147 33086
rect 46105 33083 46171 33086
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 50290 32672 50606 32673
rect 50290 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50606 32672
rect 50290 32607 50606 32608
rect 0 32466 800 32496
rect 933 32466 999 32469
rect 0 32464 999 32466
rect 0 32408 938 32464
rect 994 32408 999 32464
rect 0 32406 999 32408
rect 0 32376 800 32406
rect 933 32403 999 32406
rect 58893 32466 58959 32469
rect 59200 32466 60000 32496
rect 58893 32464 60000 32466
rect 58893 32408 58898 32464
rect 58954 32408 60000 32464
rect 58893 32406 60000 32408
rect 58893 32403 58959 32406
rect 59200 32376 60000 32406
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 58893 31650 58959 31653
rect 59200 31650 60000 31680
rect 58893 31648 60000 31650
rect 58893 31592 58898 31648
rect 58954 31592 60000 31648
rect 58893 31590 60000 31592
rect 58893 31587 58959 31590
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 50290 31584 50606 31585
rect 50290 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50606 31584
rect 59200 31560 60000 31590
rect 50290 31519 50606 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 0 30834 800 30864
rect 933 30834 999 30837
rect 0 30832 999 30834
rect 0 30776 938 30832
rect 994 30776 999 30832
rect 0 30774 999 30776
rect 0 30744 800 30774
rect 933 30771 999 30774
rect 58617 30834 58683 30837
rect 59200 30834 60000 30864
rect 58617 30832 60000 30834
rect 58617 30776 58622 30832
rect 58678 30776 60000 30832
rect 58617 30774 60000 30776
rect 58617 30771 58683 30774
rect 59200 30744 60000 30774
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 50290 30496 50606 30497
rect 50290 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50606 30496
rect 50290 30431 50606 30432
rect 58617 30018 58683 30021
rect 59200 30018 60000 30048
rect 58617 30016 60000 30018
rect 58617 29960 58622 30016
rect 58678 29960 60000 30016
rect 58617 29958 60000 29960
rect 58617 29955 58683 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 59200 29928 60000 29958
rect 34930 29887 35246 29888
rect 51533 29474 51599 29477
rect 52913 29474 52979 29477
rect 51533 29472 52979 29474
rect 51533 29416 51538 29472
rect 51594 29416 52918 29472
rect 52974 29416 52979 29472
rect 51533 29414 52979 29416
rect 51533 29411 51599 29414
rect 52913 29411 52979 29414
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 50290 29408 50606 29409
rect 50290 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50606 29408
rect 50290 29343 50606 29344
rect 0 29202 800 29232
rect 933 29202 999 29205
rect 0 29200 999 29202
rect 0 29144 938 29200
rect 994 29144 999 29200
rect 0 29142 999 29144
rect 0 29112 800 29142
rect 933 29139 999 29142
rect 51206 29140 51212 29204
rect 51276 29202 51282 29204
rect 51349 29202 51415 29205
rect 51276 29200 51415 29202
rect 51276 29144 51354 29200
rect 51410 29144 51415 29200
rect 51276 29142 51415 29144
rect 51276 29140 51282 29142
rect 51349 29139 51415 29142
rect 58525 29202 58591 29205
rect 59200 29202 60000 29232
rect 58525 29200 60000 29202
rect 58525 29144 58530 29200
rect 58586 29144 60000 29200
rect 58525 29142 60000 29144
rect 58525 29139 58591 29142
rect 59200 29112 60000 29142
rect 53465 29066 53531 29069
rect 57145 29066 57211 29069
rect 53465 29064 57211 29066
rect 53465 29008 53470 29064
rect 53526 29008 57150 29064
rect 57206 29008 57211 29064
rect 53465 29006 57211 29008
rect 53465 29003 53531 29006
rect 57145 29003 57211 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 50705 28658 50771 28661
rect 56317 28658 56383 28661
rect 50705 28656 56383 28658
rect 50705 28600 50710 28656
rect 50766 28600 56322 28656
rect 56378 28600 56383 28656
rect 50705 28598 56383 28600
rect 50705 28595 50771 28598
rect 56317 28595 56383 28598
rect 58893 28386 58959 28389
rect 59200 28386 60000 28416
rect 58893 28384 60000 28386
rect 58893 28328 58898 28384
rect 58954 28328 60000 28384
rect 58893 28326 60000 28328
rect 58893 28323 58959 28326
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 50290 28320 50606 28321
rect 50290 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50606 28320
rect 59200 28296 60000 28326
rect 50290 28255 50606 28256
rect 41321 28114 41387 28117
rect 47577 28114 47643 28117
rect 41321 28112 47643 28114
rect 41321 28056 41326 28112
rect 41382 28056 47582 28112
rect 47638 28056 47643 28112
rect 41321 28054 47643 28056
rect 41321 28051 41387 28054
rect 47577 28051 47643 28054
rect 50153 28114 50219 28117
rect 56777 28114 56843 28117
rect 50153 28112 56843 28114
rect 50153 28056 50158 28112
rect 50214 28056 56782 28112
rect 56838 28056 56843 28112
rect 50153 28054 56843 28056
rect 50153 28051 50219 28054
rect 56777 28051 56843 28054
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 50061 27708 50127 27709
rect 50061 27704 50108 27708
rect 50172 27706 50178 27708
rect 50061 27648 50066 27704
rect 50061 27644 50108 27648
rect 50172 27646 50218 27706
rect 50172 27644 50178 27646
rect 50061 27643 50127 27644
rect 0 27570 800 27600
rect 1577 27570 1643 27573
rect 0 27568 1643 27570
rect 0 27512 1582 27568
rect 1638 27512 1643 27568
rect 0 27510 1643 27512
rect 0 27480 800 27510
rect 1577 27507 1643 27510
rect 50613 27570 50679 27573
rect 51206 27570 51212 27572
rect 50613 27568 51212 27570
rect 50613 27512 50618 27568
rect 50674 27512 51212 27568
rect 50613 27510 51212 27512
rect 50613 27507 50679 27510
rect 51206 27508 51212 27510
rect 51276 27508 51282 27572
rect 58709 27570 58775 27573
rect 59200 27570 60000 27600
rect 58709 27568 60000 27570
rect 58709 27512 58714 27568
rect 58770 27512 60000 27568
rect 58709 27510 60000 27512
rect 58709 27507 58775 27510
rect 59200 27480 60000 27510
rect 48313 27434 48379 27437
rect 56225 27434 56291 27437
rect 48313 27432 56291 27434
rect 48313 27376 48318 27432
rect 48374 27376 56230 27432
rect 56286 27376 56291 27432
rect 48313 27374 56291 27376
rect 48313 27371 48379 27374
rect 56225 27371 56291 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 50290 27232 50606 27233
rect 50290 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50606 27232
rect 50290 27167 50606 27168
rect 46105 27162 46171 27165
rect 49601 27162 49667 27165
rect 46105 27160 49667 27162
rect 46105 27104 46110 27160
rect 46166 27104 49606 27160
rect 49662 27104 49667 27160
rect 46105 27102 49667 27104
rect 46105 27099 46171 27102
rect 49601 27099 49667 27102
rect 58893 26754 58959 26757
rect 59200 26754 60000 26784
rect 58893 26752 60000 26754
rect 58893 26696 58898 26752
rect 58954 26696 60000 26752
rect 58893 26694 60000 26696
rect 58893 26691 58959 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 59200 26664 60000 26694
rect 34930 26623 35246 26624
rect 44449 26346 44515 26349
rect 48129 26346 48195 26349
rect 44449 26344 48195 26346
rect 44449 26288 44454 26344
rect 44510 26288 48134 26344
rect 48190 26288 48195 26344
rect 44449 26286 48195 26288
rect 44449 26283 44515 26286
rect 48129 26283 48195 26286
rect 1577 26210 1643 26213
rect 798 26208 1643 26210
rect 798 26152 1582 26208
rect 1638 26152 1643 26208
rect 798 26150 1643 26152
rect 798 25968 858 26150
rect 1577 26147 1643 26150
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 50290 26144 50606 26145
rect 50290 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50606 26144
rect 50290 26079 50606 26080
rect 0 25878 858 25968
rect 5625 25938 5691 25941
rect 9029 25938 9095 25941
rect 5625 25936 9095 25938
rect 5625 25880 5630 25936
rect 5686 25880 9034 25936
rect 9090 25880 9095 25936
rect 5625 25878 9095 25880
rect 0 25848 800 25878
rect 5625 25875 5691 25878
rect 9029 25875 9095 25878
rect 58617 25938 58683 25941
rect 59200 25938 60000 25968
rect 58617 25936 60000 25938
rect 58617 25880 58622 25936
rect 58678 25880 60000 25936
rect 58617 25878 60000 25880
rect 58617 25875 58683 25878
rect 59200 25848 60000 25878
rect 49785 25668 49851 25669
rect 49734 25604 49740 25668
rect 49804 25666 49851 25668
rect 49804 25664 49896 25666
rect 49846 25608 49896 25664
rect 49804 25606 49896 25608
rect 49804 25604 49851 25606
rect 49785 25603 49851 25604
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 58617 25122 58683 25125
rect 59200 25122 60000 25152
rect 58617 25120 60000 25122
rect 58617 25064 58622 25120
rect 58678 25064 60000 25120
rect 58617 25062 60000 25064
rect 58617 25059 58683 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 50290 25056 50606 25057
rect 50290 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50606 25056
rect 59200 25032 60000 25062
rect 50290 24991 50606 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 0 24306 800 24336
rect 933 24306 999 24309
rect 0 24304 999 24306
rect 0 24248 938 24304
rect 994 24248 999 24304
rect 0 24246 999 24248
rect 0 24216 800 24246
rect 933 24243 999 24246
rect 58709 24306 58775 24309
rect 59200 24306 60000 24336
rect 58709 24304 60000 24306
rect 58709 24248 58714 24304
rect 58770 24248 60000 24304
rect 58709 24246 60000 24248
rect 58709 24243 58775 24246
rect 59200 24216 60000 24246
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 50290 23968 50606 23969
rect 50290 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50606 23968
rect 50290 23903 50606 23904
rect 58893 23490 58959 23493
rect 59200 23490 60000 23520
rect 58893 23488 60000 23490
rect 58893 23432 58898 23488
rect 58954 23432 60000 23488
rect 58893 23430 60000 23432
rect 58893 23427 58959 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 59200 23400 60000 23430
rect 34930 23359 35246 23360
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 50290 22880 50606 22881
rect 50290 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50606 22880
rect 50290 22815 50606 22816
rect 0 22674 800 22704
rect 933 22674 999 22677
rect 0 22672 999 22674
rect 0 22616 938 22672
rect 994 22616 999 22672
rect 0 22614 999 22616
rect 0 22584 800 22614
rect 933 22611 999 22614
rect 58801 22674 58867 22677
rect 59200 22674 60000 22704
rect 58801 22672 60000 22674
rect 58801 22616 58806 22672
rect 58862 22616 60000 22672
rect 58801 22614 60000 22616
rect 58801 22611 58867 22614
rect 59200 22584 60000 22614
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 58893 21858 58959 21861
rect 59200 21858 60000 21888
rect 58893 21856 60000 21858
rect 58893 21800 58898 21856
rect 58954 21800 60000 21856
rect 58893 21798 60000 21800
rect 58893 21795 58959 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 50290 21792 50606 21793
rect 50290 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50606 21792
rect 59200 21768 60000 21798
rect 50290 21727 50606 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 0 21042 800 21072
rect 933 21042 999 21045
rect 0 21040 999 21042
rect 0 20984 938 21040
rect 994 20984 999 21040
rect 0 20982 999 20984
rect 0 20952 800 20982
rect 933 20979 999 20982
rect 58709 21042 58775 21045
rect 59200 21042 60000 21072
rect 58709 21040 60000 21042
rect 58709 20984 58714 21040
rect 58770 20984 60000 21040
rect 58709 20982 60000 20984
rect 58709 20979 58775 20982
rect 59200 20952 60000 20982
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 50290 20704 50606 20705
rect 50290 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50606 20704
rect 50290 20639 50606 20640
rect 50102 20436 50108 20500
rect 50172 20498 50178 20500
rect 50337 20498 50403 20501
rect 50172 20496 50403 20498
rect 50172 20440 50342 20496
rect 50398 20440 50403 20496
rect 50172 20438 50403 20440
rect 50172 20436 50178 20438
rect 50337 20435 50403 20438
rect 58525 20226 58591 20229
rect 59200 20226 60000 20256
rect 58525 20224 60000 20226
rect 58525 20168 58530 20224
rect 58586 20168 60000 20224
rect 58525 20166 60000 20168
rect 58525 20163 58591 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 59200 20136 60000 20166
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 50290 19616 50606 19617
rect 50290 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50606 19616
rect 50290 19551 50606 19552
rect 0 19410 800 19440
rect 933 19410 999 19413
rect 0 19408 999 19410
rect 0 19352 938 19408
rect 994 19352 999 19408
rect 0 19350 999 19352
rect 0 19320 800 19350
rect 933 19347 999 19350
rect 56133 19410 56199 19413
rect 57605 19410 57671 19413
rect 56133 19408 57671 19410
rect 56133 19352 56138 19408
rect 56194 19352 57610 19408
rect 57666 19352 57671 19408
rect 56133 19350 57671 19352
rect 56133 19347 56199 19350
rect 57605 19347 57671 19350
rect 58893 19410 58959 19413
rect 59200 19410 60000 19440
rect 58893 19408 60000 19410
rect 58893 19352 58898 19408
rect 58954 19352 60000 19408
rect 58893 19350 60000 19352
rect 58893 19347 58959 19350
rect 59200 19320 60000 19350
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 50613 18866 50679 18869
rect 58249 18866 58315 18869
rect 50613 18864 58315 18866
rect 50613 18808 50618 18864
rect 50674 18808 58254 18864
rect 58310 18808 58315 18864
rect 50613 18806 58315 18808
rect 50613 18803 50679 18806
rect 58249 18803 58315 18806
rect 58893 18594 58959 18597
rect 59200 18594 60000 18624
rect 58893 18592 60000 18594
rect 58893 18536 58898 18592
rect 58954 18536 60000 18592
rect 58893 18534 60000 18536
rect 58893 18531 58959 18534
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 50290 18528 50606 18529
rect 50290 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50606 18528
rect 59200 18504 60000 18534
rect 50290 18463 50606 18464
rect 49601 18458 49667 18461
rect 49734 18458 49740 18460
rect 49601 18456 49740 18458
rect 49601 18400 49606 18456
rect 49662 18400 49740 18456
rect 49601 18398 49740 18400
rect 49601 18395 49667 18398
rect 49734 18396 49740 18398
rect 49804 18396 49810 18460
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 1577 17914 1643 17917
rect 798 17912 1643 17914
rect 798 17856 1582 17912
rect 1638 17856 1643 17912
rect 798 17854 1643 17856
rect 798 17808 858 17854
rect 1577 17851 1643 17854
rect 0 17718 858 17808
rect 57789 17778 57855 17781
rect 59200 17778 60000 17808
rect 57789 17776 60000 17778
rect 57789 17720 57794 17776
rect 57850 17720 60000 17776
rect 57789 17718 60000 17720
rect 0 17688 800 17718
rect 57789 17715 57855 17718
rect 59200 17688 60000 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 50290 17440 50606 17441
rect 50290 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50606 17440
rect 50290 17375 50606 17376
rect 58893 16962 58959 16965
rect 59200 16962 60000 16992
rect 58893 16960 60000 16962
rect 58893 16904 58898 16960
rect 58954 16904 60000 16960
rect 58893 16902 60000 16904
rect 58893 16899 58959 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 59200 16872 60000 16902
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 50290 16352 50606 16353
rect 50290 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50606 16352
rect 50290 16287 50606 16288
rect 0 16146 800 16176
rect 933 16146 999 16149
rect 0 16144 999 16146
rect 0 16088 938 16144
rect 994 16088 999 16144
rect 0 16086 999 16088
rect 0 16056 800 16086
rect 933 16083 999 16086
rect 58893 16146 58959 16149
rect 59200 16146 60000 16176
rect 58893 16144 60000 16146
rect 58893 16088 58898 16144
rect 58954 16088 60000 16144
rect 58893 16086 60000 16088
rect 58893 16083 58959 16086
rect 59200 16056 60000 16086
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 58893 15330 58959 15333
rect 59200 15330 60000 15360
rect 58893 15328 60000 15330
rect 58893 15272 58898 15328
rect 58954 15272 60000 15328
rect 58893 15270 60000 15272
rect 58893 15267 58959 15270
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 50290 15264 50606 15265
rect 50290 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50606 15264
rect 59200 15240 60000 15270
rect 50290 15199 50606 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 0 14514 800 14544
rect 933 14514 999 14517
rect 0 14512 999 14514
rect 0 14456 938 14512
rect 994 14456 999 14512
rect 0 14454 999 14456
rect 0 14424 800 14454
rect 933 14451 999 14454
rect 58893 14514 58959 14517
rect 59200 14514 60000 14544
rect 58893 14512 60000 14514
rect 58893 14456 58898 14512
rect 58954 14456 60000 14512
rect 58893 14454 60000 14456
rect 58893 14451 58959 14454
rect 59200 14424 60000 14454
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 50290 14176 50606 14177
rect 50290 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50606 14176
rect 50290 14111 50606 14112
rect 58893 13698 58959 13701
rect 59200 13698 60000 13728
rect 58893 13696 60000 13698
rect 58893 13640 58898 13696
rect 58954 13640 60000 13696
rect 58893 13638 60000 13640
rect 58893 13635 58959 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 59200 13608 60000 13638
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 50290 13088 50606 13089
rect 50290 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50606 13088
rect 50290 13023 50606 13024
rect 0 12882 800 12912
rect 933 12882 999 12885
rect 0 12880 999 12882
rect 0 12824 938 12880
rect 994 12824 999 12880
rect 0 12822 999 12824
rect 0 12792 800 12822
rect 933 12819 999 12822
rect 58709 12882 58775 12885
rect 59200 12882 60000 12912
rect 58709 12880 60000 12882
rect 58709 12824 58714 12880
rect 58770 12824 60000 12880
rect 58709 12822 60000 12824
rect 58709 12819 58775 12822
rect 59200 12792 60000 12822
rect 51073 12746 51139 12749
rect 54477 12746 54543 12749
rect 51073 12744 54543 12746
rect 51073 12688 51078 12744
rect 51134 12688 54482 12744
rect 54538 12688 54543 12744
rect 51073 12686 54543 12688
rect 51073 12683 51139 12686
rect 54477 12683 54543 12686
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 57973 12066 58039 12069
rect 59200 12066 60000 12096
rect 57973 12064 60000 12066
rect 57973 12008 57978 12064
rect 58034 12008 60000 12064
rect 57973 12006 60000 12008
rect 57973 12003 58039 12006
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 50290 12000 50606 12001
rect 50290 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50606 12000
rect 59200 11976 60000 12006
rect 50290 11935 50606 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 0 11250 800 11280
rect 933 11250 999 11253
rect 0 11248 999 11250
rect 0 11192 938 11248
rect 994 11192 999 11248
rect 0 11190 999 11192
rect 0 11160 800 11190
rect 933 11187 999 11190
rect 58617 11250 58683 11253
rect 59200 11250 60000 11280
rect 58617 11248 60000 11250
rect 58617 11192 58622 11248
rect 58678 11192 60000 11248
rect 58617 11190 60000 11192
rect 58617 11187 58683 11190
rect 59200 11160 60000 11190
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 50290 10912 50606 10913
rect 50290 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50606 10912
rect 50290 10847 50606 10848
rect 58893 10434 58959 10437
rect 59200 10434 60000 10464
rect 58893 10432 60000 10434
rect 58893 10376 58898 10432
rect 58954 10376 60000 10432
rect 58893 10374 60000 10376
rect 58893 10371 58959 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 59200 10344 60000 10374
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 50290 9824 50606 9825
rect 50290 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50606 9824
rect 50290 9759 50606 9760
rect 0 9618 800 9648
rect 1577 9618 1643 9621
rect 0 9616 1643 9618
rect 0 9560 1582 9616
rect 1638 9560 1643 9616
rect 0 9558 1643 9560
rect 0 9528 800 9558
rect 1577 9555 1643 9558
rect 58893 9618 58959 9621
rect 59200 9618 60000 9648
rect 58893 9616 60000 9618
rect 58893 9560 58898 9616
rect 58954 9560 60000 9616
rect 58893 9558 60000 9560
rect 58893 9555 58959 9558
rect 59200 9528 60000 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 58893 8802 58959 8805
rect 59200 8802 60000 8832
rect 58893 8800 60000 8802
rect 58893 8744 58898 8800
rect 58954 8744 60000 8800
rect 58893 8742 60000 8744
rect 58893 8739 58959 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 50290 8736 50606 8737
rect 50290 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50606 8736
rect 59200 8712 60000 8742
rect 50290 8671 50606 8672
rect 1577 8258 1643 8261
rect 798 8256 1643 8258
rect 798 8200 1582 8256
rect 1638 8200 1643 8256
rect 798 8198 1643 8200
rect 798 8016 858 8198
rect 1577 8195 1643 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 0 7926 858 8016
rect 58893 7986 58959 7989
rect 59200 7986 60000 8016
rect 58893 7984 60000 7986
rect 58893 7928 58898 7984
rect 58954 7928 60000 7984
rect 58893 7926 60000 7928
rect 0 7896 800 7926
rect 58893 7923 58959 7926
rect 59200 7896 60000 7926
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 50290 7648 50606 7649
rect 50290 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50606 7648
rect 50290 7583 50606 7584
rect 58893 7170 58959 7173
rect 59200 7170 60000 7200
rect 58893 7168 60000 7170
rect 58893 7112 58898 7168
rect 58954 7112 60000 7168
rect 58893 7110 60000 7112
rect 58893 7107 58959 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 59200 7080 60000 7110
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 50290 6560 50606 6561
rect 50290 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50606 6560
rect 50290 6495 50606 6496
rect 0 6354 800 6384
rect 933 6354 999 6357
rect 0 6352 999 6354
rect 0 6296 938 6352
rect 994 6296 999 6352
rect 0 6294 999 6296
rect 0 6264 800 6294
rect 933 6291 999 6294
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 50290 5472 50606 5473
rect 50290 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50606 5472
rect 50290 5407 50606 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 0 4722 800 4752
rect 933 4722 999 4725
rect 0 4720 999 4722
rect 0 4664 938 4720
rect 994 4664 999 4720
rect 0 4662 999 4664
rect 0 4632 800 4662
rect 933 4659 999 4662
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 50290 4384 50606 4385
rect 50290 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50606 4384
rect 50290 4319 50606 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 50290 3296 50606 3297
rect 50290 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50606 3296
rect 50290 3231 50606 3232
rect 0 3090 800 3120
rect 933 3090 999 3093
rect 0 3088 999 3090
rect 0 3032 938 3088
rect 994 3032 999 3088
rect 0 3030 999 3032
rect 0 3000 800 3030
rect 933 3027 999 3030
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 50290 2208 50606 2209
rect 50290 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50606 2208
rect 50290 2143 50606 2144
<< via3 >>
rect 19576 57692 19640 57696
rect 19576 57636 19580 57692
rect 19580 57636 19636 57692
rect 19636 57636 19640 57692
rect 19576 57632 19640 57636
rect 19656 57692 19720 57696
rect 19656 57636 19660 57692
rect 19660 57636 19716 57692
rect 19716 57636 19720 57692
rect 19656 57632 19720 57636
rect 19736 57692 19800 57696
rect 19736 57636 19740 57692
rect 19740 57636 19796 57692
rect 19796 57636 19800 57692
rect 19736 57632 19800 57636
rect 19816 57692 19880 57696
rect 19816 57636 19820 57692
rect 19820 57636 19876 57692
rect 19876 57636 19880 57692
rect 19816 57632 19880 57636
rect 50296 57692 50360 57696
rect 50296 57636 50300 57692
rect 50300 57636 50356 57692
rect 50356 57636 50360 57692
rect 50296 57632 50360 57636
rect 50376 57692 50440 57696
rect 50376 57636 50380 57692
rect 50380 57636 50436 57692
rect 50436 57636 50440 57692
rect 50376 57632 50440 57636
rect 50456 57692 50520 57696
rect 50456 57636 50460 57692
rect 50460 57636 50516 57692
rect 50516 57636 50520 57692
rect 50456 57632 50520 57636
rect 50536 57692 50600 57696
rect 50536 57636 50540 57692
rect 50540 57636 50596 57692
rect 50596 57636 50600 57692
rect 50536 57632 50600 57636
rect 4216 57148 4280 57152
rect 4216 57092 4220 57148
rect 4220 57092 4276 57148
rect 4276 57092 4280 57148
rect 4216 57088 4280 57092
rect 4296 57148 4360 57152
rect 4296 57092 4300 57148
rect 4300 57092 4356 57148
rect 4356 57092 4360 57148
rect 4296 57088 4360 57092
rect 4376 57148 4440 57152
rect 4376 57092 4380 57148
rect 4380 57092 4436 57148
rect 4436 57092 4440 57148
rect 4376 57088 4440 57092
rect 4456 57148 4520 57152
rect 4456 57092 4460 57148
rect 4460 57092 4516 57148
rect 4516 57092 4520 57148
rect 4456 57088 4520 57092
rect 34936 57148 35000 57152
rect 34936 57092 34940 57148
rect 34940 57092 34996 57148
rect 34996 57092 35000 57148
rect 34936 57088 35000 57092
rect 35016 57148 35080 57152
rect 35016 57092 35020 57148
rect 35020 57092 35076 57148
rect 35076 57092 35080 57148
rect 35016 57088 35080 57092
rect 35096 57148 35160 57152
rect 35096 57092 35100 57148
rect 35100 57092 35156 57148
rect 35156 57092 35160 57148
rect 35096 57088 35160 57092
rect 35176 57148 35240 57152
rect 35176 57092 35180 57148
rect 35180 57092 35236 57148
rect 35236 57092 35240 57148
rect 35176 57088 35240 57092
rect 19576 56604 19640 56608
rect 19576 56548 19580 56604
rect 19580 56548 19636 56604
rect 19636 56548 19640 56604
rect 19576 56544 19640 56548
rect 19656 56604 19720 56608
rect 19656 56548 19660 56604
rect 19660 56548 19716 56604
rect 19716 56548 19720 56604
rect 19656 56544 19720 56548
rect 19736 56604 19800 56608
rect 19736 56548 19740 56604
rect 19740 56548 19796 56604
rect 19796 56548 19800 56604
rect 19736 56544 19800 56548
rect 19816 56604 19880 56608
rect 19816 56548 19820 56604
rect 19820 56548 19876 56604
rect 19876 56548 19880 56604
rect 19816 56544 19880 56548
rect 50296 56604 50360 56608
rect 50296 56548 50300 56604
rect 50300 56548 50356 56604
rect 50356 56548 50360 56604
rect 50296 56544 50360 56548
rect 50376 56604 50440 56608
rect 50376 56548 50380 56604
rect 50380 56548 50436 56604
rect 50436 56548 50440 56604
rect 50376 56544 50440 56548
rect 50456 56604 50520 56608
rect 50456 56548 50460 56604
rect 50460 56548 50516 56604
rect 50516 56548 50520 56604
rect 50456 56544 50520 56548
rect 50536 56604 50600 56608
rect 50536 56548 50540 56604
rect 50540 56548 50596 56604
rect 50596 56548 50600 56604
rect 50536 56544 50600 56548
rect 4216 56060 4280 56064
rect 4216 56004 4220 56060
rect 4220 56004 4276 56060
rect 4276 56004 4280 56060
rect 4216 56000 4280 56004
rect 4296 56060 4360 56064
rect 4296 56004 4300 56060
rect 4300 56004 4356 56060
rect 4356 56004 4360 56060
rect 4296 56000 4360 56004
rect 4376 56060 4440 56064
rect 4376 56004 4380 56060
rect 4380 56004 4436 56060
rect 4436 56004 4440 56060
rect 4376 56000 4440 56004
rect 4456 56060 4520 56064
rect 4456 56004 4460 56060
rect 4460 56004 4516 56060
rect 4516 56004 4520 56060
rect 4456 56000 4520 56004
rect 34936 56060 35000 56064
rect 34936 56004 34940 56060
rect 34940 56004 34996 56060
rect 34996 56004 35000 56060
rect 34936 56000 35000 56004
rect 35016 56060 35080 56064
rect 35016 56004 35020 56060
rect 35020 56004 35076 56060
rect 35076 56004 35080 56060
rect 35016 56000 35080 56004
rect 35096 56060 35160 56064
rect 35096 56004 35100 56060
rect 35100 56004 35156 56060
rect 35156 56004 35160 56060
rect 35096 56000 35160 56004
rect 35176 56060 35240 56064
rect 35176 56004 35180 56060
rect 35180 56004 35236 56060
rect 35236 56004 35240 56060
rect 35176 56000 35240 56004
rect 19576 55516 19640 55520
rect 19576 55460 19580 55516
rect 19580 55460 19636 55516
rect 19636 55460 19640 55516
rect 19576 55456 19640 55460
rect 19656 55516 19720 55520
rect 19656 55460 19660 55516
rect 19660 55460 19716 55516
rect 19716 55460 19720 55516
rect 19656 55456 19720 55460
rect 19736 55516 19800 55520
rect 19736 55460 19740 55516
rect 19740 55460 19796 55516
rect 19796 55460 19800 55516
rect 19736 55456 19800 55460
rect 19816 55516 19880 55520
rect 19816 55460 19820 55516
rect 19820 55460 19876 55516
rect 19876 55460 19880 55516
rect 19816 55456 19880 55460
rect 50296 55516 50360 55520
rect 50296 55460 50300 55516
rect 50300 55460 50356 55516
rect 50356 55460 50360 55516
rect 50296 55456 50360 55460
rect 50376 55516 50440 55520
rect 50376 55460 50380 55516
rect 50380 55460 50436 55516
rect 50436 55460 50440 55516
rect 50376 55456 50440 55460
rect 50456 55516 50520 55520
rect 50456 55460 50460 55516
rect 50460 55460 50516 55516
rect 50516 55460 50520 55516
rect 50456 55456 50520 55460
rect 50536 55516 50600 55520
rect 50536 55460 50540 55516
rect 50540 55460 50596 55516
rect 50596 55460 50600 55516
rect 50536 55456 50600 55460
rect 4216 54972 4280 54976
rect 4216 54916 4220 54972
rect 4220 54916 4276 54972
rect 4276 54916 4280 54972
rect 4216 54912 4280 54916
rect 4296 54972 4360 54976
rect 4296 54916 4300 54972
rect 4300 54916 4356 54972
rect 4356 54916 4360 54972
rect 4296 54912 4360 54916
rect 4376 54972 4440 54976
rect 4376 54916 4380 54972
rect 4380 54916 4436 54972
rect 4436 54916 4440 54972
rect 4376 54912 4440 54916
rect 4456 54972 4520 54976
rect 4456 54916 4460 54972
rect 4460 54916 4516 54972
rect 4516 54916 4520 54972
rect 4456 54912 4520 54916
rect 34936 54972 35000 54976
rect 34936 54916 34940 54972
rect 34940 54916 34996 54972
rect 34996 54916 35000 54972
rect 34936 54912 35000 54916
rect 35016 54972 35080 54976
rect 35016 54916 35020 54972
rect 35020 54916 35076 54972
rect 35076 54916 35080 54972
rect 35016 54912 35080 54916
rect 35096 54972 35160 54976
rect 35096 54916 35100 54972
rect 35100 54916 35156 54972
rect 35156 54916 35160 54972
rect 35096 54912 35160 54916
rect 35176 54972 35240 54976
rect 35176 54916 35180 54972
rect 35180 54916 35236 54972
rect 35236 54916 35240 54972
rect 35176 54912 35240 54916
rect 19576 54428 19640 54432
rect 19576 54372 19580 54428
rect 19580 54372 19636 54428
rect 19636 54372 19640 54428
rect 19576 54368 19640 54372
rect 19656 54428 19720 54432
rect 19656 54372 19660 54428
rect 19660 54372 19716 54428
rect 19716 54372 19720 54428
rect 19656 54368 19720 54372
rect 19736 54428 19800 54432
rect 19736 54372 19740 54428
rect 19740 54372 19796 54428
rect 19796 54372 19800 54428
rect 19736 54368 19800 54372
rect 19816 54428 19880 54432
rect 19816 54372 19820 54428
rect 19820 54372 19876 54428
rect 19876 54372 19880 54428
rect 19816 54368 19880 54372
rect 50296 54428 50360 54432
rect 50296 54372 50300 54428
rect 50300 54372 50356 54428
rect 50356 54372 50360 54428
rect 50296 54368 50360 54372
rect 50376 54428 50440 54432
rect 50376 54372 50380 54428
rect 50380 54372 50436 54428
rect 50436 54372 50440 54428
rect 50376 54368 50440 54372
rect 50456 54428 50520 54432
rect 50456 54372 50460 54428
rect 50460 54372 50516 54428
rect 50516 54372 50520 54428
rect 50456 54368 50520 54372
rect 50536 54428 50600 54432
rect 50536 54372 50540 54428
rect 50540 54372 50596 54428
rect 50596 54372 50600 54428
rect 50536 54368 50600 54372
rect 4216 53884 4280 53888
rect 4216 53828 4220 53884
rect 4220 53828 4276 53884
rect 4276 53828 4280 53884
rect 4216 53824 4280 53828
rect 4296 53884 4360 53888
rect 4296 53828 4300 53884
rect 4300 53828 4356 53884
rect 4356 53828 4360 53884
rect 4296 53824 4360 53828
rect 4376 53884 4440 53888
rect 4376 53828 4380 53884
rect 4380 53828 4436 53884
rect 4436 53828 4440 53884
rect 4376 53824 4440 53828
rect 4456 53884 4520 53888
rect 4456 53828 4460 53884
rect 4460 53828 4516 53884
rect 4516 53828 4520 53884
rect 4456 53824 4520 53828
rect 34936 53884 35000 53888
rect 34936 53828 34940 53884
rect 34940 53828 34996 53884
rect 34996 53828 35000 53884
rect 34936 53824 35000 53828
rect 35016 53884 35080 53888
rect 35016 53828 35020 53884
rect 35020 53828 35076 53884
rect 35076 53828 35080 53884
rect 35016 53824 35080 53828
rect 35096 53884 35160 53888
rect 35096 53828 35100 53884
rect 35100 53828 35156 53884
rect 35156 53828 35160 53884
rect 35096 53824 35160 53828
rect 35176 53884 35240 53888
rect 35176 53828 35180 53884
rect 35180 53828 35236 53884
rect 35236 53828 35240 53884
rect 35176 53824 35240 53828
rect 19576 53340 19640 53344
rect 19576 53284 19580 53340
rect 19580 53284 19636 53340
rect 19636 53284 19640 53340
rect 19576 53280 19640 53284
rect 19656 53340 19720 53344
rect 19656 53284 19660 53340
rect 19660 53284 19716 53340
rect 19716 53284 19720 53340
rect 19656 53280 19720 53284
rect 19736 53340 19800 53344
rect 19736 53284 19740 53340
rect 19740 53284 19796 53340
rect 19796 53284 19800 53340
rect 19736 53280 19800 53284
rect 19816 53340 19880 53344
rect 19816 53284 19820 53340
rect 19820 53284 19876 53340
rect 19876 53284 19880 53340
rect 19816 53280 19880 53284
rect 50296 53340 50360 53344
rect 50296 53284 50300 53340
rect 50300 53284 50356 53340
rect 50356 53284 50360 53340
rect 50296 53280 50360 53284
rect 50376 53340 50440 53344
rect 50376 53284 50380 53340
rect 50380 53284 50436 53340
rect 50436 53284 50440 53340
rect 50376 53280 50440 53284
rect 50456 53340 50520 53344
rect 50456 53284 50460 53340
rect 50460 53284 50516 53340
rect 50516 53284 50520 53340
rect 50456 53280 50520 53284
rect 50536 53340 50600 53344
rect 50536 53284 50540 53340
rect 50540 53284 50596 53340
rect 50596 53284 50600 53340
rect 50536 53280 50600 53284
rect 4216 52796 4280 52800
rect 4216 52740 4220 52796
rect 4220 52740 4276 52796
rect 4276 52740 4280 52796
rect 4216 52736 4280 52740
rect 4296 52796 4360 52800
rect 4296 52740 4300 52796
rect 4300 52740 4356 52796
rect 4356 52740 4360 52796
rect 4296 52736 4360 52740
rect 4376 52796 4440 52800
rect 4376 52740 4380 52796
rect 4380 52740 4436 52796
rect 4436 52740 4440 52796
rect 4376 52736 4440 52740
rect 4456 52796 4520 52800
rect 4456 52740 4460 52796
rect 4460 52740 4516 52796
rect 4516 52740 4520 52796
rect 4456 52736 4520 52740
rect 34936 52796 35000 52800
rect 34936 52740 34940 52796
rect 34940 52740 34996 52796
rect 34996 52740 35000 52796
rect 34936 52736 35000 52740
rect 35016 52796 35080 52800
rect 35016 52740 35020 52796
rect 35020 52740 35076 52796
rect 35076 52740 35080 52796
rect 35016 52736 35080 52740
rect 35096 52796 35160 52800
rect 35096 52740 35100 52796
rect 35100 52740 35156 52796
rect 35156 52740 35160 52796
rect 35096 52736 35160 52740
rect 35176 52796 35240 52800
rect 35176 52740 35180 52796
rect 35180 52740 35236 52796
rect 35236 52740 35240 52796
rect 35176 52736 35240 52740
rect 19576 52252 19640 52256
rect 19576 52196 19580 52252
rect 19580 52196 19636 52252
rect 19636 52196 19640 52252
rect 19576 52192 19640 52196
rect 19656 52252 19720 52256
rect 19656 52196 19660 52252
rect 19660 52196 19716 52252
rect 19716 52196 19720 52252
rect 19656 52192 19720 52196
rect 19736 52252 19800 52256
rect 19736 52196 19740 52252
rect 19740 52196 19796 52252
rect 19796 52196 19800 52252
rect 19736 52192 19800 52196
rect 19816 52252 19880 52256
rect 19816 52196 19820 52252
rect 19820 52196 19876 52252
rect 19876 52196 19880 52252
rect 19816 52192 19880 52196
rect 50296 52252 50360 52256
rect 50296 52196 50300 52252
rect 50300 52196 50356 52252
rect 50356 52196 50360 52252
rect 50296 52192 50360 52196
rect 50376 52252 50440 52256
rect 50376 52196 50380 52252
rect 50380 52196 50436 52252
rect 50436 52196 50440 52252
rect 50376 52192 50440 52196
rect 50456 52252 50520 52256
rect 50456 52196 50460 52252
rect 50460 52196 50516 52252
rect 50516 52196 50520 52252
rect 50456 52192 50520 52196
rect 50536 52252 50600 52256
rect 50536 52196 50540 52252
rect 50540 52196 50596 52252
rect 50596 52196 50600 52252
rect 50536 52192 50600 52196
rect 4216 51708 4280 51712
rect 4216 51652 4220 51708
rect 4220 51652 4276 51708
rect 4276 51652 4280 51708
rect 4216 51648 4280 51652
rect 4296 51708 4360 51712
rect 4296 51652 4300 51708
rect 4300 51652 4356 51708
rect 4356 51652 4360 51708
rect 4296 51648 4360 51652
rect 4376 51708 4440 51712
rect 4376 51652 4380 51708
rect 4380 51652 4436 51708
rect 4436 51652 4440 51708
rect 4376 51648 4440 51652
rect 4456 51708 4520 51712
rect 4456 51652 4460 51708
rect 4460 51652 4516 51708
rect 4516 51652 4520 51708
rect 4456 51648 4520 51652
rect 34936 51708 35000 51712
rect 34936 51652 34940 51708
rect 34940 51652 34996 51708
rect 34996 51652 35000 51708
rect 34936 51648 35000 51652
rect 35016 51708 35080 51712
rect 35016 51652 35020 51708
rect 35020 51652 35076 51708
rect 35076 51652 35080 51708
rect 35016 51648 35080 51652
rect 35096 51708 35160 51712
rect 35096 51652 35100 51708
rect 35100 51652 35156 51708
rect 35156 51652 35160 51708
rect 35096 51648 35160 51652
rect 35176 51708 35240 51712
rect 35176 51652 35180 51708
rect 35180 51652 35236 51708
rect 35236 51652 35240 51708
rect 35176 51648 35240 51652
rect 19576 51164 19640 51168
rect 19576 51108 19580 51164
rect 19580 51108 19636 51164
rect 19636 51108 19640 51164
rect 19576 51104 19640 51108
rect 19656 51164 19720 51168
rect 19656 51108 19660 51164
rect 19660 51108 19716 51164
rect 19716 51108 19720 51164
rect 19656 51104 19720 51108
rect 19736 51164 19800 51168
rect 19736 51108 19740 51164
rect 19740 51108 19796 51164
rect 19796 51108 19800 51164
rect 19736 51104 19800 51108
rect 19816 51164 19880 51168
rect 19816 51108 19820 51164
rect 19820 51108 19876 51164
rect 19876 51108 19880 51164
rect 19816 51104 19880 51108
rect 50296 51164 50360 51168
rect 50296 51108 50300 51164
rect 50300 51108 50356 51164
rect 50356 51108 50360 51164
rect 50296 51104 50360 51108
rect 50376 51164 50440 51168
rect 50376 51108 50380 51164
rect 50380 51108 50436 51164
rect 50436 51108 50440 51164
rect 50376 51104 50440 51108
rect 50456 51164 50520 51168
rect 50456 51108 50460 51164
rect 50460 51108 50516 51164
rect 50516 51108 50520 51164
rect 50456 51104 50520 51108
rect 50536 51164 50600 51168
rect 50536 51108 50540 51164
rect 50540 51108 50596 51164
rect 50596 51108 50600 51164
rect 50536 51104 50600 51108
rect 4216 50620 4280 50624
rect 4216 50564 4220 50620
rect 4220 50564 4276 50620
rect 4276 50564 4280 50620
rect 4216 50560 4280 50564
rect 4296 50620 4360 50624
rect 4296 50564 4300 50620
rect 4300 50564 4356 50620
rect 4356 50564 4360 50620
rect 4296 50560 4360 50564
rect 4376 50620 4440 50624
rect 4376 50564 4380 50620
rect 4380 50564 4436 50620
rect 4436 50564 4440 50620
rect 4376 50560 4440 50564
rect 4456 50620 4520 50624
rect 4456 50564 4460 50620
rect 4460 50564 4516 50620
rect 4516 50564 4520 50620
rect 4456 50560 4520 50564
rect 34936 50620 35000 50624
rect 34936 50564 34940 50620
rect 34940 50564 34996 50620
rect 34996 50564 35000 50620
rect 34936 50560 35000 50564
rect 35016 50620 35080 50624
rect 35016 50564 35020 50620
rect 35020 50564 35076 50620
rect 35076 50564 35080 50620
rect 35016 50560 35080 50564
rect 35096 50620 35160 50624
rect 35096 50564 35100 50620
rect 35100 50564 35156 50620
rect 35156 50564 35160 50620
rect 35096 50560 35160 50564
rect 35176 50620 35240 50624
rect 35176 50564 35180 50620
rect 35180 50564 35236 50620
rect 35236 50564 35240 50620
rect 35176 50560 35240 50564
rect 19576 50076 19640 50080
rect 19576 50020 19580 50076
rect 19580 50020 19636 50076
rect 19636 50020 19640 50076
rect 19576 50016 19640 50020
rect 19656 50076 19720 50080
rect 19656 50020 19660 50076
rect 19660 50020 19716 50076
rect 19716 50020 19720 50076
rect 19656 50016 19720 50020
rect 19736 50076 19800 50080
rect 19736 50020 19740 50076
rect 19740 50020 19796 50076
rect 19796 50020 19800 50076
rect 19736 50016 19800 50020
rect 19816 50076 19880 50080
rect 19816 50020 19820 50076
rect 19820 50020 19876 50076
rect 19876 50020 19880 50076
rect 19816 50016 19880 50020
rect 50296 50076 50360 50080
rect 50296 50020 50300 50076
rect 50300 50020 50356 50076
rect 50356 50020 50360 50076
rect 50296 50016 50360 50020
rect 50376 50076 50440 50080
rect 50376 50020 50380 50076
rect 50380 50020 50436 50076
rect 50436 50020 50440 50076
rect 50376 50016 50440 50020
rect 50456 50076 50520 50080
rect 50456 50020 50460 50076
rect 50460 50020 50516 50076
rect 50516 50020 50520 50076
rect 50456 50016 50520 50020
rect 50536 50076 50600 50080
rect 50536 50020 50540 50076
rect 50540 50020 50596 50076
rect 50596 50020 50600 50076
rect 50536 50016 50600 50020
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 50296 48988 50360 48992
rect 50296 48932 50300 48988
rect 50300 48932 50356 48988
rect 50356 48932 50360 48988
rect 50296 48928 50360 48932
rect 50376 48988 50440 48992
rect 50376 48932 50380 48988
rect 50380 48932 50436 48988
rect 50436 48932 50440 48988
rect 50376 48928 50440 48932
rect 50456 48988 50520 48992
rect 50456 48932 50460 48988
rect 50460 48932 50516 48988
rect 50516 48932 50520 48988
rect 50456 48928 50520 48932
rect 50536 48988 50600 48992
rect 50536 48932 50540 48988
rect 50540 48932 50596 48988
rect 50596 48932 50600 48988
rect 50536 48928 50600 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 50296 47900 50360 47904
rect 50296 47844 50300 47900
rect 50300 47844 50356 47900
rect 50356 47844 50360 47900
rect 50296 47840 50360 47844
rect 50376 47900 50440 47904
rect 50376 47844 50380 47900
rect 50380 47844 50436 47900
rect 50436 47844 50440 47900
rect 50376 47840 50440 47844
rect 50456 47900 50520 47904
rect 50456 47844 50460 47900
rect 50460 47844 50516 47900
rect 50516 47844 50520 47900
rect 50456 47840 50520 47844
rect 50536 47900 50600 47904
rect 50536 47844 50540 47900
rect 50540 47844 50596 47900
rect 50596 47844 50600 47900
rect 50536 47840 50600 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 50296 46812 50360 46816
rect 50296 46756 50300 46812
rect 50300 46756 50356 46812
rect 50356 46756 50360 46812
rect 50296 46752 50360 46756
rect 50376 46812 50440 46816
rect 50376 46756 50380 46812
rect 50380 46756 50436 46812
rect 50436 46756 50440 46812
rect 50376 46752 50440 46756
rect 50456 46812 50520 46816
rect 50456 46756 50460 46812
rect 50460 46756 50516 46812
rect 50516 46756 50520 46812
rect 50456 46752 50520 46756
rect 50536 46812 50600 46816
rect 50536 46756 50540 46812
rect 50540 46756 50596 46812
rect 50596 46756 50600 46812
rect 50536 46752 50600 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 50296 45724 50360 45728
rect 50296 45668 50300 45724
rect 50300 45668 50356 45724
rect 50356 45668 50360 45724
rect 50296 45664 50360 45668
rect 50376 45724 50440 45728
rect 50376 45668 50380 45724
rect 50380 45668 50436 45724
rect 50436 45668 50440 45724
rect 50376 45664 50440 45668
rect 50456 45724 50520 45728
rect 50456 45668 50460 45724
rect 50460 45668 50516 45724
rect 50516 45668 50520 45724
rect 50456 45664 50520 45668
rect 50536 45724 50600 45728
rect 50536 45668 50540 45724
rect 50540 45668 50596 45724
rect 50596 45668 50600 45724
rect 50536 45664 50600 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 50296 44636 50360 44640
rect 50296 44580 50300 44636
rect 50300 44580 50356 44636
rect 50356 44580 50360 44636
rect 50296 44576 50360 44580
rect 50376 44636 50440 44640
rect 50376 44580 50380 44636
rect 50380 44580 50436 44636
rect 50436 44580 50440 44636
rect 50376 44576 50440 44580
rect 50456 44636 50520 44640
rect 50456 44580 50460 44636
rect 50460 44580 50516 44636
rect 50516 44580 50520 44636
rect 50456 44576 50520 44580
rect 50536 44636 50600 44640
rect 50536 44580 50540 44636
rect 50540 44580 50596 44636
rect 50596 44580 50600 44636
rect 50536 44576 50600 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 50296 43548 50360 43552
rect 50296 43492 50300 43548
rect 50300 43492 50356 43548
rect 50356 43492 50360 43548
rect 50296 43488 50360 43492
rect 50376 43548 50440 43552
rect 50376 43492 50380 43548
rect 50380 43492 50436 43548
rect 50436 43492 50440 43548
rect 50376 43488 50440 43492
rect 50456 43548 50520 43552
rect 50456 43492 50460 43548
rect 50460 43492 50516 43548
rect 50516 43492 50520 43548
rect 50456 43488 50520 43492
rect 50536 43548 50600 43552
rect 50536 43492 50540 43548
rect 50540 43492 50596 43548
rect 50596 43492 50600 43548
rect 50536 43488 50600 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 50296 42460 50360 42464
rect 50296 42404 50300 42460
rect 50300 42404 50356 42460
rect 50356 42404 50360 42460
rect 50296 42400 50360 42404
rect 50376 42460 50440 42464
rect 50376 42404 50380 42460
rect 50380 42404 50436 42460
rect 50436 42404 50440 42460
rect 50376 42400 50440 42404
rect 50456 42460 50520 42464
rect 50456 42404 50460 42460
rect 50460 42404 50516 42460
rect 50516 42404 50520 42460
rect 50456 42400 50520 42404
rect 50536 42460 50600 42464
rect 50536 42404 50540 42460
rect 50540 42404 50596 42460
rect 50596 42404 50600 42460
rect 50536 42400 50600 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 50296 41372 50360 41376
rect 50296 41316 50300 41372
rect 50300 41316 50356 41372
rect 50356 41316 50360 41372
rect 50296 41312 50360 41316
rect 50376 41372 50440 41376
rect 50376 41316 50380 41372
rect 50380 41316 50436 41372
rect 50436 41316 50440 41372
rect 50376 41312 50440 41316
rect 50456 41372 50520 41376
rect 50456 41316 50460 41372
rect 50460 41316 50516 41372
rect 50516 41316 50520 41372
rect 50456 41312 50520 41316
rect 50536 41372 50600 41376
rect 50536 41316 50540 41372
rect 50540 41316 50596 41372
rect 50596 41316 50600 41372
rect 50536 41312 50600 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 50296 40284 50360 40288
rect 50296 40228 50300 40284
rect 50300 40228 50356 40284
rect 50356 40228 50360 40284
rect 50296 40224 50360 40228
rect 50376 40284 50440 40288
rect 50376 40228 50380 40284
rect 50380 40228 50436 40284
rect 50436 40228 50440 40284
rect 50376 40224 50440 40228
rect 50456 40284 50520 40288
rect 50456 40228 50460 40284
rect 50460 40228 50516 40284
rect 50516 40228 50520 40284
rect 50456 40224 50520 40228
rect 50536 40284 50600 40288
rect 50536 40228 50540 40284
rect 50540 40228 50596 40284
rect 50596 40228 50600 40284
rect 50536 40224 50600 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 50296 39196 50360 39200
rect 50296 39140 50300 39196
rect 50300 39140 50356 39196
rect 50356 39140 50360 39196
rect 50296 39136 50360 39140
rect 50376 39196 50440 39200
rect 50376 39140 50380 39196
rect 50380 39140 50436 39196
rect 50436 39140 50440 39196
rect 50376 39136 50440 39140
rect 50456 39196 50520 39200
rect 50456 39140 50460 39196
rect 50460 39140 50516 39196
rect 50516 39140 50520 39196
rect 50456 39136 50520 39140
rect 50536 39196 50600 39200
rect 50536 39140 50540 39196
rect 50540 39140 50596 39196
rect 50596 39140 50600 39196
rect 50536 39136 50600 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 50296 38108 50360 38112
rect 50296 38052 50300 38108
rect 50300 38052 50356 38108
rect 50356 38052 50360 38108
rect 50296 38048 50360 38052
rect 50376 38108 50440 38112
rect 50376 38052 50380 38108
rect 50380 38052 50436 38108
rect 50436 38052 50440 38108
rect 50376 38048 50440 38052
rect 50456 38108 50520 38112
rect 50456 38052 50460 38108
rect 50460 38052 50516 38108
rect 50516 38052 50520 38108
rect 50456 38048 50520 38052
rect 50536 38108 50600 38112
rect 50536 38052 50540 38108
rect 50540 38052 50596 38108
rect 50596 38052 50600 38108
rect 50536 38048 50600 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 51212 29140 51276 29204
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 50108 27704 50172 27708
rect 50108 27648 50122 27704
rect 50122 27648 50172 27704
rect 50108 27644 50172 27648
rect 51212 27508 51276 27572
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 49740 25664 49804 25668
rect 49740 25608 49790 25664
rect 49790 25608 49804 25664
rect 49740 25604 49804 25608
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 50108 20436 50172 20500
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 49740 18396 49804 18460
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 57152 4528 57712
rect 4208 57088 4216 57152
rect 4280 57088 4296 57152
rect 4360 57088 4376 57152
rect 4440 57088 4456 57152
rect 4520 57088 4528 57152
rect 4208 56064 4528 57088
rect 4208 56000 4216 56064
rect 4280 56000 4296 56064
rect 4360 56000 4376 56064
rect 4440 56000 4456 56064
rect 4520 56000 4528 56064
rect 4208 54976 4528 56000
rect 4208 54912 4216 54976
rect 4280 54912 4296 54976
rect 4360 54912 4376 54976
rect 4440 54912 4456 54976
rect 4520 54912 4528 54976
rect 4208 53888 4528 54912
rect 4208 53824 4216 53888
rect 4280 53824 4296 53888
rect 4360 53824 4376 53888
rect 4440 53824 4456 53888
rect 4520 53824 4528 53888
rect 4208 52800 4528 53824
rect 4208 52736 4216 52800
rect 4280 52736 4296 52800
rect 4360 52736 4376 52800
rect 4440 52736 4456 52800
rect 4520 52736 4528 52800
rect 4208 51712 4528 52736
rect 4208 51648 4216 51712
rect 4280 51648 4296 51712
rect 4360 51648 4376 51712
rect 4440 51648 4456 51712
rect 4520 51648 4528 51712
rect 4208 50624 4528 51648
rect 4208 50560 4216 50624
rect 4280 50560 4296 50624
rect 4360 50560 4376 50624
rect 4440 50560 4456 50624
rect 4520 50560 4528 50624
rect 4208 49536 4528 50560
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 57696 19888 57712
rect 19568 57632 19576 57696
rect 19640 57632 19656 57696
rect 19720 57632 19736 57696
rect 19800 57632 19816 57696
rect 19880 57632 19888 57696
rect 19568 56608 19888 57632
rect 19568 56544 19576 56608
rect 19640 56544 19656 56608
rect 19720 56544 19736 56608
rect 19800 56544 19816 56608
rect 19880 56544 19888 56608
rect 19568 55520 19888 56544
rect 19568 55456 19576 55520
rect 19640 55456 19656 55520
rect 19720 55456 19736 55520
rect 19800 55456 19816 55520
rect 19880 55456 19888 55520
rect 19568 54432 19888 55456
rect 19568 54368 19576 54432
rect 19640 54368 19656 54432
rect 19720 54368 19736 54432
rect 19800 54368 19816 54432
rect 19880 54368 19888 54432
rect 19568 53344 19888 54368
rect 19568 53280 19576 53344
rect 19640 53280 19656 53344
rect 19720 53280 19736 53344
rect 19800 53280 19816 53344
rect 19880 53280 19888 53344
rect 19568 52256 19888 53280
rect 19568 52192 19576 52256
rect 19640 52192 19656 52256
rect 19720 52192 19736 52256
rect 19800 52192 19816 52256
rect 19880 52192 19888 52256
rect 19568 51168 19888 52192
rect 19568 51104 19576 51168
rect 19640 51104 19656 51168
rect 19720 51104 19736 51168
rect 19800 51104 19816 51168
rect 19880 51104 19888 51168
rect 19568 50080 19888 51104
rect 19568 50016 19576 50080
rect 19640 50016 19656 50080
rect 19720 50016 19736 50080
rect 19800 50016 19816 50080
rect 19880 50016 19888 50080
rect 19568 48992 19888 50016
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 57152 35248 57712
rect 34928 57088 34936 57152
rect 35000 57088 35016 57152
rect 35080 57088 35096 57152
rect 35160 57088 35176 57152
rect 35240 57088 35248 57152
rect 34928 56064 35248 57088
rect 34928 56000 34936 56064
rect 35000 56000 35016 56064
rect 35080 56000 35096 56064
rect 35160 56000 35176 56064
rect 35240 56000 35248 56064
rect 34928 54976 35248 56000
rect 34928 54912 34936 54976
rect 35000 54912 35016 54976
rect 35080 54912 35096 54976
rect 35160 54912 35176 54976
rect 35240 54912 35248 54976
rect 34928 53888 35248 54912
rect 34928 53824 34936 53888
rect 35000 53824 35016 53888
rect 35080 53824 35096 53888
rect 35160 53824 35176 53888
rect 35240 53824 35248 53888
rect 34928 52800 35248 53824
rect 34928 52736 34936 52800
rect 35000 52736 35016 52800
rect 35080 52736 35096 52800
rect 35160 52736 35176 52800
rect 35240 52736 35248 52800
rect 34928 51712 35248 52736
rect 34928 51648 34936 51712
rect 35000 51648 35016 51712
rect 35080 51648 35096 51712
rect 35160 51648 35176 51712
rect 35240 51648 35248 51712
rect 34928 50624 35248 51648
rect 34928 50560 34936 50624
rect 35000 50560 35016 50624
rect 35080 50560 35096 50624
rect 35160 50560 35176 50624
rect 35240 50560 35248 50624
rect 34928 49536 35248 50560
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 50288 57696 50608 57712
rect 50288 57632 50296 57696
rect 50360 57632 50376 57696
rect 50440 57632 50456 57696
rect 50520 57632 50536 57696
rect 50600 57632 50608 57696
rect 50288 56608 50608 57632
rect 50288 56544 50296 56608
rect 50360 56544 50376 56608
rect 50440 56544 50456 56608
rect 50520 56544 50536 56608
rect 50600 56544 50608 56608
rect 50288 55520 50608 56544
rect 50288 55456 50296 55520
rect 50360 55456 50376 55520
rect 50440 55456 50456 55520
rect 50520 55456 50536 55520
rect 50600 55456 50608 55520
rect 50288 54432 50608 55456
rect 50288 54368 50296 54432
rect 50360 54368 50376 54432
rect 50440 54368 50456 54432
rect 50520 54368 50536 54432
rect 50600 54368 50608 54432
rect 50288 53344 50608 54368
rect 50288 53280 50296 53344
rect 50360 53280 50376 53344
rect 50440 53280 50456 53344
rect 50520 53280 50536 53344
rect 50600 53280 50608 53344
rect 50288 52256 50608 53280
rect 50288 52192 50296 52256
rect 50360 52192 50376 52256
rect 50440 52192 50456 52256
rect 50520 52192 50536 52256
rect 50600 52192 50608 52256
rect 50288 51168 50608 52192
rect 50288 51104 50296 51168
rect 50360 51104 50376 51168
rect 50440 51104 50456 51168
rect 50520 51104 50536 51168
rect 50600 51104 50608 51168
rect 50288 50080 50608 51104
rect 50288 50016 50296 50080
rect 50360 50016 50376 50080
rect 50440 50016 50456 50080
rect 50520 50016 50536 50080
rect 50600 50016 50608 50080
rect 50288 48992 50608 50016
rect 50288 48928 50296 48992
rect 50360 48928 50376 48992
rect 50440 48928 50456 48992
rect 50520 48928 50536 48992
rect 50600 48928 50608 48992
rect 50288 47904 50608 48928
rect 50288 47840 50296 47904
rect 50360 47840 50376 47904
rect 50440 47840 50456 47904
rect 50520 47840 50536 47904
rect 50600 47840 50608 47904
rect 50288 46816 50608 47840
rect 50288 46752 50296 46816
rect 50360 46752 50376 46816
rect 50440 46752 50456 46816
rect 50520 46752 50536 46816
rect 50600 46752 50608 46816
rect 50288 45728 50608 46752
rect 50288 45664 50296 45728
rect 50360 45664 50376 45728
rect 50440 45664 50456 45728
rect 50520 45664 50536 45728
rect 50600 45664 50608 45728
rect 50288 44640 50608 45664
rect 50288 44576 50296 44640
rect 50360 44576 50376 44640
rect 50440 44576 50456 44640
rect 50520 44576 50536 44640
rect 50600 44576 50608 44640
rect 50288 43552 50608 44576
rect 50288 43488 50296 43552
rect 50360 43488 50376 43552
rect 50440 43488 50456 43552
rect 50520 43488 50536 43552
rect 50600 43488 50608 43552
rect 50288 42464 50608 43488
rect 50288 42400 50296 42464
rect 50360 42400 50376 42464
rect 50440 42400 50456 42464
rect 50520 42400 50536 42464
rect 50600 42400 50608 42464
rect 50288 41376 50608 42400
rect 50288 41312 50296 41376
rect 50360 41312 50376 41376
rect 50440 41312 50456 41376
rect 50520 41312 50536 41376
rect 50600 41312 50608 41376
rect 50288 40288 50608 41312
rect 50288 40224 50296 40288
rect 50360 40224 50376 40288
rect 50440 40224 50456 40288
rect 50520 40224 50536 40288
rect 50600 40224 50608 40288
rect 50288 39200 50608 40224
rect 50288 39136 50296 39200
rect 50360 39136 50376 39200
rect 50440 39136 50456 39200
rect 50520 39136 50536 39200
rect 50600 39136 50608 39200
rect 50288 38112 50608 39136
rect 50288 38048 50296 38112
rect 50360 38048 50376 38112
rect 50440 38048 50456 38112
rect 50520 38048 50536 38112
rect 50600 38048 50608 38112
rect 50288 37024 50608 38048
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 51211 29204 51277 29205
rect 51211 29140 51212 29204
rect 51276 29140 51277 29204
rect 51211 29139 51277 29140
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50107 27708 50173 27709
rect 50107 27644 50108 27708
rect 50172 27644 50173 27708
rect 50107 27643 50173 27644
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 49739 25668 49805 25669
rect 49739 25604 49740 25668
rect 49804 25604 49805 25668
rect 49739 25603 49805 25604
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 49742 18461 49802 25603
rect 50110 20501 50170 27643
rect 50288 27232 50608 28256
rect 51214 27573 51274 29139
rect 51211 27572 51277 27573
rect 51211 27508 51212 27572
rect 51276 27508 51277 27572
rect 51211 27507 51277 27508
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50107 20500 50173 20501
rect 50107 20436 50108 20500
rect 50172 20436 50173 20500
rect 50107 20435 50173 20436
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 49739 18460 49805 18461
rect 49739 18396 49740 18460
rect 49804 18396 49805 18460
rect 49739 18395 49805 18396
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__nand2_1  _0779_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11132 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0780_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12236 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0781_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12512 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0782_
timestamp 1688980957
transform -1 0 13064 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0783_
timestamp 1688980957
transform 1 0 12512 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0784_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 42320 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _0785_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12604 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0786_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0787_
timestamp 1688980957
transform -1 0 10856 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1688980957
transform -1 0 10212 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1688980957
transform -1 0 9016 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0790_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 8832 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0791_
timestamp 1688980957
transform 1 0 7820 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0792_
timestamp 1688980957
transform -1 0 8556 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1688980957
transform -1 0 9200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0794_
timestamp 1688980957
transform -1 0 8832 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0795_
timestamp 1688980957
transform 1 0 6992 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0796_
timestamp 1688980957
transform -1 0 8004 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0797_
timestamp 1688980957
transform -1 0 11868 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0798_
timestamp 1688980957
transform 1 0 9844 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0799_
timestamp 1688980957
transform -1 0 10396 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0800_
timestamp 1688980957
transform -1 0 10488 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1688980957
transform -1 0 12328 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _0802_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9568 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _0803_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 9476 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0804_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 5336 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0805_
timestamp 1688980957
transform 1 0 4600 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0806_
timestamp 1688980957
transform 1 0 4508 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0807_
timestamp 1688980957
transform -1 0 6808 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0808_
timestamp 1688980957
transform 1 0 5612 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0809_
timestamp 1688980957
transform -1 0 6716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0810_
timestamp 1688980957
transform -1 0 5060 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0811_
timestamp 1688980957
transform 1 0 4508 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0812_
timestamp 1688980957
transform 1 0 4508 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0813_
timestamp 1688980957
transform -1 0 8740 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0814_
timestamp 1688980957
transform 1 0 7912 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0815_
timestamp 1688980957
transform 1 0 7912 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0816_
timestamp 1688980957
transform 1 0 11224 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _0817_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11776 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _0818_
timestamp 1688980957
transform -1 0 5336 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0819_
timestamp 1688980957
transform 1 0 5428 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0820_
timestamp 1688980957
transform 1 0 5060 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0821_
timestamp 1688980957
transform 1 0 8556 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0822_
timestamp 1688980957
transform -1 0 10028 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0823_
timestamp 1688980957
transform 1 0 9108 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0824_
timestamp 1688980957
transform -1 0 8556 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0825_
timestamp 1688980957
transform 1 0 6992 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0826_
timestamp 1688980957
transform -1 0 7820 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _0827_
timestamp 1688980957
transform -1 0 9660 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0828_
timestamp 1688980957
transform -1 0 6624 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0829_
timestamp 1688980957
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _0830_
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _0831_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10396 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0832_
timestamp 1688980957
transform 1 0 9936 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0833_
timestamp 1688980957
transform 1 0 9660 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0834_
timestamp 1688980957
transform -1 0 10488 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0835_
timestamp 1688980957
transform 1 0 6072 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0836_
timestamp 1688980957
transform -1 0 7176 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0837_
timestamp 1688980957
transform 1 0 6532 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0838_
timestamp 1688980957
transform -1 0 5060 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0839_
timestamp 1688980957
transform 1 0 4140 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0840_
timestamp 1688980957
transform -1 0 4876 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _0841_
timestamp 1688980957
transform 1 0 10212 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0842_
timestamp 1688980957
transform 1 0 10580 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0843_
timestamp 1688980957
transform -1 0 12512 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0844_
timestamp 1688980957
transform -1 0 11224 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0845_
timestamp 1688980957
transform 1 0 46736 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0846_
timestamp 1688980957
transform 1 0 57868 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0847_
timestamp 1688980957
transform 1 0 58052 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _0848_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 57868 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _0849_
timestamp 1688980957
transform 1 0 57868 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0850_
timestamp 1688980957
transform 1 0 58236 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _0851_
timestamp 1688980957
transform -1 0 58420 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _0852_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 57868 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_2  _0853_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 58420 0 1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0854_
timestamp 1688980957
transform 1 0 47012 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0855_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 45632 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0856_
timestamp 1688980957
transform 1 0 47932 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0857_
timestamp 1688980957
transform -1 0 50416 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0858_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 50048 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _0859_
timestamp 1688980957
transform 1 0 49312 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _0860_
timestamp 1688980957
transform -1 0 48208 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0861_
timestamp 1688980957
transform -1 0 47840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _0862_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 50968 0 -1 26112
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2_1  _0863_
timestamp 1688980957
transform -1 0 47472 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3_2  _0864_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 47196 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1688980957
transform -1 0 44712 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0866_
timestamp 1688980957
transform 1 0 43332 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _0867_
timestamp 1688980957
transform 1 0 36800 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1688980957
transform 1 0 37904 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0869_
timestamp 1688980957
transform 1 0 39192 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0870_
timestamp 1688980957
transform -1 0 40020 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1688980957
transform 1 0 40388 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0872_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 41216 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1688980957
transform -1 0 48024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0874_
timestamp 1688980957
transform 1 0 47196 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0875_
timestamp 1688980957
transform -1 0 46368 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _0876_
timestamp 1688980957
transform -1 0 46276 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _0877_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44988 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_8  _0878_
timestamp 1688980957
transform 1 0 24564 0 1 27200
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2_1  _0879_
timestamp 1688980957
transform 1 0 46092 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0880_
timestamp 1688980957
transform -1 0 46644 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0881_
timestamp 1688980957
transform 1 0 47748 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0882_
timestamp 1688980957
transform 1 0 47104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0883_
timestamp 1688980957
transform 1 0 46736 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _0884_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 46460 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _0885_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 43516 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _0886_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 41768 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0887_
timestamp 1688980957
transform -1 0 15548 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0888_
timestamp 1688980957
transform -1 0 38916 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1688980957
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0890_
timestamp 1688980957
transform -1 0 39284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1688980957
transform 1 0 12880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0892_
timestamp 1688980957
transform -1 0 39468 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1688980957
transform 1 0 39468 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0894_
timestamp 1688980957
transform -1 0 39468 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1688980957
transform -1 0 41400 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0896_
timestamp 1688980957
transform -1 0 41216 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__buf_8  _0897_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _0898_
timestamp 1688980957
transform 1 0 37720 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0899_
timestamp 1688980957
transform 1 0 37352 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0900_
timestamp 1688980957
transform 1 0 50784 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _0901_
timestamp 1688980957
transform 1 0 52716 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1688980957
transform 1 0 49128 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0903_
timestamp 1688980957
transform -1 0 51704 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1688980957
transform -1 0 50048 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0905_
timestamp 1688980957
transform -1 0 49128 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0906_
timestamp 1688980957
transform -1 0 49128 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0907_
timestamp 1688980957
transform 1 0 48576 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1688980957
transform -1 0 49680 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0909_
timestamp 1688980957
transform -1 0 41400 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1688980957
transform 1 0 39836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0911_
timestamp 1688980957
transform -1 0 39744 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0912_
timestamp 1688980957
transform -1 0 39100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0913_
timestamp 1688980957
transform 1 0 38732 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1688980957
transform -1 0 39284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0915_
timestamp 1688980957
transform -1 0 39192 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1688980957
transform -1 0 40112 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0917_
timestamp 1688980957
transform -1 0 39744 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1688980957
transform 1 0 40388 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _0919_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 40204 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0920_
timestamp 1688980957
transform 1 0 43976 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_1  _0921_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _0922_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 47840 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1688980957
transform 1 0 42964 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1688980957
transform -1 0 43792 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  _0925_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44436 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _0926_
timestamp 1688980957
transform -1 0 45724 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_2  _0927_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42780 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1688980957
transform 1 0 44160 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_2  _0929_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 44068 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _0930_
timestamp 1688980957
transform -1 0 40204 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _0931_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 43700 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _0932_
timestamp 1688980957
transform -1 0 44160 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _0933_
timestamp 1688980957
transform 1 0 43700 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1688980957
transform 1 0 44252 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _0935_
timestamp 1688980957
transform 1 0 44528 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _0936_
timestamp 1688980957
transform 1 0 51428 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _0937_
timestamp 1688980957
transform -1 0 51428 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _0938_
timestamp 1688980957
transform -1 0 45816 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _0939_
timestamp 1688980957
transform -1 0 46368 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0940_
timestamp 1688980957
transform -1 0 43976 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _0941_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 41400 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 40296 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0943_
timestamp 1688980957
transform 1 0 47196 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0944_
timestamp 1688980957
transform 1 0 47288 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _0945_
timestamp 1688980957
transform 1 0 45632 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0946_
timestamp 1688980957
transform 1 0 43424 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0947_
timestamp 1688980957
transform -1 0 43516 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1688980957
transform 1 0 44252 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0949_
timestamp 1688980957
transform 1 0 45264 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0950_
timestamp 1688980957
transform -1 0 44896 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1688980957
transform 1 0 46368 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _0952_
timestamp 1688980957
transform -1 0 47196 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _0953_
timestamp 1688980957
transform -1 0 45540 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  _0954_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44988 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _0955_
timestamp 1688980957
transform 1 0 43700 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _0956_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 43148 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _0957_
timestamp 1688980957
transform 1 0 43976 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0958_
timestamp 1688980957
transform -1 0 44528 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _0959_
timestamp 1688980957
transform -1 0 43976 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _0960_
timestamp 1688980957
transform 1 0 42504 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0961_
timestamp 1688980957
transform 1 0 42780 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _0962_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 43240 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _0963_
timestamp 1688980957
transform 1 0 44344 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _0964_
timestamp 1688980957
transform -1 0 46000 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _0965_
timestamp 1688980957
transform 1 0 44252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1688980957
transform 1 0 51888 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _0967_
timestamp 1688980957
transform -1 0 52256 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _0968_
timestamp 1688980957
transform -1 0 48116 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _0969_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 50140 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1688980957
transform 1 0 51704 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0971_
timestamp 1688980957
transform 1 0 49404 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _0972_
timestamp 1688980957
transform 1 0 48852 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _0973_
timestamp 1688980957
transform 1 0 9844 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0974_
timestamp 1688980957
transform -1 0 10856 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0975_
timestamp 1688980957
transform -1 0 4692 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0976_
timestamp 1688980957
transform -1 0 4324 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0977_
timestamp 1688980957
transform -1 0 6072 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0978_
timestamp 1688980957
transform -1 0 6808 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0979_
timestamp 1688980957
transform -1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0980_
timestamp 1688980957
transform 1 0 10488 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0981_
timestamp 1688980957
transform 1 0 5704 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0982_
timestamp 1688980957
transform 1 0 5336 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0983_
timestamp 1688980957
transform 1 0 6348 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0984_
timestamp 1688980957
transform -1 0 7268 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0985_
timestamp 1688980957
transform 1 0 8188 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0986_
timestamp 1688980957
transform -1 0 8832 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0987_
timestamp 1688980957
transform 1 0 4508 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0988_
timestamp 1688980957
transform -1 0 5060 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0989_
timestamp 1688980957
transform 1 0 8280 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0990_
timestamp 1688980957
transform 1 0 7912 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0991_
timestamp 1688980957
transform 1 0 3496 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0992_
timestamp 1688980957
transform -1 0 4784 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0993_
timestamp 1688980957
transform 1 0 6716 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0994_
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0995_
timestamp 1688980957
transform 1 0 4600 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0996_
timestamp 1688980957
transform -1 0 4968 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0997_
timestamp 1688980957
transform 1 0 9936 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _0998_
timestamp 1688980957
transform -1 0 10488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _0999_
timestamp 1688980957
transform 1 0 7360 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1000_
timestamp 1688980957
transform 1 0 7176 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1001_
timestamp 1688980957
transform 1 0 7176 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1002_
timestamp 1688980957
transform -1 0 7728 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1003_
timestamp 1688980957
transform 1 0 12696 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1004_
timestamp 1688980957
transform -1 0 13892 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1005_
timestamp 1688980957
transform 1 0 12880 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1688980957
transform 1 0 13340 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1007_
timestamp 1688980957
transform 1 0 10304 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1688980957
transform -1 0 11960 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12144 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1010_
timestamp 1688980957
transform -1 0 11408 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1011_
timestamp 1688980957
transform 1 0 12144 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1012_
timestamp 1688980957
transform -1 0 12420 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1013_
timestamp 1688980957
transform -1 0 13248 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014__1
timestamp 1688980957
transform 1 0 39468 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1688980957
transform 1 0 3864 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1688980957
transform 1 0 6072 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1688980957
transform 1 0 10212 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1688980957
transform 1 0 5336 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1688980957
transform 1 0 6716 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1688980957
transform -1 0 9752 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1688980957
transform 1 0 3312 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1688980957
transform 1 0 8188 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1688980957
transform 1 0 3864 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1688980957
transform 1 0 5888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1688980957
transform 1 0 10396 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1688980957
transform 1 0 7268 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1688980957
transform -1 0 8372 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1030_
timestamp 1688980957
transform 1 0 9108 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1031_
timestamp 1688980957
transform -1 0 9936 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _1032_
timestamp 1688980957
transform 1 0 41676 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_6  _1033_
timestamp 1688980957
transform -1 0 10212 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _1034_
timestamp 1688980957
transform -1 0 10764 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1035_
timestamp 1688980957
transform 1 0 9752 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1036_
timestamp 1688980957
transform 1 0 8372 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1037_
timestamp 1688980957
transform -1 0 6256 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1038_
timestamp 1688980957
transform -1 0 5888 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1039_
timestamp 1688980957
transform -1 0 6440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1040_
timestamp 1688980957
transform 1 0 4416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1041_
timestamp 1688980957
transform 1 0 6808 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1042_
timestamp 1688980957
transform -1 0 7084 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1043_
timestamp 1688980957
transform -1 0 7176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1044_
timestamp 1688980957
transform 1 0 6532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1045_
timestamp 1688980957
transform -1 0 12880 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1046_
timestamp 1688980957
transform -1 0 12328 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1047_
timestamp 1688980957
transform 1 0 10948 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1048_
timestamp 1688980957
transform 1 0 9568 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1049_
timestamp 1688980957
transform -1 0 10396 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1050_
timestamp 1688980957
transform -1 0 10120 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1051_
timestamp 1688980957
transform 1 0 10948 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1052_
timestamp 1688980957
transform 1 0 9568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1053_
timestamp 1688980957
transform -1 0 6716 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1054_
timestamp 1688980957
transform -1 0 6716 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1055_
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1056_
timestamp 1688980957
transform 1 0 2392 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1057_
timestamp 1688980957
transform -1 0 7728 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1058_
timestamp 1688980957
transform -1 0 6992 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1059_
timestamp 1688980957
transform -1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1060_
timestamp 1688980957
transform 1 0 6440 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1061_
timestamp 1688980957
transform -1 0 12144 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1062_
timestamp 1688980957
transform -1 0 11868 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1063_
timestamp 1688980957
transform 1 0 10856 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1064_
timestamp 1688980957
transform 1 0 9568 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1065_
timestamp 1688980957
transform 1 0 4508 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1066_
timestamp 1688980957
transform -1 0 5060 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1067_
timestamp 1688980957
transform -1 0 4784 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1068_
timestamp 1688980957
transform 1 0 4508 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1069_
timestamp 1688980957
transform -1 0 4324 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1070_
timestamp 1688980957
transform -1 0 3680 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1071_
timestamp 1688980957
transform -1 0 3588 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1072_
timestamp 1688980957
transform -1 0 4048 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1073_
timestamp 1688980957
transform 1 0 3956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1074_
timestamp 1688980957
transform 1 0 2116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1075_
timestamp 1688980957
transform -1 0 4048 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1076_
timestamp 1688980957
transform 1 0 3772 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1077_
timestamp 1688980957
transform -1 0 3588 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1078_
timestamp 1688980957
transform -1 0 3680 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1079_
timestamp 1688980957
transform 1 0 3956 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1080_
timestamp 1688980957
transform 1 0 2208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1081_
timestamp 1688980957
transform -1 0 4324 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1082_
timestamp 1688980957
transform 1 0 3772 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1083_
timestamp 1688980957
transform 1 0 3220 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1084_
timestamp 1688980957
transform -1 0 4324 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1085_
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1086_
timestamp 1688980957
transform 1 0 2300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1087_
timestamp 1688980957
transform -1 0 4232 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1088_
timestamp 1688980957
transform -1 0 3496 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1089_
timestamp 1688980957
transform -1 0 3128 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1090_
timestamp 1688980957
transform -1 0 4784 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1091_
timestamp 1688980957
transform -1 0 8832 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  _1092_
timestamp 1688980957
transform -1 0 9476 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1093_
timestamp 1688980957
transform -1 0 3496 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1094_
timestamp 1688980957
transform 1 0 3404 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1095_
timestamp 1688980957
transform -1 0 4140 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1096_
timestamp 1688980957
transform 1 0 4140 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1097_
timestamp 1688980957
transform 1 0 3220 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1098_
timestamp 1688980957
transform -1 0 4508 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1099_
timestamp 1688980957
transform 1 0 3404 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1100_
timestamp 1688980957
transform 1 0 2116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1101_
timestamp 1688980957
transform -1 0 4232 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1102_
timestamp 1688980957
transform 1 0 3220 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1103_
timestamp 1688980957
transform 1 0 2852 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1104_
timestamp 1688980957
transform -1 0 4784 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1105_
timestamp 1688980957
transform -1 0 5704 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1106_
timestamp 1688980957
transform 1 0 4048 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1107_
timestamp 1688980957
transform -1 0 3588 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1108_
timestamp 1688980957
transform -1 0 3496 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1109_
timestamp 1688980957
transform 1 0 1932 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1110_
timestamp 1688980957
transform -1 0 4324 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1111_
timestamp 1688980957
transform -1 0 3680 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1112_
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1113_
timestamp 1688980957
transform -1 0 4048 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1114_
timestamp 1688980957
transform 1 0 3220 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1115_
timestamp 1688980957
transform 1 0 1840 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1116_
timestamp 1688980957
transform -1 0 9476 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1117_
timestamp 1688980957
transform 1 0 8280 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1118_
timestamp 1688980957
transform 1 0 7636 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1119_
timestamp 1688980957
transform -1 0 4140 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1120_
timestamp 1688980957
transform -1 0 4508 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1121_
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1122_
timestamp 1688980957
transform -1 0 6256 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1123_
timestamp 1688980957
transform 1 0 7360 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1124_
timestamp 1688980957
transform 1 0 5612 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1125_
timestamp 1688980957
transform -1 0 9016 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1126_
timestamp 1688980957
transform -1 0 8648 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1127_
timestamp 1688980957
transform 1 0 7728 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1128_
timestamp 1688980957
transform -1 0 9200 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1129_
timestamp 1688980957
transform 1 0 8464 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1130_
timestamp 1688980957
transform 1 0 7176 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1131_
timestamp 1688980957
transform -1 0 4416 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1132_
timestamp 1688980957
transform -1 0 3588 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1133_
timestamp 1688980957
transform 1 0 1840 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1134_
timestamp 1688980957
transform -1 0 7268 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1135_
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1136_
timestamp 1688980957
transform 1 0 6624 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1137_
timestamp 1688980957
transform -1 0 8740 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1138_
timestamp 1688980957
transform -1 0 8740 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1139_
timestamp 1688980957
transform 1 0 8004 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1140_
timestamp 1688980957
transform 1 0 49588 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1141_
timestamp 1688980957
transform 1 0 50876 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1142_
timestamp 1688980957
transform -1 0 47196 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1143_
timestamp 1688980957
transform -1 0 43056 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1144_
timestamp 1688980957
transform 1 0 43056 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1145_
timestamp 1688980957
transform -1 0 44160 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1146_
timestamp 1688980957
transform -1 0 45264 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1147_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42964 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1148_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 41768 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1149_
timestamp 1688980957
transform 1 0 40756 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1150_
timestamp 1688980957
transform 1 0 57776 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1151_
timestamp 1688980957
transform 1 0 58144 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1152_
timestamp 1688980957
transform -1 0 56580 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1153_
timestamp 1688980957
transform -1 0 55200 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1154_
timestamp 1688980957
transform 1 0 48300 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1155_
timestamp 1688980957
transform 1 0 53544 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1156_
timestamp 1688980957
transform 1 0 58144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1157_
timestamp 1688980957
transform 1 0 55292 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1158_
timestamp 1688980957
transform -1 0 56028 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1159_
timestamp 1688980957
transform 1 0 53084 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1160_
timestamp 1688980957
transform 1 0 53176 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1161_
timestamp 1688980957
transform 1 0 52808 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1162_
timestamp 1688980957
transform 1 0 58236 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1163_
timestamp 1688980957
transform -1 0 58236 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1164_
timestamp 1688980957
transform 1 0 57500 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1165_
timestamp 1688980957
transform 1 0 55568 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1166_
timestamp 1688980957
transform -1 0 57500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1167_
timestamp 1688980957
transform -1 0 57224 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1168_
timestamp 1688980957
transform -1 0 55660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1169_
timestamp 1688980957
transform 1 0 55108 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1170_
timestamp 1688980957
transform 1 0 55292 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1171_
timestamp 1688980957
transform 1 0 52716 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1172_
timestamp 1688980957
transform 1 0 52716 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1173_
timestamp 1688980957
transform 1 0 50508 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1174_
timestamp 1688980957
transform -1 0 58144 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1175_
timestamp 1688980957
transform -1 0 58420 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1176_
timestamp 1688980957
transform 1 0 57316 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1177_
timestamp 1688980957
transform 1 0 57868 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1178_
timestamp 1688980957
transform 1 0 57040 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1179_
timestamp 1688980957
transform 1 0 57500 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1180_
timestamp 1688980957
transform -1 0 58420 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1181_
timestamp 1688980957
transform 1 0 50416 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1182_
timestamp 1688980957
transform 1 0 49128 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1183_
timestamp 1688980957
transform 1 0 47104 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1184_
timestamp 1688980957
transform -1 0 49404 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1185_
timestamp 1688980957
transform -1 0 48392 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1186_
timestamp 1688980957
transform 1 0 47564 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1187_
timestamp 1688980957
transform -1 0 48668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1188_
timestamp 1688980957
transform -1 0 48484 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1189_
timestamp 1688980957
transform -1 0 48208 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1190_
timestamp 1688980957
transform 1 0 47564 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1191_
timestamp 1688980957
transform -1 0 49404 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1192_
timestamp 1688980957
transform 1 0 50232 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1193_
timestamp 1688980957
transform -1 0 49404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1194_
timestamp 1688980957
transform -1 0 49128 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1195_
timestamp 1688980957
transform 1 0 50140 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1196_
timestamp 1688980957
transform -1 0 49956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1197_
timestamp 1688980957
transform 1 0 49128 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1198_
timestamp 1688980957
transform 1 0 48484 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1199_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 49220 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1200_
timestamp 1688980957
transform 1 0 49404 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1201_
timestamp 1688980957
transform -1 0 49864 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1202_
timestamp 1688980957
transform -1 0 55936 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1203_
timestamp 1688980957
transform 1 0 56764 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1204_
timestamp 1688980957
transform -1 0 58420 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1205_
timestamp 1688980957
transform -1 0 58144 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1206_
timestamp 1688980957
transform -1 0 58604 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1207_
timestamp 1688980957
transform 1 0 57500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1208_
timestamp 1688980957
transform 1 0 57224 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1209_
timestamp 1688980957
transform 1 0 56304 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1210_
timestamp 1688980957
transform 1 0 42412 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1211_
timestamp 1688980957
transform -1 0 47472 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_4  _1212_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 49128 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1213_
timestamp 1688980957
transform 1 0 47932 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1214_
timestamp 1688980957
transform -1 0 48760 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1215_
timestamp 1688980957
transform -1 0 47472 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1216_
timestamp 1688980957
transform 1 0 48300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1217_
timestamp 1688980957
transform 1 0 50876 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _1218_
timestamp 1688980957
transform -1 0 53268 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1219_
timestamp 1688980957
transform 1 0 58144 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1220_
timestamp 1688980957
transform 1 0 52256 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1221_
timestamp 1688980957
transform 1 0 52716 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1222_
timestamp 1688980957
transform 1 0 52072 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1223_
timestamp 1688980957
transform -1 0 52164 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1224_
timestamp 1688980957
transform -1 0 51888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1225_
timestamp 1688980957
transform -1 0 51888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1226_
timestamp 1688980957
transform 1 0 50968 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1227_
timestamp 1688980957
transform 1 0 51336 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1228_
timestamp 1688980957
transform -1 0 51704 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1229_
timestamp 1688980957
transform -1 0 51980 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1230_
timestamp 1688980957
transform -1 0 53820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1231_
timestamp 1688980957
transform -1 0 54372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1232_
timestamp 1688980957
transform -1 0 53912 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1233_
timestamp 1688980957
transform 1 0 53268 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1234_
timestamp 1688980957
transform -1 0 54004 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1235_
timestamp 1688980957
transform -1 0 53912 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1236_
timestamp 1688980957
transform -1 0 54188 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1237_
timestamp 1688980957
transform 1 0 52072 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1238_
timestamp 1688980957
transform 1 0 51796 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1239_
timestamp 1688980957
transform -1 0 51796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1240_
timestamp 1688980957
transform 1 0 51336 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1241_
timestamp 1688980957
transform 1 0 58144 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1242_
timestamp 1688980957
transform -1 0 52164 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1243_
timestamp 1688980957
transform -1 0 52440 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1244_
timestamp 1688980957
transform 1 0 51980 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1245_
timestamp 1688980957
transform 1 0 58052 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1246_
timestamp 1688980957
transform -1 0 52164 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1247_
timestamp 1688980957
transform -1 0 52440 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1248_
timestamp 1688980957
transform -1 0 51888 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1249_
timestamp 1688980957
transform 1 0 51612 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1250_
timestamp 1688980957
transform 1 0 51244 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1251_
timestamp 1688980957
transform -1 0 52532 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1252_
timestamp 1688980957
transform 1 0 51520 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1253_
timestamp 1688980957
transform 1 0 57868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1254_
timestamp 1688980957
transform -1 0 55200 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1255_
timestamp 1688980957
transform -1 0 54924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1256_
timestamp 1688980957
transform 1 0 54004 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1257_
timestamp 1688980957
transform 1 0 54648 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1258_
timestamp 1688980957
transform 1 0 54372 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1259_
timestamp 1688980957
transform 1 0 58236 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1260_
timestamp 1688980957
transform -1 0 55200 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1261_
timestamp 1688980957
transform 1 0 54188 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1262_
timestamp 1688980957
transform 1 0 54280 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1263_
timestamp 1688980957
transform 1 0 54648 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1264_
timestamp 1688980957
transform 1 0 53452 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1265_
timestamp 1688980957
transform 1 0 53452 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1266_
timestamp 1688980957
transform 1 0 52440 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1267_
timestamp 1688980957
transform -1 0 52164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1268_
timestamp 1688980957
transform 1 0 51612 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1269_
timestamp 1688980957
transform -1 0 51980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1270_
timestamp 1688980957
transform 1 0 50692 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1271_
timestamp 1688980957
transform -1 0 50692 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1272_
timestamp 1688980957
transform 1 0 50324 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1273_
timestamp 1688980957
transform 1 0 50324 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1274_
timestamp 1688980957
transform 1 0 50416 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1275_
timestamp 1688980957
transform 1 0 57592 0 1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1276_
timestamp 1688980957
transform 1 0 57040 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _1277_
timestamp 1688980957
transform 1 0 57316 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1278_
timestamp 1688980957
transform -1 0 58236 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1279_
timestamp 1688980957
transform 1 0 55844 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1280_
timestamp 1688980957
transform 1 0 56948 0 -1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1281_
timestamp 1688980957
transform 1 0 56120 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1282_
timestamp 1688980957
transform -1 0 55844 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1283_
timestamp 1688980957
transform 1 0 49128 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_1  _1284_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 50140 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1285_
timestamp 1688980957
transform -1 0 50416 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1286_
timestamp 1688980957
transform 1 0 49312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1287_
timestamp 1688980957
transform 1 0 47012 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1288_
timestamp 1688980957
transform 1 0 47104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1289_
timestamp 1688980957
transform -1 0 58420 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1290_
timestamp 1688980957
transform -1 0 57592 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1291_
timestamp 1688980957
transform 1 0 56948 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1292_
timestamp 1688980957
transform 1 0 56948 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1293_
timestamp 1688980957
transform -1 0 58420 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1294_
timestamp 1688980957
transform -1 0 58144 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1295_
timestamp 1688980957
transform -1 0 57776 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1296_
timestamp 1688980957
transform 1 0 57224 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1297_
timestamp 1688980957
transform -1 0 57224 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1298_
timestamp 1688980957
transform 1 0 51888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1299_
timestamp 1688980957
transform 1 0 58144 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1300_
timestamp 1688980957
transform -1 0 57868 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1301_
timestamp 1688980957
transform 1 0 57132 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1302_
timestamp 1688980957
transform 1 0 56948 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1303_
timestamp 1688980957
transform 1 0 58236 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1304_
timestamp 1688980957
transform -1 0 58236 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1305_
timestamp 1688980957
transform -1 0 57776 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1306_
timestamp 1688980957
transform 1 0 57224 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1307_
timestamp 1688980957
transform -1 0 57132 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1308_
timestamp 1688980957
transform 1 0 51612 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1309_
timestamp 1688980957
transform 1 0 51244 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1310_
timestamp 1688980957
transform -1 0 51612 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1311_
timestamp 1688980957
transform -1 0 58420 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1312_
timestamp 1688980957
transform -1 0 58144 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1313_
timestamp 1688980957
transform 1 0 57868 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1314_
timestamp 1688980957
transform 1 0 57868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1315_
timestamp 1688980957
transform -1 0 57500 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1316_
timestamp 1688980957
transform -1 0 58236 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1317_
timestamp 1688980957
transform -1 0 58236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1318_
timestamp 1688980957
transform 1 0 51520 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1319_
timestamp 1688980957
transform 1 0 51244 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1320_
timestamp 1688980957
transform 1 0 58144 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1321_
timestamp 1688980957
transform -1 0 49588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1322_
timestamp 1688980957
transform 1 0 48668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1323_
timestamp 1688980957
transform -1 0 49312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1324_
timestamp 1688980957
transform -1 0 50140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1325_
timestamp 1688980957
transform -1 0 49588 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1326_
timestamp 1688980957
transform 1 0 49036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1327_
timestamp 1688980957
transform 1 0 49128 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1328_
timestamp 1688980957
transform -1 0 49496 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1329_
timestamp 1688980957
transform 1 0 50140 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1330_
timestamp 1688980957
transform 1 0 50140 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1331_
timestamp 1688980957
transform 1 0 49588 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1332_
timestamp 1688980957
transform -1 0 49496 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1333_
timestamp 1688980957
transform -1 0 49772 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1334_
timestamp 1688980957
transform 1 0 50140 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1335_
timestamp 1688980957
transform -1 0 49864 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1336_
timestamp 1688980957
transform 1 0 56120 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1337_
timestamp 1688980957
transform 1 0 55476 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1338_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 58512 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1339_
timestamp 1688980957
transform 1 0 50876 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1340_
timestamp 1688980957
transform 1 0 49772 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1341_
timestamp 1688980957
transform -1 0 49588 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1342_
timestamp 1688980957
transform -1 0 49220 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1343_
timestamp 1688980957
transform -1 0 48944 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1344_
timestamp 1688980957
transform 1 0 49220 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1345_
timestamp 1688980957
transform 1 0 52348 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1346_
timestamp 1688980957
transform -1 0 57868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1347_
timestamp 1688980957
transform 1 0 52072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1348_
timestamp 1688980957
transform 1 0 52808 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1349_
timestamp 1688980957
transform -1 0 53544 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1350_
timestamp 1688980957
transform -1 0 54832 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1351_
timestamp 1688980957
transform -1 0 54004 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1352_
timestamp 1688980957
transform -1 0 54740 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1353_
timestamp 1688980957
transform 1 0 53820 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1354_
timestamp 1688980957
transform -1 0 54464 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1355_
timestamp 1688980957
transform 1 0 52992 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1356_
timestamp 1688980957
transform 1 0 52900 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1357_
timestamp 1688980957
transform -1 0 53820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1358_
timestamp 1688980957
transform -1 0 54464 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1359_
timestamp 1688980957
transform -1 0 54004 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1360_
timestamp 1688980957
transform -1 0 55200 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1361_
timestamp 1688980957
transform -1 0 54372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _1362_
timestamp 1688980957
transform -1 0 53912 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1363_
timestamp 1688980957
transform -1 0 53544 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1364_
timestamp 1688980957
transform 1 0 51980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1365_
timestamp 1688980957
transform 1 0 51704 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1366_
timestamp 1688980957
transform 1 0 51796 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _1367_
timestamp 1688980957
transform 1 0 52992 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1368_
timestamp 1688980957
transform -1 0 58420 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1369_
timestamp 1688980957
transform 1 0 52900 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1370_
timestamp 1688980957
transform 1 0 53268 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1371_
timestamp 1688980957
transform 1 0 52992 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1372_
timestamp 1688980957
transform 1 0 57500 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1373_
timestamp 1688980957
transform -1 0 55016 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1374_
timestamp 1688980957
transform -1 0 54648 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1375_
timestamp 1688980957
transform 1 0 54096 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1376_
timestamp 1688980957
transform 1 0 54280 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1377_
timestamp 1688980957
transform 1 0 53544 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1378_
timestamp 1688980957
transform -1 0 53544 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1379_
timestamp 1688980957
transform 1 0 53268 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1380_
timestamp 1688980957
transform 1 0 58144 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1381_
timestamp 1688980957
transform -1 0 54740 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1382_
timestamp 1688980957
transform 1 0 53820 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1383_
timestamp 1688980957
transform 1 0 53452 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1384_
timestamp 1688980957
transform -1 0 53728 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1385_
timestamp 1688980957
transform 1 0 53176 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1386_
timestamp 1688980957
transform 1 0 58144 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1387_
timestamp 1688980957
transform -1 0 54832 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1388_
timestamp 1688980957
transform -1 0 54832 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1389_
timestamp 1688980957
transform -1 0 54464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1390_
timestamp 1688980957
transform 1 0 54188 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1391_
timestamp 1688980957
transform 1 0 53728 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1392_
timestamp 1688980957
transform -1 0 53728 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1393_
timestamp 1688980957
transform 1 0 52716 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1394_
timestamp 1688980957
transform 1 0 52992 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1395_
timestamp 1688980957
transform 1 0 52164 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1396_
timestamp 1688980957
transform -1 0 51704 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1397_
timestamp 1688980957
transform 1 0 50784 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1398_
timestamp 1688980957
transform -1 0 51336 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1399_
timestamp 1688980957
transform 1 0 50232 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1400_
timestamp 1688980957
transform 1 0 50416 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1401_
timestamp 1688980957
transform 1 0 50508 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1402_
timestamp 1688980957
transform 1 0 57500 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1403_
timestamp 1688980957
transform 1 0 57224 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1404_
timestamp 1688980957
transform 1 0 56948 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1405_
timestamp 1688980957
transform -1 0 57500 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1406_
timestamp 1688980957
transform -1 0 58144 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1407_
timestamp 1688980957
transform 1 0 56580 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1408_
timestamp 1688980957
transform 1 0 57132 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1409_
timestamp 1688980957
transform 1 0 56672 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1410_
timestamp 1688980957
transform -1 0 56580 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1411_
timestamp 1688980957
transform 1 0 49588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1412_
timestamp 1688980957
transform 1 0 49680 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1413_
timestamp 1688980957
transform 1 0 49864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1414_
timestamp 1688980957
transform 1 0 49312 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1415_
timestamp 1688980957
transform -1 0 48576 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1416_
timestamp 1688980957
transform 1 0 47196 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _1417_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 41768 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1418_
timestamp 1688980957
transform 1 0 41492 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_2  _1419_
timestamp 1688980957
transform 1 0 41676 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  _1420_
timestamp 1688980957
transform -1 0 49312 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1421_
timestamp 1688980957
transform -1 0 51704 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1422_
timestamp 1688980957
transform -1 0 48024 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1423_
timestamp 1688980957
transform -1 0 47196 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1424_
timestamp 1688980957
transform -1 0 51336 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1425_
timestamp 1688980957
transform 1 0 50324 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1426_
timestamp 1688980957
transform -1 0 49956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1427_
timestamp 1688980957
transform -1 0 48760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1428_
timestamp 1688980957
transform 1 0 56028 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1429_
timestamp 1688980957
transform 1 0 54188 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1430_
timestamp 1688980957
transform -1 0 48116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1431_
timestamp 1688980957
transform -1 0 46920 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1432_
timestamp 1688980957
transform -1 0 52256 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1433_
timestamp 1688980957
transform 1 0 52256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1434_
timestamp 1688980957
transform -1 0 47840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1435_
timestamp 1688980957
transform -1 0 47288 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1436_
timestamp 1688980957
transform -1 0 51336 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1437_
timestamp 1688980957
transform 1 0 49680 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1438_
timestamp 1688980957
transform -1 0 57040 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1439_
timestamp 1688980957
transform -1 0 57776 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1440_
timestamp 1688980957
transform 1 0 56304 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1441_
timestamp 1688980957
transform -1 0 55200 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1442_
timestamp 1688980957
transform 1 0 56212 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1443_
timestamp 1688980957
transform 1 0 54832 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1444_
timestamp 1688980957
transform -1 0 58328 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1445_
timestamp 1688980957
transform -1 0 57776 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1446_
timestamp 1688980957
transform 1 0 56488 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1447_
timestamp 1688980957
transform -1 0 55660 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1448_
timestamp 1688980957
transform -1 0 56856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1449_
timestamp 1688980957
transform 1 0 55292 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1450_
timestamp 1688980957
transform -1 0 56028 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1451_
timestamp 1688980957
transform -1 0 56580 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1452_
timestamp 1688980957
transform 1 0 54832 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1453_
timestamp 1688980957
transform -1 0 53176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1454_
timestamp 1688980957
transform 1 0 54740 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1455_
timestamp 1688980957
transform 1 0 52164 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1456_
timestamp 1688980957
transform -1 0 57776 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1457_
timestamp 1688980957
transform -1 0 57592 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1458_
timestamp 1688980957
transform -1 0 57316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1459_
timestamp 1688980957
transform -1 0 55568 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1460_
timestamp 1688980957
transform 1 0 56212 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1461_
timestamp 1688980957
transform 1 0 54740 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _1462_
timestamp 1688980957
transform 1 0 51152 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  _1463_
timestamp 1688980957
transform 1 0 51704 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1464_
timestamp 1688980957
transform 1 0 56672 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1465_
timestamp 1688980957
transform -1 0 55108 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1466_
timestamp 1688980957
transform -1 0 52716 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1467_
timestamp 1688980957
transform 1 0 52164 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1468_
timestamp 1688980957
transform -1 0 58052 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1469_
timestamp 1688980957
transform 1 0 56028 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1470_
timestamp 1688980957
transform 1 0 56028 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1471_
timestamp 1688980957
transform 1 0 54832 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1472_
timestamp 1688980957
transform -1 0 57224 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1473_
timestamp 1688980957
transform -1 0 56764 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1474_
timestamp 1688980957
transform 1 0 56028 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1475_
timestamp 1688980957
transform 1 0 54648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1476_
timestamp 1688980957
transform -1 0 56948 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1477_
timestamp 1688980957
transform -1 0 57316 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1478_
timestamp 1688980957
transform -1 0 53728 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1479_
timestamp 1688980957
transform -1 0 51612 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1480_
timestamp 1688980957
transform -1 0 55108 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1481_
timestamp 1688980957
transform -1 0 54096 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1482_
timestamp 1688980957
transform -1 0 52624 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1483_
timestamp 1688980957
transform -1 0 51796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1484_
timestamp 1688980957
transform -1 0 57684 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1485_
timestamp 1688980957
transform -1 0 56672 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1486_
timestamp 1688980957
transform 1 0 54924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1487_
timestamp 1688980957
transform 1 0 54648 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1488_
timestamp 1688980957
transform -1 0 55200 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1489_
timestamp 1688980957
transform -1 0 56304 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1490_
timestamp 1688980957
transform 1 0 51336 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1491_
timestamp 1688980957
transform 1 0 52072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1492_
timestamp 1688980957
transform -1 0 56488 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1493_
timestamp 1688980957
transform 1 0 56488 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1494_
timestamp 1688980957
transform -1 0 53084 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1495_
timestamp 1688980957
transform 1 0 52808 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1496_
timestamp 1688980957
transform 1 0 46828 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1497_
timestamp 1688980957
transform -1 0 45632 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1498_
timestamp 1688980957
transform -1 0 49128 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1499_
timestamp 1688980957
transform -1 0 47748 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1500_
timestamp 1688980957
transform 1 0 45264 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1501_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 47748 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1502_
timestamp 1688980957
transform -1 0 48484 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1503_
timestamp 1688980957
transform -1 0 39744 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1504_
timestamp 1688980957
transform -1 0 40204 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1505_
timestamp 1688980957
transform -1 0 38548 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1506_
timestamp 1688980957
transform 1 0 38180 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1507_
timestamp 1688980957
transform 1 0 38272 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1508_
timestamp 1688980957
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1509_
timestamp 1688980957
transform 1 0 39192 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1510_
timestamp 1688980957
transform 1 0 39284 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1511_
timestamp 1688980957
transform 1 0 39100 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1512_
timestamp 1688980957
transform -1 0 40020 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_1  _1513_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39836 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1514_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 38548 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o22a_1  _1515_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39836 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1516_
timestamp 1688980957
transform -1 0 38364 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1517_
timestamp 1688980957
transform 1 0 38456 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1518_
timestamp 1688980957
transform 1 0 37904 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1519_
timestamp 1688980957
transform 1 0 38548 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1520_
timestamp 1688980957
transform -1 0 40940 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1521_
timestamp 1688980957
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1522_
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1523_
timestamp 1688980957
transform 1 0 40572 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_2  _1524_
timestamp 1688980957
transform -1 0 38824 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1525_
timestamp 1688980957
transform 1 0 36800 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1526_
timestamp 1688980957
transform -1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1527_
timestamp 1688980957
transform -1 0 37904 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1528_
timestamp 1688980957
transform 1 0 37076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1529_
timestamp 1688980957
transform 1 0 36432 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1530_
timestamp 1688980957
transform -1 0 37536 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1531_
timestamp 1688980957
transform 1 0 35420 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1532_
timestamp 1688980957
transform -1 0 38732 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1533_
timestamp 1688980957
transform 1 0 37996 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1534_
timestamp 1688980957
transform -1 0 39836 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1535_
timestamp 1688980957
transform 1 0 37352 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1536_
timestamp 1688980957
transform -1 0 43148 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1537_
timestamp 1688980957
transform -1 0 43148 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1538_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 42596 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1539_
timestamp 1688980957
transform -1 0 42872 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1540_
timestamp 1688980957
transform 1 0 41308 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1541_
timestamp 1688980957
transform -1 0 43424 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1542_
timestamp 1688980957
transform 1 0 44988 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1543_
timestamp 1688980957
transform -1 0 44712 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _1544_
timestamp 1688980957
transform 1 0 41768 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1545_
timestamp 1688980957
transform 1 0 45080 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1546_
timestamp 1688980957
transform 1 0 43884 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1547_
timestamp 1688980957
transform 1 0 48024 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1548_
timestamp 1688980957
transform -1 0 46460 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1549_
timestamp 1688980957
transform 1 0 46276 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1550_
timestamp 1688980957
transform 1 0 48484 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1551_
timestamp 1688980957
transform 1 0 48300 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_1  _1552_
timestamp 1688980957
transform 1 0 48208 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1553_
timestamp 1688980957
transform -1 0 50232 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1554_
timestamp 1688980957
transform 1 0 48852 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1555_
timestamp 1688980957
transform -1 0 48116 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1556_
timestamp 1688980957
transform 1 0 47196 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1557_
timestamp 1688980957
transform 1 0 47564 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1558_
timestamp 1688980957
transform -1 0 46920 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1559_
timestamp 1688980957
transform -1 0 46644 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dfstp_1  _1560_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 47472 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1561_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42964 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1562_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 50784 0 -1 30464
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1563_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 44988 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1564_
timestamp 1688980957
transform 1 0 47472 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1565_
timestamp 1688980957
transform 1 0 42504 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1566_
timestamp 1688980957
transform 1 0 37352 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1567_
timestamp 1688980957
transform 1 0 46644 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1568_
timestamp 1688980957
transform 1 0 40204 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1569_
timestamp 1688980957
transform 1 0 43792 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _1570_
timestamp 1688980957
transform 1 0 45632 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1571_
timestamp 1688980957
transform -1 0 42320 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1572_
timestamp 1688980957
transform 1 0 41308 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1573_
timestamp 1688980957
transform 1 0 40940 0 1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1574_
timestamp 1688980957
transform -1 0 46460 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1575_
timestamp 1688980957
transform -1 0 51152 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1576_
timestamp 1688980957
transform 1 0 47564 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  _1577_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 10488 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1578_
timestamp 1688980957
transform -1 0 5796 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1579_
timestamp 1688980957
transform -1 0 8004 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1580_
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1581_
timestamp 1688980957
transform -1 0 5336 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1582_
timestamp 1688980957
transform -1 0 8096 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1583_
timestamp 1688980957
transform -1 0 10304 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1584_
timestamp 1688980957
transform -1 0 6256 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1585_
timestamp 1688980957
transform -1 0 8832 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1586_
timestamp 1688980957
transform -1 0 5704 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1587_
timestamp 1688980957
transform -1 0 7360 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1588_
timestamp 1688980957
transform -1 0 5796 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1589_
timestamp 1688980957
transform -1 0 11408 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1590_
timestamp 1688980957
transform -1 0 7360 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1591_
timestamp 1688980957
transform -1 0 7820 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1592_
timestamp 1688980957
transform -1 0 14444 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1593_
timestamp 1688980957
transform 1 0 13156 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1594_
timestamp 1688980957
transform -1 0 12420 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1595_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13984 0 1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1596_
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _1597_
timestamp 1688980957
transform 1 0 39836 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_1  _1598_
timestamp 1688980957
transform -1 0 13064 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1599_
timestamp 1688980957
transform 1 0 4416 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1600_
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1601_
timestamp 1688980957
transform 1 0 10488 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1688980957
transform 1 0 5612 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1603_
timestamp 1688980957
transform 1 0 7268 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1604_
timestamp 1688980957
transform 1 0 9292 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1605_
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1606_
timestamp 1688980957
transform -1 0 8832 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1607_
timestamp 1688980957
transform 1 0 4140 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1608_
timestamp 1688980957
transform -1 0 7360 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1609_
timestamp 1688980957
transform 1 0 4048 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1610_
timestamp 1688980957
transform 1 0 10488 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1688980957
transform 1 0 7544 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 1688980957
transform 1 0 8096 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1688980957
transform 1 0 12512 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_2  _1614_
timestamp 1688980957
transform -1 0 10856 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1615_
timestamp 1688980957
transform -1 0 6164 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1616_
timestamp 1688980957
transform -1 0 8832 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1617_
timestamp 1688980957
transform -1 0 10948 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1618_
timestamp 1688980957
transform -1 0 12052 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1619_
timestamp 1688980957
transform -1 0 3496 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1620_
timestamp 1688980957
transform -1 0 8556 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1621_
timestamp 1688980957
transform -1 0 11960 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1622_
timestamp 1688980957
transform -1 0 6256 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1623_
timestamp 1688980957
transform -1 0 3220 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1624_
timestamp 1688980957
transform -1 0 3220 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1625_
timestamp 1688980957
transform -1 0 3220 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1626_
timestamp 1688980957
transform -1 0 3220 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1627_
timestamp 1688980957
transform -1 0 3220 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1628_
timestamp 1688980957
transform -1 0 3220 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1629_
timestamp 1688980957
transform -1 0 3220 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1630_
timestamp 1688980957
transform -1 0 3220 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1631_
timestamp 1688980957
transform -1 0 3220 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1632_
timestamp 1688980957
transform -1 0 3220 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1633_
timestamp 1688980957
transform -1 0 3220 0 -1 34816
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1634_
timestamp 1688980957
transform 1 0 4416 0 -1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1635_
timestamp 1688980957
transform -1 0 3220 0 1 35904
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1636_
timestamp 1688980957
transform -1 0 5796 0 -1 36992
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1637_
timestamp 1688980957
transform -1 0 3220 0 1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1638_
timestamp 1688980957
transform -1 0 10212 0 -1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _1639_
timestamp 1688980957
transform -1 0 5612 0 -1 39168
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _1640_
timestamp 1688980957
transform -1 0 8280 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1641_
timestamp 1688980957
transform -1 0 10856 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1642_
timestamp 1688980957
transform -1 0 8280 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1643_
timestamp 1688980957
transform -1 0 3312 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _1644_
timestamp 1688980957
transform -1 0 7452 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _1645_
timestamp 1688980957
transform -1 0 10580 0 -1 36992
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _1646_
timestamp 1688980957
transform 1 0 40204 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfxtp_2  _1647_
timestamp 1688980957
transform -1 0 47104 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1688980957
transform -1 0 47104 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1688980957
transform 1 0 46184 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1688980957
transform 1 0 47564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1688980957
transform 1 0 46276 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1688980957
transform 1 0 50232 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1688980957
transform 1 0 48208 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1654_
timestamp 1688980957
transform 1 0 53728 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1655_
timestamp 1688980957
transform 1 0 46000 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1656_
timestamp 1688980957
transform 1 0 52716 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1657_
timestamp 1688980957
transform 1 0 46644 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1658_
timestamp 1688980957
transform 1 0 50140 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1659_
timestamp 1688980957
transform 1 0 56212 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1660_
timestamp 1688980957
transform 1 0 55292 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1661_
timestamp 1688980957
transform 1 0 56856 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1662_
timestamp 1688980957
transform 1 0 55108 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1663_
timestamp 1688980957
transform 1 0 55292 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1664_
timestamp 1688980957
transform 1 0 52532 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1665_
timestamp 1688980957
transform 1 0 56764 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1666_
timestamp 1688980957
transform 1 0 55292 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1667_
timestamp 1688980957
transform 1 0 54464 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1668_
timestamp 1688980957
transform 1 0 52716 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1669_
timestamp 1688980957
transform 1 0 56396 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1670_
timestamp 1688980957
transform 1 0 55292 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1671_
timestamp 1688980957
transform 1 0 56212 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1672_
timestamp 1688980957
transform 1 0 55016 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1673_
timestamp 1688980957
transform 1 0 56764 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1674_
timestamp 1688980957
transform 1 0 51060 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1675_
timestamp 1688980957
transform 1 0 53452 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1676_
timestamp 1688980957
transform 1 0 51152 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1677_
timestamp 1688980957
transform 1 0 56120 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1678_
timestamp 1688980957
transform 1 0 55292 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1679_
timestamp 1688980957
transform -1 0 56764 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1680_
timestamp 1688980957
transform -1 0 52072 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1681_
timestamp 1688980957
transform 1 0 56764 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1682_
timestamp 1688980957
transform 1 0 52532 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_1  _1683_
timestamp 1688980957
transform -1 0 47196 0 -1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1684_
timestamp 1688980957
transform 1 0 48208 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1685_
timestamp 1688980957
transform 1 0 36432 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1686_
timestamp 1688980957
transform -1 0 41676 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1687_
timestamp 1688980957
transform 1 0 36708 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1688_
timestamp 1688980957
transform 1 0 35144 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1689_
timestamp 1688980957
transform 1 0 35420 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1690_
timestamp 1688980957
transform 1 0 37444 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1691_
timestamp 1688980957
transform 1 0 40296 0 1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1692_
timestamp 1688980957
transform 1 0 41584 0 1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1693_
timestamp 1688980957
transform -1 0 46368 0 -1 33728
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1694_
timestamp 1688980957
transform 1 0 48668 0 -1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1695_
timestamp 1688980957
transform -1 0 50876 0 -1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _1696_
timestamp 1688980957
transform 1 0 44988 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12512 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A
timestamp 1688980957
transform 1 0 13340 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A
timestamp 1688980957
transform -1 0 8740 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A
timestamp 1688980957
transform -1 0 9384 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A
timestamp 1688980957
transform -1 0 12236 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A
timestamp 1688980957
transform 1 0 12972 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B
timestamp 1688980957
transform 1 0 5520 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A
timestamp 1688980957
transform 1 0 5704 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A
timestamp 1688980957
transform 1 0 10212 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A
timestamp 1688980957
transform 1 0 7268 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A
timestamp 1688980957
transform 1 0 6624 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A
timestamp 1688980957
transform 1 0 11868 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__C_N
timestamp 1688980957
transform 1 0 57592 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A1
timestamp 1688980957
transform -1 0 45632 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1688980957
transform 1 0 50968 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__B
timestamp 1688980957
transform 1 0 50600 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__B
timestamp 1688980957
transform 1 0 47656 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B
timestamp 1688980957
transform 1 0 41952 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__C
timestamp 1688980957
transform 1 0 41676 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A
timestamp 1688980957
transform 1 0 48024 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1688980957
transform 1 0 47196 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B
timestamp 1688980957
transform 1 0 46460 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A
timestamp 1688980957
transform 1 0 25760 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A3
timestamp 1688980957
transform 1 0 46276 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A
timestamp 1688980957
transform 1 0 15732 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__B
timestamp 1688980957
transform 1 0 39008 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A
timestamp 1688980957
transform -1 0 42780 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B
timestamp 1688980957
transform -1 0 41400 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B
timestamp 1688980957
transform -1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A
timestamp 1688980957
transform 1 0 52440 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1688980957
transform 1 0 51244 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B
timestamp 1688980957
transform 1 0 39192 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A2
timestamp 1688980957
transform -1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A
timestamp 1688980957
transform 1 0 40296 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A
timestamp 1688980957
transform -1 0 44160 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A
timestamp 1688980957
transform -1 0 45080 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1688980957
transform 1 0 45908 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__B
timestamp 1688980957
transform 1 0 46276 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__C
timestamp 1688980957
transform 1 0 45080 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A2
timestamp 1688980957
transform 1 0 43424 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A
timestamp 1688980957
transform 1 0 52440 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A
timestamp 1688980957
transform 1 0 52072 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A1
timestamp 1688980957
transform 1 0 46000 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A
timestamp 1688980957
transform -1 0 47012 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1688980957
transform -1 0 44068 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__C
timestamp 1688980957
transform 1 0 45724 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A
timestamp 1688980957
transform 1 0 52440 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A
timestamp 1688980957
transform 1 0 5980 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A
timestamp 1688980957
transform 1 0 6164 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A
timestamp 1688980957
transform 1 0 8004 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A
timestamp 1688980957
transform 1 0 4784 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__B1
timestamp 1688980957
transform 1 0 14260 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__B
timestamp 1688980957
transform 1 0 13800 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1688980957
transform 1 0 12420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__1_A
timestamp 1688980957
transform 1 0 39284 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A
timestamp 1688980957
transform 1 0 4876 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A
timestamp 1688980957
transform 1 0 6532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1688980957
transform 1 0 10028 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1688980957
transform -1 0 5336 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A
timestamp 1688980957
transform -1 0 7452 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A
timestamp 1688980957
transform 1 0 10580 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A
timestamp 1688980957
transform -1 0 3312 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A
timestamp 1688980957
transform 1 0 8648 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A
timestamp 1688980957
transform -1 0 4324 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A
timestamp 1688980957
transform -1 0 7084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A
timestamp 1688980957
transform 1 0 4048 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1688980957
transform 1 0 10856 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A
timestamp 1688980957
transform 1 0 8188 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A
timestamp 1688980957
transform 1 0 8556 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A
timestamp 1688980957
transform 1 0 12052 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B
timestamp 1688980957
transform 1 0 9568 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A2
timestamp 1688980957
transform 1 0 9936 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A
timestamp 1688980957
transform 1 0 10212 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A
timestamp 1688980957
transform 1 0 10764 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B
timestamp 1688980957
transform 1 0 6256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A2
timestamp 1688980957
transform 1 0 5888 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B
timestamp 1688980957
transform -1 0 7452 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A2
timestamp 1688980957
transform 1 0 7912 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__B
timestamp 1688980957
transform 1 0 13432 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A2
timestamp 1688980957
transform 1 0 12328 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B
timestamp 1688980957
transform -1 0 11132 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A2
timestamp 1688980957
transform 1 0 10120 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__B
timestamp 1688980957
transform -1 0 6900 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A2
timestamp 1688980957
transform 1 0 6716 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__B
timestamp 1688980957
transform 1 0 7912 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A2
timestamp 1688980957
transform 1 0 7636 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__B
timestamp 1688980957
transform -1 0 12972 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A2
timestamp 1688980957
transform 1 0 11868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1688980957
transform 1 0 5244 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__A
timestamp 1688980957
transform 1 0 8832 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__A
timestamp 1688980957
transform 1 0 9660 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__A
timestamp 1688980957
transform 1 0 9476 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A
timestamp 1688980957
transform 1 0 5244 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__A
timestamp 1688980957
transform 1 0 6532 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A
timestamp 1688980957
transform 1 0 9200 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A
timestamp 1688980957
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__A
timestamp 1688980957
transform 1 0 5060 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A
timestamp 1688980957
transform 1 0 7452 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1688980957
transform 1 0 9568 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__B1
timestamp 1688980957
transform 1 0 42872 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__A
timestamp 1688980957
transform 1 0 49588 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__B
timestamp 1688980957
transform 1 0 53360 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__B
timestamp 1688980957
transform 1 0 56028 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__B
timestamp 1688980957
transform 1 0 54924 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A
timestamp 1688980957
transform 1 0 56396 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__C
timestamp 1688980957
transform 1 0 57132 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A
timestamp 1688980957
transform 1 0 57684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__C
timestamp 1688980957
transform -1 0 57684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__B
timestamp 1688980957
transform 1 0 49588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__B
timestamp 1688980957
transform -1 0 50324 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__C1
timestamp 1688980957
transform -1 0 48484 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__S
timestamp 1688980957
transform -1 0 56396 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__C
timestamp 1688980957
transform 1 0 57776 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A
timestamp 1688980957
transform 1 0 57592 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__B
timestamp 1688980957
transform 1 0 57592 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__B1
timestamp 1688980957
transform 1 0 47564 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__B
timestamp 1688980957
transform 1 0 52532 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__B
timestamp 1688980957
transform 1 0 53360 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1235__B
timestamp 1688980957
transform 1 0 53084 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__B
timestamp 1688980957
transform -1 0 52900 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__B
timestamp 1688980957
transform -1 0 51244 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__B
timestamp 1688980957
transform 1 0 53820 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__B
timestamp 1688980957
transform 1 0 53268 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__B
timestamp 1688980957
transform 1 0 51152 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__C1
timestamp 1688980957
transform -1 0 51060 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__S
timestamp 1688980957
transform 1 0 57132 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__A
timestamp 1688980957
transform 1 0 56856 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__S
timestamp 1688980957
transform 1 0 56764 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1283__A
timestamp 1688980957
transform 1 0 48944 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__B
timestamp 1688980957
transform 1 0 56764 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1296__B
timestamp 1688980957
transform 1 0 57040 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__B
timestamp 1688980957
transform 1 0 56764 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1306__B
timestamp 1688980957
transform 1 0 56764 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__A
timestamp 1688980957
transform -1 0 57040 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__C
timestamp 1688980957
transform 1 0 56396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1314__A
timestamp 1688980957
transform 1 0 57040 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__C
timestamp 1688980957
transform 1 0 57316 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1323__B
timestamp 1688980957
transform 1 0 48852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__B
timestamp 1688980957
transform 1 0 49404 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__C1
timestamp 1688980957
transform 1 0 49680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__S
timestamp 1688980957
transform 1 0 55936 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__A1
timestamp 1688980957
transform 1 0 57592 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__B
timestamp 1688980957
transform 1 0 53084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__B
timestamp 1688980957
transform 1 0 54188 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__B
timestamp 1688980957
transform 1 0 53084 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__B
timestamp 1688980957
transform 1 0 52900 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__B
timestamp 1688980957
transform 1 0 54004 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__B
timestamp 1688980957
transform 1 0 52992 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__C
timestamp 1688980957
transform 1 0 54464 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__B
timestamp 1688980957
transform 1 0 53728 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__B
timestamp 1688980957
transform -1 0 51428 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__C1
timestamp 1688980957
transform 1 0 50048 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__S
timestamp 1688980957
transform 1 0 57040 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__S
timestamp 1688980957
transform 1 0 56764 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__S
timestamp 1688980957
transform -1 0 56764 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__A
timestamp 1688980957
transform 1 0 50048 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__C
timestamp 1688980957
transform 1 0 41952 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__B
timestamp 1688980957
transform -1 0 47472 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__A1
timestamp 1688980957
transform 1 0 48852 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__A1
timestamp 1688980957
transform 1 0 48668 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__A
timestamp 1688980957
transform 1 0 39192 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__A2
timestamp 1688980957
transform 1 0 38272 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1565__RESET_B
timestamp 1688980957
transform 1 0 44528 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1566__CLK
timestamp 1688980957
transform 1 0 37168 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1568__CLK
timestamp 1688980957
transform 1 0 40020 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1568__RESET_B
timestamp 1688980957
transform 1 0 42136 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1572__RESET_B
timestamp 1688980957
transform 1 0 43700 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1573__RESET_B
timestamp 1688980957
transform 1 0 43240 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1574__RESET_B
timestamp 1688980957
transform -1 0 46828 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__CLK
timestamp 1688980957
transform 1 0 8280 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1583__CLK
timestamp 1688980957
transform 1 0 10488 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1584__CLK
timestamp 1688980957
transform 1 0 6532 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1594__CLK
timestamp 1688980957
transform 1 0 12420 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1595__CLK
timestamp 1688980957
transform -1 0 14444 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1596__CLK
timestamp 1688980957
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1597__RESET_B
timestamp 1688980957
transform 1 0 42596 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1598__CLK
timestamp 1688980957
transform 1 0 13248 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1617__CLK
timestamp 1688980957
transform 1 0 11684 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1618__CLK
timestamp 1688980957
transform 1 0 12236 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1621__CLK
timestamp 1688980957
transform 1 0 12420 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1631__CLK
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1641__CLK
timestamp 1688980957
transform -1 0 11224 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1642__CLK
timestamp 1688980957
transform 1 0 9200 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1645__CLK
timestamp 1688980957
transform 1 0 10764 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1646__CLK
timestamp 1688980957
transform 1 0 40020 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1683__RESET_B
timestamp 1688980957
transform 1 0 47196 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1684__RESET_B
timestamp 1688980957
transform 1 0 48484 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1685__CLK
timestamp 1688980957
transform 1 0 36248 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1685__RESET_B
timestamp 1688980957
transform 1 0 38272 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1687__CLK
timestamp 1688980957
transform 1 0 36524 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1687__RESET_B
timestamp 1688980957
transform 1 0 39376 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1688__CLK
timestamp 1688980957
transform 1 0 34960 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1688__RESET_B
timestamp 1688980957
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1689__CLK
timestamp 1688980957
transform 1 0 35236 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1689__RESET_B
timestamp 1688980957
transform 1 0 37444 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1690__CLK
timestamp 1688980957
transform 1 0 37260 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1690__RESET_B
timestamp 1688980957
transform 1 0 39652 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1693__RESET_B
timestamp 1688980957
transform -1 0 46552 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1694__RESET_B
timestamp 1688980957
transform 1 0 48484 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1695__RESET_B
timestamp 1688980957
transform 1 0 48852 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1696__RESET_B
timestamp 1688980957
transform 1 0 47288 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_clk_i_A
timestamp 1688980957
transform 1 0 14260 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_clk_i_A
timestamp 1688980957
transform 1 0 20240 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_clk_i_A
timestamp 1688980957
transform -1 0 12604 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_clk_i_A
timestamp 1688980957
transform -1 0 17848 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_clk_i_A
timestamp 1688980957
transform -1 0 44160 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_clk_i_A
timestamp 1688980957
transform 1 0 49680 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_clk_i_A
timestamp 1688980957
transform 1 0 43976 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_clk_i_A
timestamp 1688980957
transform 1 0 49772 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout103_A
timestamp 1688980957
transform 1 0 12788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout104_A
timestamp 1688980957
transform -1 0 13340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout105_A
timestamp 1688980957
transform 1 0 11684 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout106_A
timestamp 1688980957
transform -1 0 44804 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_fanout107_A
timestamp 1688980957
transform 1 0 46184 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold85_A
timestamp 1688980957
transform 1 0 46092 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold88_A
timestamp 1688980957
transform 1 0 48944 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold156_A
timestamp 1688980957
transform 1 0 47012 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold215_A
timestamp 1688980957
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold234_A
timestamp 1688980957
transform -1 0 42964 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold241_A
timestamp 1688980957
transform -1 0 42412 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output63_A
timestamp 1688980957
transform 1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output64_A
timestamp 1688980957
transform 1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output65_A
timestamp 1688980957
transform 1 0 29164 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output66_A
timestamp 1688980957
transform 1 0 39100 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output68_A
timestamp 1688980957
transform 1 0 56120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output93_A
timestamp 1688980957
transform 1 0 3036 0 -1 54400
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1688980957
transform -1 0 3220 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output95_A
timestamp 1688980957
transform 1 0 3036 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29808 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk_i
timestamp 1688980957
transform -1 0 13800 0 1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk_i
timestamp 1688980957
transform 1 0 18216 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk_i
timestamp 1688980957
transform -1 0 12236 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk_i
timestamp 1688980957
transform 1 0 15640 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk_i
timestamp 1688980957
transform 1 0 44160 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk_i
timestamp 1688980957
transform 1 0 49404 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk_i
timestamp 1688980957
transform 1 0 44160 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk_i
timestamp 1688980957
transform 1 0 50140 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_4  fanout103
timestamp 1688980957
transform -1 0 13524 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout104
timestamp 1688980957
transform -1 0 12972 0 -1 20672
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout105
timestamp 1688980957
transform -1 0 11224 0 -1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout106
timestamp 1688980957
transform 1 0 43424 0 1 33728
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  fanout107
timestamp 1688980957
transform 1 0 46368 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_11 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_33 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_45
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_89
timestamp 1688980957
transform 1 0 9292 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_101
timestamp 1688980957
transform 1 0 10396 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_129
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_182
timestamp 1688980957
transform 1 0 17848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_194
timestamp 1688980957
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_243
timestamp 1688980957
transform 1 0 23460 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_281 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_303
timestamp 1688980957
transform 1 0 28980 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_337 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_345
timestamp 1688980957
transform 1 0 32844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_357
timestamp 1688980957
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_411
timestamp 1688980957
transform 1 0 38916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_415
timestamp 1688980957
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_419
timestamp 1688980957
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_453
timestamp 1688980957
transform 1 0 42780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_465
timestamp 1688980957
transform 1 0 43884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_473
timestamp 1688980957
transform 1 0 44620 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_477
timestamp 1688980957
transform 1 0 44988 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_489
timestamp 1688980957
transform 1 0 46092 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_501
timestamp 1688980957
transform 1 0 47196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_521
timestamp 1688980957
transform 1 0 49036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_529
timestamp 1688980957
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_533
timestamp 1688980957
transform 1 0 50140 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_545
timestamp 1688980957
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_557
timestamp 1688980957
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_565
timestamp 1688980957
transform 1 0 53084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_577
timestamp 1688980957
transform 1 0 54188 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_585
timestamp 1688980957
transform 1 0 54924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_589
timestamp 1688980957
transform 1 0 55292 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_597
timestamp 1688980957
transform 1 0 56028 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_617
timestamp 1688980957
transform 1 0 57868 0 1 2176
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_473
timestamp 1688980957
transform 1 0 44620 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_485
timestamp 1688980957
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_497
timestamp 1688980957
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_503
timestamp 1688980957
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_505
timestamp 1688980957
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_517
timestamp 1688980957
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_529
timestamp 1688980957
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_541
timestamp 1688980957
transform 1 0 50876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_553
timestamp 1688980957
transform 1 0 51980 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_559
timestamp 1688980957
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_561
timestamp 1688980957
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_573
timestamp 1688980957
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_585
timestamp 1688980957
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_597
timestamp 1688980957
transform 1 0 56028 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_609
timestamp 1688980957
transform 1 0 57132 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_615
timestamp 1688980957
transform 1 0 57684 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_617
timestamp 1688980957
transform 1 0 57868 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_19
timestamp 1688980957
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_469
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_475
timestamp 1688980957
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_477
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_489
timestamp 1688980957
transform 1 0 46092 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_501
timestamp 1688980957
transform 1 0 47196 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_513
timestamp 1688980957
transform 1 0 48300 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_525
timestamp 1688980957
transform 1 0 49404 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_531
timestamp 1688980957
transform 1 0 49956 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_533
timestamp 1688980957
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_545
timestamp 1688980957
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_557
timestamp 1688980957
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_569
timestamp 1688980957
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_581
timestamp 1688980957
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_587
timestamp 1688980957
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_589
timestamp 1688980957
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_601
timestamp 1688980957
transform 1 0 56396 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_613
timestamp 1688980957
transform 1 0 57500 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_473
timestamp 1688980957
transform 1 0 44620 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_485
timestamp 1688980957
transform 1 0 45724 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_497
timestamp 1688980957
transform 1 0 46828 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_503
timestamp 1688980957
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_505
timestamp 1688980957
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_517
timestamp 1688980957
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_529
timestamp 1688980957
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_541
timestamp 1688980957
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_553
timestamp 1688980957
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_559
timestamp 1688980957
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_561
timestamp 1688980957
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_573
timestamp 1688980957
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_585
timestamp 1688980957
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_597
timestamp 1688980957
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_609
timestamp 1688980957
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_615
timestamp 1688980957
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_617
timestamp 1688980957
transform 1 0 57868 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 1688980957
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1688980957
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_477
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_489
timestamp 1688980957
transform 1 0 46092 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_501
timestamp 1688980957
transform 1 0 47196 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_513
timestamp 1688980957
transform 1 0 48300 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_525
timestamp 1688980957
transform 1 0 49404 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_531
timestamp 1688980957
transform 1 0 49956 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_533
timestamp 1688980957
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_545
timestamp 1688980957
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_557
timestamp 1688980957
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_569
timestamp 1688980957
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_581
timestamp 1688980957
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_587
timestamp 1688980957
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_589
timestamp 1688980957
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_601
timestamp 1688980957
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_613
timestamp 1688980957
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_19
timestamp 1688980957
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_31
timestamp 1688980957
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_43
timestamp 1688980957
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_473
timestamp 1688980957
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_485
timestamp 1688980957
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_497
timestamp 1688980957
transform 1 0 46828 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_503
timestamp 1688980957
transform 1 0 47380 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_505
timestamp 1688980957
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_517
timestamp 1688980957
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_529
timestamp 1688980957
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_541
timestamp 1688980957
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_553
timestamp 1688980957
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_559
timestamp 1688980957
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_561
timestamp 1688980957
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_573
timestamp 1688980957
transform 1 0 53820 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_585
timestamp 1688980957
transform 1 0 54924 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_597
timestamp 1688980957
transform 1 0 56028 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_609
timestamp 1688980957
transform 1 0 57132 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_615
timestamp 1688980957
transform 1 0 57684 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_617
timestamp 1688980957
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_469
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 1688980957
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_489
timestamp 1688980957
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_501
timestamp 1688980957
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_513
timestamp 1688980957
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_525
timestamp 1688980957
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_531
timestamp 1688980957
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_533
timestamp 1688980957
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_545
timestamp 1688980957
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_557
timestamp 1688980957
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_569
timestamp 1688980957
transform 1 0 53452 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_581
timestamp 1688980957
transform 1 0 54556 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_587
timestamp 1688980957
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_589
timestamp 1688980957
transform 1 0 55292 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_601
timestamp 1688980957
transform 1 0 56396 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_613
timestamp 1688980957
transform 1 0 57500 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_473
timestamp 1688980957
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_485
timestamp 1688980957
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_497
timestamp 1688980957
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_503
timestamp 1688980957
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_505
timestamp 1688980957
transform 1 0 47564 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_517
timestamp 1688980957
transform 1 0 48668 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_529
timestamp 1688980957
transform 1 0 49772 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_541
timestamp 1688980957
transform 1 0 50876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_553
timestamp 1688980957
transform 1 0 51980 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_559
timestamp 1688980957
transform 1 0 52532 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_561
timestamp 1688980957
transform 1 0 52716 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_573
timestamp 1688980957
transform 1 0 53820 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_585
timestamp 1688980957
transform 1 0 54924 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_597
timestamp 1688980957
transform 1 0 56028 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_609
timestamp 1688980957
transform 1 0 57132 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_615
timestamp 1688980957
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_617
timestamp 1688980957
transform 1 0 57868 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_19
timestamp 1688980957
transform 1 0 2852 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 1688980957
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 1688980957
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_477
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_489
timestamp 1688980957
transform 1 0 46092 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_501
timestamp 1688980957
transform 1 0 47196 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_513
timestamp 1688980957
transform 1 0 48300 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_525
timestamp 1688980957
transform 1 0 49404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_531
timestamp 1688980957
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_533
timestamp 1688980957
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_545
timestamp 1688980957
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_557
timestamp 1688980957
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_569
timestamp 1688980957
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_581
timestamp 1688980957
transform 1 0 54556 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_587
timestamp 1688980957
transform 1 0 55108 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_589
timestamp 1688980957
transform 1 0 55292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_601
timestamp 1688980957
transform 1 0 56396 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_613
timestamp 1688980957
transform 1 0 57500 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_473
timestamp 1688980957
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_485
timestamp 1688980957
transform 1 0 45724 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_497
timestamp 1688980957
transform 1 0 46828 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_503
timestamp 1688980957
transform 1 0 47380 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_505
timestamp 1688980957
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_517
timestamp 1688980957
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_529
timestamp 1688980957
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_541
timestamp 1688980957
transform 1 0 50876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_553
timestamp 1688980957
transform 1 0 51980 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_559
timestamp 1688980957
transform 1 0 52532 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_561
timestamp 1688980957
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_573
timestamp 1688980957
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_585
timestamp 1688980957
transform 1 0 54924 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_597
timestamp 1688980957
transform 1 0 56028 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_609
timestamp 1688980957
transform 1 0 57132 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_615
timestamp 1688980957
transform 1 0 57684 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_617
timestamp 1688980957
transform 1 0 57868 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_621
timestamp 1688980957
transform 1 0 58236 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_469
timestamp 1688980957
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_475
timestamp 1688980957
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_477
timestamp 1688980957
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_489
timestamp 1688980957
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_501
timestamp 1688980957
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_513
timestamp 1688980957
transform 1 0 48300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_525
timestamp 1688980957
transform 1 0 49404 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_531
timestamp 1688980957
transform 1 0 49956 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_533
timestamp 1688980957
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_545
timestamp 1688980957
transform 1 0 51244 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_557
timestamp 1688980957
transform 1 0 52348 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_569
timestamp 1688980957
transform 1 0 53452 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_581
timestamp 1688980957
transform 1 0 54556 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_587
timestamp 1688980957
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_589
timestamp 1688980957
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_601
timestamp 1688980957
transform 1 0 56396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_613
timestamp 1688980957
transform 1 0 57500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_19
timestamp 1688980957
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_31
timestamp 1688980957
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_43
timestamp 1688980957
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 1688980957
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_461
timestamp 1688980957
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_473
timestamp 1688980957
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_485
timestamp 1688980957
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_497
timestamp 1688980957
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_503
timestamp 1688980957
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_505
timestamp 1688980957
transform 1 0 47564 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_517
timestamp 1688980957
transform 1 0 48668 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_529
timestamp 1688980957
transform 1 0 49772 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_541
timestamp 1688980957
transform 1 0 50876 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_553
timestamp 1688980957
transform 1 0 51980 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_559
timestamp 1688980957
transform 1 0 52532 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_561
timestamp 1688980957
transform 1 0 52716 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_573
timestamp 1688980957
transform 1 0 53820 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_585
timestamp 1688980957
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_597
timestamp 1688980957
transform 1 0 56028 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_609
timestamp 1688980957
transform 1 0 57132 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_615
timestamp 1688980957
transform 1 0 57684 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_617
timestamp 1688980957
transform 1 0 57868 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_621
timestamp 1688980957
transform 1 0 58236 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 1688980957
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 1688980957
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 1688980957
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 1688980957
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 1688980957
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 1688980957
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 1688980957
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 1688980957
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_221
timestamp 1688980957
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_233
timestamp 1688980957
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_253
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_265
timestamp 1688980957
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_289
timestamp 1688980957
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1688980957
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_457
timestamp 1688980957
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_469
timestamp 1688980957
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_475
timestamp 1688980957
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_477
timestamp 1688980957
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_489
timestamp 1688980957
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_501
timestamp 1688980957
transform 1 0 47196 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_513
timestamp 1688980957
transform 1 0 48300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_525
timestamp 1688980957
transform 1 0 49404 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_531
timestamp 1688980957
transform 1 0 49956 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_533
timestamp 1688980957
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_545
timestamp 1688980957
transform 1 0 51244 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_557
timestamp 1688980957
transform 1 0 52348 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_569
timestamp 1688980957
transform 1 0 53452 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_581
timestamp 1688980957
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_587
timestamp 1688980957
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_589
timestamp 1688980957
transform 1 0 55292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_601
timestamp 1688980957
transform 1 0 56396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_613
timestamp 1688980957
transform 1 0 57500 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_621
timestamp 1688980957
transform 1 0 58236 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 1688980957
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 1688980957
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 1688980957
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 1688980957
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 1688980957
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 1688980957
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 1688980957
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1688980957
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_237
timestamp 1688980957
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_261
timestamp 1688980957
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_273
timestamp 1688980957
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_279
timestamp 1688980957
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 1688980957
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_305
timestamp 1688980957
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_317
timestamp 1688980957
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_335
timestamp 1688980957
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 1688980957
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 1688980957
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_361
timestamp 1688980957
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 1688980957
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 1688980957
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 1688980957
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_405
timestamp 1688980957
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_417
timestamp 1688980957
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_429
timestamp 1688980957
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_441
timestamp 1688980957
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1688980957
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_449
timestamp 1688980957
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_461
timestamp 1688980957
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_473
timestamp 1688980957
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_485
timestamp 1688980957
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_497
timestamp 1688980957
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_503
timestamp 1688980957
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_505
timestamp 1688980957
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_517
timestamp 1688980957
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_529
timestamp 1688980957
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_541
timestamp 1688980957
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_553
timestamp 1688980957
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_559
timestamp 1688980957
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_561
timestamp 1688980957
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_573
timestamp 1688980957
transform 1 0 53820 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_585
timestamp 1688980957
transform 1 0 54924 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_597
timestamp 1688980957
transform 1 0 56028 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_609
timestamp 1688980957
transform 1 0 57132 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_615
timestamp 1688980957
transform 1 0 57684 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_617
timestamp 1688980957
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_19
timestamp 1688980957
transform 1 0 2852 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 1688980957
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 1688980957
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 1688980957
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 1688980957
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 1688980957
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 1688980957
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 1688980957
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_209
timestamp 1688980957
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_221
timestamp 1688980957
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_233
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_245
timestamp 1688980957
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_289
timestamp 1688980957
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_301
timestamp 1688980957
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 1688980957
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_321
timestamp 1688980957
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_333
timestamp 1688980957
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_345
timestamp 1688980957
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_357
timestamp 1688980957
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_363
timestamp 1688980957
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1688980957
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 1688980957
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_401
timestamp 1688980957
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_413
timestamp 1688980957
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_419
timestamp 1688980957
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_421
timestamp 1688980957
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_433
timestamp 1688980957
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_445
timestamp 1688980957
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_457
timestamp 1688980957
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_469
timestamp 1688980957
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_475
timestamp 1688980957
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_477
timestamp 1688980957
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_489
timestamp 1688980957
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_501
timestamp 1688980957
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_513
timestamp 1688980957
transform 1 0 48300 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_525
timestamp 1688980957
transform 1 0 49404 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_531
timestamp 1688980957
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_533
timestamp 1688980957
transform 1 0 50140 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_545
timestamp 1688980957
transform 1 0 51244 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_557
timestamp 1688980957
transform 1 0 52348 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_569
timestamp 1688980957
transform 1 0 53452 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_581
timestamp 1688980957
transform 1 0 54556 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_587
timestamp 1688980957
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_589
timestamp 1688980957
transform 1 0 55292 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_601
timestamp 1688980957
transform 1 0 56396 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_613
timestamp 1688980957
transform 1 0 57500 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_621
timestamp 1688980957
transform 1 0 58236 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 1688980957
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 1688980957
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 1688980957
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 1688980957
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 1688980957
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 1688980957
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 1688980957
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 1688980957
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_217
timestamp 1688980957
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_223
timestamp 1688980957
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_225
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_237
timestamp 1688980957
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_249
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_261
timestamp 1688980957
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_273
timestamp 1688980957
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_279
timestamp 1688980957
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 1688980957
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_305
timestamp 1688980957
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_317
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_329
timestamp 1688980957
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_335
timestamp 1688980957
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 1688980957
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 1688980957
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_361
timestamp 1688980957
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_373
timestamp 1688980957
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_385
timestamp 1688980957
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 1688980957
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_405
timestamp 1688980957
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_417
timestamp 1688980957
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_429
timestamp 1688980957
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_441
timestamp 1688980957
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_447
timestamp 1688980957
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_449
timestamp 1688980957
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_461
timestamp 1688980957
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_473
timestamp 1688980957
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_485
timestamp 1688980957
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_497
timestamp 1688980957
transform 1 0 46828 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_503
timestamp 1688980957
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_505
timestamp 1688980957
transform 1 0 47564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_517
timestamp 1688980957
transform 1 0 48668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_521
timestamp 1688980957
transform 1 0 49036 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_525
timestamp 1688980957
transform 1 0 49404 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_537
timestamp 1688980957
transform 1 0 50508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_549
timestamp 1688980957
transform 1 0 51612 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_557
timestamp 1688980957
transform 1 0 52348 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_561
timestamp 1688980957
transform 1 0 52716 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_573
timestamp 1688980957
transform 1 0 53820 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_585
timestamp 1688980957
transform 1 0 54924 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_597
timestamp 1688980957
transform 1 0 56028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_609
timestamp 1688980957
transform 1 0 57132 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_615
timestamp 1688980957
transform 1 0 57684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_617
timestamp 1688980957
transform 1 0 57868 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_621
timestamp 1688980957
transform 1 0 58236 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 1688980957
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 1688980957
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 1688980957
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 1688980957
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 1688980957
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 1688980957
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 1688980957
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 1688980957
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 1688980957
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 1688980957
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_221
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_233
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_245
timestamp 1688980957
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 1688980957
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 1688980957
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_289
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_301
timestamp 1688980957
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_307
timestamp 1688980957
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_333
timestamp 1688980957
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_345
timestamp 1688980957
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_357
timestamp 1688980957
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 1688980957
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 1688980957
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_389
timestamp 1688980957
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_401
timestamp 1688980957
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_413
timestamp 1688980957
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_419
timestamp 1688980957
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_421
timestamp 1688980957
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_433
timestamp 1688980957
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_445
timestamp 1688980957
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_457
timestamp 1688980957
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_469
timestamp 1688980957
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_475
timestamp 1688980957
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_477
timestamp 1688980957
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_489
timestamp 1688980957
transform 1 0 46092 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_501
timestamp 1688980957
transform 1 0 47196 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_513
timestamp 1688980957
transform 1 0 48300 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_525
timestamp 1688980957
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_531
timestamp 1688980957
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_533
timestamp 1688980957
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_545
timestamp 1688980957
transform 1 0 51244 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_557
timestamp 1688980957
transform 1 0 52348 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_569
timestamp 1688980957
transform 1 0 53452 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_581
timestamp 1688980957
transform 1 0 54556 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_587
timestamp 1688980957
transform 1 0 55108 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_589
timestamp 1688980957
transform 1 0 55292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_601
timestamp 1688980957
transform 1 0 56396 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_613
timestamp 1688980957
transform 1 0 57500 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_19
timestamp 1688980957
transform 1 0 2852 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_31
timestamp 1688980957
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_43
timestamp 1688980957
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 1688980957
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 1688980957
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 1688980957
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 1688980957
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1688980957
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1688980957
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 1688980957
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_293
timestamp 1688980957
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_305
timestamp 1688980957
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_317
timestamp 1688980957
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_329
timestamp 1688980957
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_335
timestamp 1688980957
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 1688980957
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_361
timestamp 1688980957
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_373
timestamp 1688980957
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_385
timestamp 1688980957
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 1688980957
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_405
timestamp 1688980957
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_417
timestamp 1688980957
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_429
timestamp 1688980957
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_441
timestamp 1688980957
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_447
timestamp 1688980957
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_449
timestamp 1688980957
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_461
timestamp 1688980957
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_473
timestamp 1688980957
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_485
timestamp 1688980957
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_497
timestamp 1688980957
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_503
timestamp 1688980957
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_505
timestamp 1688980957
transform 1 0 47564 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_517
timestamp 1688980957
transform 1 0 48668 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_525
timestamp 1688980957
transform 1 0 49404 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_536
timestamp 1688980957
transform 1 0 50416 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_548
timestamp 1688980957
transform 1 0 51520 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_561
timestamp 1688980957
transform 1 0 52716 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_573
timestamp 1688980957
transform 1 0 53820 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_585
timestamp 1688980957
transform 1 0 54924 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_597
timestamp 1688980957
transform 1 0 56028 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_609
timestamp 1688980957
transform 1 0 57132 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_615
timestamp 1688980957
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_623
timestamp 1688980957
transform 1 0 58420 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 1688980957
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 1688980957
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 1688980957
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 1688980957
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 1688980957
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 1688980957
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 1688980957
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 1688980957
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1688980957
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1688980957
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 1688980957
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_177
timestamp 1688980957
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_189
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 1688980957
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 1688980957
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 1688980957
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 1688980957
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 1688980957
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 1688980957
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_289
timestamp 1688980957
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_301
timestamp 1688980957
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 1688980957
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 1688980957
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 1688980957
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 1688980957
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1688980957
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1688980957
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_401
timestamp 1688980957
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_413
timestamp 1688980957
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_419
timestamp 1688980957
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_421
timestamp 1688980957
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_433
timestamp 1688980957
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_445
timestamp 1688980957
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_457
timestamp 1688980957
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_469
timestamp 1688980957
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_475
timestamp 1688980957
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_477
timestamp 1688980957
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_489
timestamp 1688980957
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_501
timestamp 1688980957
transform 1 0 47196 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_509
timestamp 1688980957
transform 1 0 47932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_531
timestamp 1688980957
transform 1 0 49956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_533
timestamp 1688980957
transform 1 0 50140 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_550
timestamp 1688980957
transform 1 0 51704 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_556
timestamp 1688980957
transform 1 0 52256 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_568
timestamp 1688980957
transform 1 0 53360 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_600
timestamp 1688980957
transform 1 0 56304 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_604
timestamp 1688980957
transform 1 0 56672 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_616
timestamp 1688980957
transform 1 0 57776 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_623
timestamp 1688980957
transform 1 0 58420 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 1688980957
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 1688980957
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 1688980957
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 1688980957
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 1688980957
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 1688980957
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 1688980957
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 1688980957
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 1688980957
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 1688980957
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 1688980957
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_193
timestamp 1688980957
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_205
timestamp 1688980957
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_217
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 1688980957
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 1688980957
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 1688980957
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 1688980957
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 1688980957
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_305
timestamp 1688980957
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_317
timestamp 1688980957
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_329
timestamp 1688980957
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1688980957
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1688980957
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 1688980957
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 1688980957
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 1688980957
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 1688980957
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_405
timestamp 1688980957
transform 1 0 38364 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_417
timestamp 1688980957
transform 1 0 39468 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_429
timestamp 1688980957
transform 1 0 40572 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_441
timestamp 1688980957
transform 1 0 41676 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_447
timestamp 1688980957
transform 1 0 42228 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_449
timestamp 1688980957
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_461
timestamp 1688980957
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_473
timestamp 1688980957
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_485
timestamp 1688980957
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_501
timestamp 1688980957
transform 1 0 47196 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_505
timestamp 1688980957
transform 1 0 47564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_510
timestamp 1688980957
transform 1 0 48024 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_518
timestamp 1688980957
transform 1 0 48760 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_533
timestamp 1688980957
transform 1 0 50140 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_539
timestamp 1688980957
transform 1 0 50692 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_546
timestamp 1688980957
transform 1 0 51336 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_555
timestamp 1688980957
transform 1 0 52164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_584
timestamp 1688980957
transform 1 0 54832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_594
timestamp 1688980957
transform 1 0 55752 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_598
timestamp 1688980957
transform 1 0 56120 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_615
timestamp 1688980957
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_19
timestamp 1688980957
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 1688980957
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 1688980957
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1688980957
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1688980957
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1688980957
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 1688980957
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 1688980957
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 1688980957
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 1688980957
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 1688980957
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 1688980957
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 1688980957
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 1688980957
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 1688980957
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 1688980957
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 1688980957
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_289
timestamp 1688980957
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_301
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 1688980957
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 1688980957
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 1688980957
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 1688980957
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 1688980957
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1688980957
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 1688980957
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 1688980957
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_401
timestamp 1688980957
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_413
timestamp 1688980957
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_419
timestamp 1688980957
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_421
timestamp 1688980957
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_433
timestamp 1688980957
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_445
timestamp 1688980957
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_457
timestamp 1688980957
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_469
timestamp 1688980957
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_475
timestamp 1688980957
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_477
timestamp 1688980957
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_489
timestamp 1688980957
transform 1 0 46092 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_523
timestamp 1688980957
transform 1 0 49220 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_527
timestamp 1688980957
transform 1 0 49588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_531
timestamp 1688980957
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_533
timestamp 1688980957
transform 1 0 50140 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_571
timestamp 1688980957
transform 1 0 53636 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_575
timestamp 1688980957
transform 1 0 54004 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_579
timestamp 1688980957
transform 1 0 54372 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_583
timestamp 1688980957
transform 1 0 54740 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_587
timestamp 1688980957
transform 1 0 55108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_589
timestamp 1688980957
transform 1 0 55292 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_597
timestamp 1688980957
transform 1 0 56028 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_604
timestamp 1688980957
transform 1 0 56672 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_608
timestamp 1688980957
transform 1 0 57040 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_620
timestamp 1688980957
transform 1 0 58144 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 1688980957
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 1688980957
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 1688980957
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1688980957
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1688980957
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 1688980957
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 1688980957
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 1688980957
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1688980957
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 1688980957
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 1688980957
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 1688980957
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 1688980957
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 1688980957
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 1688980957
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_293
timestamp 1688980957
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_305
timestamp 1688980957
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_317
timestamp 1688980957
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_329
timestamp 1688980957
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_335
timestamp 1688980957
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 1688980957
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_361
timestamp 1688980957
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_373
timestamp 1688980957
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_385
timestamp 1688980957
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 1688980957
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_405
timestamp 1688980957
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_417
timestamp 1688980957
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_429
timestamp 1688980957
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_441
timestamp 1688980957
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_447
timestamp 1688980957
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_449
timestamp 1688980957
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_461
timestamp 1688980957
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_473
timestamp 1688980957
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_485
timestamp 1688980957
transform 1 0 45724 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_497
timestamp 1688980957
transform 1 0 46828 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_503
timestamp 1688980957
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_515
timestamp 1688980957
transform 1 0 48484 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_525
timestamp 1688980957
transform 1 0 49404 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_537
timestamp 1688980957
transform 1 0 50508 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_541
timestamp 1688980957
transform 1 0 50876 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_552
timestamp 1688980957
transform 1 0 51888 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_567
timestamp 1688980957
transform 1 0 53268 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_580
timestamp 1688980957
transform 1 0 54464 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_588
timestamp 1688980957
transform 1 0 55200 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_606
timestamp 1688980957
transform 1 0 56856 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_614
timestamp 1688980957
transform 1 0 57592 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_617
timestamp 1688980957
transform 1 0 57868 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1688980957
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 1688980957
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 1688980957
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 1688980957
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 1688980957
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 1688980957
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 1688980957
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 1688980957
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 1688980957
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1688980957
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1688980957
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 1688980957
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 1688980957
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 1688980957
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1688980957
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1688980957
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 1688980957
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 1688980957
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 1688980957
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 1688980957
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 1688980957
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 1688980957
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_401
timestamp 1688980957
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_413
timestamp 1688980957
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_419
timestamp 1688980957
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_421
timestamp 1688980957
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_433
timestamp 1688980957
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_445
timestamp 1688980957
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_457
timestamp 1688980957
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_469
timestamp 1688980957
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_475
timestamp 1688980957
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_477
timestamp 1688980957
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_489
timestamp 1688980957
transform 1 0 46092 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_501
timestamp 1688980957
transform 1 0 47196 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_518
timestamp 1688980957
transform 1 0 48760 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_525
timestamp 1688980957
transform 1 0 49404 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_531
timestamp 1688980957
transform 1 0 49956 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_533
timestamp 1688980957
transform 1 0 50140 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_539
timestamp 1688980957
transform 1 0 50692 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_543
timestamp 1688980957
transform 1 0 51060 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_555
timestamp 1688980957
transform 1 0 52164 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_559
timestamp 1688980957
transform 1 0 52532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_571
timestamp 1688980957
transform 1 0 53636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_583
timestamp 1688980957
transform 1 0 54740 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_605
timestamp 1688980957
transform 1 0 56764 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_19
timestamp 1688980957
transform 1 0 2852 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_31
timestamp 1688980957
transform 1 0 3956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_43
timestamp 1688980957
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 1688980957
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 1688980957
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 1688980957
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 1688980957
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 1688980957
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 1688980957
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 1688980957
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 1688980957
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1688980957
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1688980957
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 1688980957
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 1688980957
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 1688980957
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 1688980957
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 1688980957
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 1688980957
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 1688980957
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 1688980957
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 1688980957
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 1688980957
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 1688980957
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_361
timestamp 1688980957
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_373
timestamp 1688980957
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_385
timestamp 1688980957
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 1688980957
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_405
timestamp 1688980957
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_417
timestamp 1688980957
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_429
timestamp 1688980957
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_441
timestamp 1688980957
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_447
timestamp 1688980957
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_449
timestamp 1688980957
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_461
timestamp 1688980957
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_473
timestamp 1688980957
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_485
timestamp 1688980957
transform 1 0 45724 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_493
timestamp 1688980957
transform 1 0 46460 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_498
timestamp 1688980957
transform 1 0 46920 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_509
timestamp 1688980957
transform 1 0 47932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_514
timestamp 1688980957
transform 1 0 48392 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_526
timestamp 1688980957
transform 1 0 49496 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_530
timestamp 1688980957
transform 1 0 49864 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_534
timestamp 1688980957
transform 1 0 50232 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_546
timestamp 1688980957
transform 1 0 51336 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_550
timestamp 1688980957
transform 1 0 51704 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_558
timestamp 1688980957
transform 1 0 52440 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_567
timestamp 1688980957
transform 1 0 53268 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_573
timestamp 1688980957
transform 1 0 53820 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_579
timestamp 1688980957
transform 1 0 54372 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_599
timestamp 1688980957
transform 1 0 56212 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_605
timestamp 1688980957
transform 1 0 56764 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 1688980957
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 1688980957
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 1688980957
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 1688980957
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 1688980957
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 1688980957
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 1688980957
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 1688980957
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 1688980957
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 1688980957
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 1688980957
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 1688980957
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 1688980957
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 1688980957
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 1688980957
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 1688980957
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_289
timestamp 1688980957
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1688980957
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1688980957
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 1688980957
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 1688980957
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 1688980957
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 1688980957
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 1688980957
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 1688980957
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 1688980957
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_401
timestamp 1688980957
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_413
timestamp 1688980957
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_419
timestamp 1688980957
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_421
timestamp 1688980957
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_433
timestamp 1688980957
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_445
timestamp 1688980957
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_457
timestamp 1688980957
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_469
timestamp 1688980957
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_475
timestamp 1688980957
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_477
timestamp 1688980957
transform 1 0 44988 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_485
timestamp 1688980957
transform 1 0 45724 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_520
timestamp 1688980957
transform 1 0 48944 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_529
timestamp 1688980957
transform 1 0 49772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_533
timestamp 1688980957
transform 1 0 50140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_542
timestamp 1688980957
transform 1 0 50968 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_548
timestamp 1688980957
transform 1 0 51520 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_553
timestamp 1688980957
transform 1 0 51980 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_557
timestamp 1688980957
transform 1 0 52348 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_561
timestamp 1688980957
transform 1 0 52716 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_567
timestamp 1688980957
transform 1 0 53268 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_574
timestamp 1688980957
transform 1 0 53912 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_586
timestamp 1688980957
transform 1 0 55016 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_593
timestamp 1688980957
transform 1 0 55660 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_606
timestamp 1688980957
transform 1 0 56856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_611
timestamp 1688980957
transform 1 0 57316 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_616
timestamp 1688980957
transform 1 0 57776 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_623
timestamp 1688980957
transform 1 0 58420 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 1688980957
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 1688980957
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 1688980957
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_65
timestamp 1688980957
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_73
timestamp 1688980957
transform 1 0 7820 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_82
timestamp 1688980957
transform 1 0 8648 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_94
timestamp 1688980957
transform 1 0 9752 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_106
timestamp 1688980957
transform 1 0 10856 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1688980957
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 1688980957
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 1688980957
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 1688980957
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 1688980957
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 1688980957
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 1688980957
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 1688980957
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 1688980957
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 1688980957
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 1688980957
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 1688980957
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 1688980957
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_361
timestamp 1688980957
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_373
timestamp 1688980957
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_385
timestamp 1688980957
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 1688980957
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_405
timestamp 1688980957
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_417
timestamp 1688980957
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_429
timestamp 1688980957
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_441
timestamp 1688980957
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_447
timestamp 1688980957
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_449
timestamp 1688980957
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_461
timestamp 1688980957
transform 1 0 43516 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_465
timestamp 1688980957
transform 1 0 43884 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_488
timestamp 1688980957
transform 1 0 46000 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_500
timestamp 1688980957
transform 1 0 47104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_505
timestamp 1688980957
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_511
timestamp 1688980957
transform 1 0 48116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_517
timestamp 1688980957
transform 1 0 48668 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_525
timestamp 1688980957
transform 1 0 49404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_529
timestamp 1688980957
transform 1 0 49772 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_546
timestamp 1688980957
transform 1 0 51336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_557
timestamp 1688980957
transform 1 0 52348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_561
timestamp 1688980957
transform 1 0 52716 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_565
timestamp 1688980957
transform 1 0 53084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_569
timestamp 1688980957
transform 1 0 53452 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_573
timestamp 1688980957
transform 1 0 53820 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_580
timestamp 1688980957
transform 1 0 54464 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_586
timestamp 1688980957
transform 1 0 55016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_615
timestamp 1688980957
transform 1 0 57684 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_623
timestamp 1688980957
transform 1 0 58420 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_26
timestamp 1688980957
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_32
timestamp 1688980957
transform 1 0 4048 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_58
timestamp 1688980957
transform 1 0 6440 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_81
timestamp 1688980957
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_106
timestamp 1688980957
transform 1 0 10856 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_118
timestamp 1688980957
transform 1 0 11960 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_130
timestamp 1688980957
transform 1 0 13064 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1688980957
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 1688980957
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 1688980957
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 1688980957
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 1688980957
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 1688980957
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 1688980957
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 1688980957
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 1688980957
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 1688980957
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 1688980957
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 1688980957
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 1688980957
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 1688980957
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 1688980957
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 1688980957
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 1688980957
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 1688980957
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 1688980957
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 1688980957
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 1688980957
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_401
timestamp 1688980957
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_413
timestamp 1688980957
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_419
timestamp 1688980957
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_421
timestamp 1688980957
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_433
timestamp 1688980957
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_445
timestamp 1688980957
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_457
timestamp 1688980957
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_469
timestamp 1688980957
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_475
timestamp 1688980957
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_477
timestamp 1688980957
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_489
timestamp 1688980957
transform 1 0 46092 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_511
timestamp 1688980957
transform 1 0 48116 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_521
timestamp 1688980957
transform 1 0 49036 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_527
timestamp 1688980957
transform 1 0 49588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_570
timestamp 1688980957
transform 1 0 53544 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_575
timestamp 1688980957
transform 1 0 54004 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_579
timestamp 1688980957
transform 1 0 54372 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_587
timestamp 1688980957
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_589
timestamp 1688980957
transform 1 0 55292 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_593
timestamp 1688980957
transform 1 0 55660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_611
timestamp 1688980957
transform 1 0 57316 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_621
timestamp 1688980957
transform 1 0 58236 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_11
timestamp 1688980957
transform 1 0 2116 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_34
timestamp 1688980957
transform 1 0 4232 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_97
timestamp 1688980957
transform 1 0 10028 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_110
timestamp 1688980957
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1688980957
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 1688980957
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 1688980957
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 1688980957
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 1688980957
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 1688980957
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 1688980957
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 1688980957
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 1688980957
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 1688980957
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 1688980957
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 1688980957
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 1688980957
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 1688980957
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 1688980957
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 1688980957
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_361
timestamp 1688980957
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_373
timestamp 1688980957
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_385
timestamp 1688980957
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1688980957
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_405
timestamp 1688980957
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_417
timestamp 1688980957
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_429
timestamp 1688980957
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_441
timestamp 1688980957
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_447
timestamp 1688980957
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_449
timestamp 1688980957
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_461
timestamp 1688980957
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_473
timestamp 1688980957
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_485
timestamp 1688980957
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_497
timestamp 1688980957
transform 1 0 46828 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_502
timestamp 1688980957
transform 1 0 47288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_508
timestamp 1688980957
transform 1 0 47840 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_527
timestamp 1688980957
transform 1 0 49588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_539
timestamp 1688980957
transform 1 0 50692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_551
timestamp 1688980957
transform 1 0 51796 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_559
timestamp 1688980957
transform 1 0 52532 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_561
timestamp 1688980957
transform 1 0 52716 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_567
timestamp 1688980957
transform 1 0 53268 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_579
timestamp 1688980957
transform 1 0 54372 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_591
timestamp 1688980957
transform 1 0 55476 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_603
timestamp 1688980957
transform 1 0 56580 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_607
timestamp 1688980957
transform 1 0 56948 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_611
timestamp 1688980957
transform 1 0 57316 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_615
timestamp 1688980957
transform 1 0 57684 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_617
timestamp 1688980957
transform 1 0 57868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_621
timestamp 1688980957
transform 1 0 58236 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1688980957
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_56
timestamp 1688980957
transform 1 0 6256 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_68
timestamp 1688980957
transform 1 0 7360 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_76
timestamp 1688980957
transform 1 0 8096 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 1688980957
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_88
timestamp 1688980957
transform 1 0 9200 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_119
timestamp 1688980957
transform 1 0 12052 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_123
timestamp 1688980957
transform 1 0 12420 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_135
timestamp 1688980957
transform 1 0 13524 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 1688980957
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 1688980957
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 1688980957
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 1688980957
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 1688980957
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 1688980957
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 1688980957
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 1688980957
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 1688980957
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 1688980957
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 1688980957
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 1688980957
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 1688980957
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 1688980957
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 1688980957
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 1688980957
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 1688980957
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 1688980957
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 1688980957
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_401
timestamp 1688980957
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_413
timestamp 1688980957
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_419
timestamp 1688980957
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_421
timestamp 1688980957
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_433
timestamp 1688980957
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_445
timestamp 1688980957
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_457
timestamp 1688980957
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_469
timestamp 1688980957
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_475
timestamp 1688980957
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_477
timestamp 1688980957
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_489
timestamp 1688980957
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_501
timestamp 1688980957
transform 1 0 47196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_510
timestamp 1688980957
transform 1 0 48024 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_526
timestamp 1688980957
transform 1 0 49496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_530
timestamp 1688980957
transform 1 0 49864 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_536
timestamp 1688980957
transform 1 0 50416 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_548
timestamp 1688980957
transform 1 0 51520 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_560
timestamp 1688980957
transform 1 0 52624 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_564
timestamp 1688980957
transform 1 0 52992 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_577
timestamp 1688980957
transform 1 0 54188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_583
timestamp 1688980957
transform 1 0 54740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_623
timestamp 1688980957
transform 1 0 58420 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_19
timestamp 1688980957
transform 1 0 2852 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_82
timestamp 1688980957
transform 1 0 8648 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_90
timestamp 1688980957
transform 1 0 9384 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_96
timestamp 1688980957
transform 1 0 9936 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_106
timestamp 1688980957
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_121
timestamp 1688980957
transform 1 0 12236 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_133
timestamp 1688980957
transform 1 0 13340 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_145
timestamp 1688980957
transform 1 0 14444 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_157
timestamp 1688980957
transform 1 0 15548 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_165
timestamp 1688980957
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 1688980957
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1688980957
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 1688980957
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 1688980957
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 1688980957
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 1688980957
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 1688980957
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 1688980957
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 1688980957
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 1688980957
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_361
timestamp 1688980957
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_373
timestamp 1688980957
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_385
timestamp 1688980957
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_391
timestamp 1688980957
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_405
timestamp 1688980957
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_417
timestamp 1688980957
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_429
timestamp 1688980957
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_441
timestamp 1688980957
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_447
timestamp 1688980957
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_449
timestamp 1688980957
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_461
timestamp 1688980957
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_473
timestamp 1688980957
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_485
timestamp 1688980957
transform 1 0 45724 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_502
timestamp 1688980957
transform 1 0 47288 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_516
timestamp 1688980957
transform 1 0 48576 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_557
timestamp 1688980957
transform 1 0 52348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_561
timestamp 1688980957
transform 1 0 52716 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_566
timestamp 1688980957
transform 1 0 53176 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_570
timestamp 1688980957
transform 1 0 53544 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_583
timestamp 1688980957
transform 1 0 54740 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_591
timestamp 1688980957
transform 1 0 55476 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_597
timestamp 1688980957
transform 1 0 56028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_609
timestamp 1688980957
transform 1 0 57132 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_621
timestamp 1688980957
transform 1 0 58236 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_3
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_15
timestamp 1688980957
transform 1 0 2484 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_91
timestamp 1688980957
transform 1 0 9476 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_96
timestamp 1688980957
transform 1 0 9936 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_110
timestamp 1688980957
transform 1 0 11224 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_122
timestamp 1688980957
transform 1 0 12328 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_134
timestamp 1688980957
transform 1 0 13432 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 1688980957
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 1688980957
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 1688980957
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 1688980957
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 1688980957
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1688980957
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 1688980957
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 1688980957
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 1688980957
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1688980957
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 1688980957
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_389
timestamp 1688980957
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_401
timestamp 1688980957
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_413
timestamp 1688980957
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_419
timestamp 1688980957
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_421
timestamp 1688980957
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_433
timestamp 1688980957
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_445
timestamp 1688980957
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_457
timestamp 1688980957
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_469
timestamp 1688980957
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_475
timestamp 1688980957
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_477
timestamp 1688980957
transform 1 0 44988 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_483
timestamp 1688980957
transform 1 0 45540 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_503
timestamp 1688980957
transform 1 0 47380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_521
timestamp 1688980957
transform 1 0 49036 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_530
timestamp 1688980957
transform 1 0 49864 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_539
timestamp 1688980957
transform 1 0 50692 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_547
timestamp 1688980957
transform 1 0 51428 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_551
timestamp 1688980957
transform 1 0 51796 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_586
timestamp 1688980957
transform 1 0 55016 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_589
timestamp 1688980957
transform 1 0 55292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_601
timestamp 1688980957
transform 1 0 56396 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_607
timestamp 1688980957
transform 1 0 56948 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_616
timestamp 1688980957
transform 1 0 57776 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_620
timestamp 1688980957
transform 1 0 58144 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_34
timestamp 1688980957
transform 1 0 4232 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_46
timestamp 1688980957
transform 1 0 5336 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_54
timestamp 1688980957
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_79
timestamp 1688980957
transform 1 0 8372 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_110
timestamp 1688980957
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_117
timestamp 1688980957
transform 1 0 11868 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_129
timestamp 1688980957
transform 1 0 12972 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_141
timestamp 1688980957
transform 1 0 14076 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_153
timestamp 1688980957
transform 1 0 15180 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_165
timestamp 1688980957
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 1688980957
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 1688980957
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 1688980957
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 1688980957
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 1688980957
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 1688980957
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 1688980957
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 1688980957
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 1688980957
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1688980957
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 1688980957
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 1688980957
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 1688980957
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_373
timestamp 1688980957
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_385
timestamp 1688980957
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 1688980957
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_405
timestamp 1688980957
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_417
timestamp 1688980957
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_429
timestamp 1688980957
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_441
timestamp 1688980957
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_447
timestamp 1688980957
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_449
timestamp 1688980957
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_461
timestamp 1688980957
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_473
timestamp 1688980957
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_485
timestamp 1688980957
transform 1 0 45724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_497
timestamp 1688980957
transform 1 0 46828 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_521
timestamp 1688980957
transform 1 0 49036 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_531
timestamp 1688980957
transform 1 0 49956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_538
timestamp 1688980957
transform 1 0 50600 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_553
timestamp 1688980957
transform 1 0 51980 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_559
timestamp 1688980957
transform 1 0 52532 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_561
timestamp 1688980957
transform 1 0 52716 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_573
timestamp 1688980957
transform 1 0 53820 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_581
timestamp 1688980957
transform 1 0 54556 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_587
timestamp 1688980957
transform 1 0 55108 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_592
timestamp 1688980957
transform 1 0 55568 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_604
timestamp 1688980957
transform 1 0 56672 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_614
timestamp 1688980957
transform 1 0 57592 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_35
timestamp 1688980957
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_43
timestamp 1688980957
transform 1 0 5060 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_51
timestamp 1688980957
transform 1 0 5796 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_97
timestamp 1688980957
transform 1 0 10028 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_117
timestamp 1688980957
transform 1 0 11868 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1688980957
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 1688980957
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 1688980957
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 1688980957
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 1688980957
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 1688980957
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 1688980957
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 1688980957
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 1688980957
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 1688980957
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 1688980957
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 1688980957
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 1688980957
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 1688980957
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 1688980957
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 1688980957
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 1688980957
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 1688980957
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_377
timestamp 1688980957
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 1688980957
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_401
timestamp 1688980957
transform 1 0 37996 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_413
timestamp 1688980957
transform 1 0 39100 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_419
timestamp 1688980957
transform 1 0 39652 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_421
timestamp 1688980957
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_433
timestamp 1688980957
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_445
timestamp 1688980957
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_457
timestamp 1688980957
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_469
timestamp 1688980957
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_475
timestamp 1688980957
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_477
timestamp 1688980957
transform 1 0 44988 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_500
timestamp 1688980957
transform 1 0 47104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_530
timestamp 1688980957
transform 1 0 49864 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_542
timestamp 1688980957
transform 1 0 50968 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_546
timestamp 1688980957
transform 1 0 51336 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_556
timestamp 1688980957
transform 1 0 52256 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_564
timestamp 1688980957
transform 1 0 52992 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_574
timestamp 1688980957
transform 1 0 53912 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_579
timestamp 1688980957
transform 1 0 54372 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_624
timestamp 1688980957
transform 1 0 58512 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_25
timestamp 1688980957
transform 1 0 3404 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_32
timestamp 1688980957
transform 1 0 4048 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_50
timestamp 1688980957
transform 1 0 5704 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_64
timestamp 1688980957
transform 1 0 6992 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_72
timestamp 1688980957
transform 1 0 7728 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 1688980957
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_93
timestamp 1688980957
transform 1 0 9660 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_97
timestamp 1688980957
transform 1 0 10028 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_109
timestamp 1688980957
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_117
timestamp 1688980957
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_129
timestamp 1688980957
transform 1 0 12972 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_133
timestamp 1688980957
transform 1 0 13340 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_145
timestamp 1688980957
transform 1 0 14444 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_157
timestamp 1688980957
transform 1 0 15548 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1688980957
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_181
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_185
timestamp 1688980957
transform 1 0 18124 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_206
timestamp 1688980957
transform 1 0 20056 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_210
timestamp 1688980957
transform 1 0 20424 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_222
timestamp 1688980957
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 1688980957
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 1688980957
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1688980957
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 1688980957
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 1688980957
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 1688980957
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 1688980957
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 1688980957
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 1688980957
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_361
timestamp 1688980957
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_373
timestamp 1688980957
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 1688980957
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 1688980957
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_405
timestamp 1688980957
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_417
timestamp 1688980957
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_429
timestamp 1688980957
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_441
timestamp 1688980957
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_447
timestamp 1688980957
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_449
timestamp 1688980957
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_461
timestamp 1688980957
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_473
timestamp 1688980957
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_485
timestamp 1688980957
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_497
timestamp 1688980957
transform 1 0 46828 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_520
timestamp 1688980957
transform 1 0 48944 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_524
timestamp 1688980957
transform 1 0 49312 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_527
timestamp 1688980957
transform 1 0 49588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_539
timestamp 1688980957
transform 1 0 50692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_554
timestamp 1688980957
transform 1 0 52072 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_567
timestamp 1688980957
transform 1 0 53268 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_579
timestamp 1688980957
transform 1 0 54372 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_602
timestamp 1688980957
transform 1 0 56488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_37
timestamp 1688980957
transform 1 0 4508 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_43
timestamp 1688980957
transform 1 0 5060 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_55
timestamp 1688980957
transform 1 0 6164 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_62
timestamp 1688980957
transform 1 0 6808 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_74
timestamp 1688980957
transform 1 0 7912 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_91
timestamp 1688980957
transform 1 0 9476 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_96
timestamp 1688980957
transform 1 0 9936 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_138
timestamp 1688980957
transform 1 0 13800 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_145
timestamp 1688980957
transform 1 0 14444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_157
timestamp 1688980957
transform 1 0 15548 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_169
timestamp 1688980957
transform 1 0 16652 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_181
timestamp 1688980957
transform 1 0 17756 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_193
timestamp 1688980957
transform 1 0 18860 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 1688980957
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 1688980957
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 1688980957
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 1688980957
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 1688980957
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 1688980957
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 1688980957
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 1688980957
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 1688980957
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 1688980957
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 1688980957
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 1688980957
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 1688980957
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 1688980957
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 1688980957
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_389
timestamp 1688980957
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_401
timestamp 1688980957
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_413
timestamp 1688980957
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_419
timestamp 1688980957
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_421
timestamp 1688980957
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_433
timestamp 1688980957
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_445
timestamp 1688980957
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_457
timestamp 1688980957
transform 1 0 43148 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_465
timestamp 1688980957
transform 1 0 43884 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_469
timestamp 1688980957
transform 1 0 44252 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_475
timestamp 1688980957
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_480
timestamp 1688980957
transform 1 0 45264 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_484
timestamp 1688980957
transform 1 0 45632 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_488
timestamp 1688980957
transform 1 0 46000 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_506
timestamp 1688980957
transform 1 0 47656 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_530
timestamp 1688980957
transform 1 0 49864 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_539
timestamp 1688980957
transform 1 0 50692 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_550
timestamp 1688980957
transform 1 0 51704 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_562
timestamp 1688980957
transform 1 0 52808 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_574
timestamp 1688980957
transform 1 0 53912 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_582
timestamp 1688980957
transform 1 0 54648 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_587
timestamp 1688980957
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_617
timestamp 1688980957
transform 1 0 57868 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_624
timestamp 1688980957
transform 1 0 58512 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_19
timestamp 1688980957
transform 1 0 2852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_30
timestamp 1688980957
transform 1 0 3864 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_35
timestamp 1688980957
transform 1 0 4324 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_41
timestamp 1688980957
transform 1 0 4876 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_49
timestamp 1688980957
transform 1 0 5612 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_61
timestamp 1688980957
transform 1 0 6716 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_65
timestamp 1688980957
transform 1 0 7084 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_73
timestamp 1688980957
transform 1 0 7820 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_78
timestamp 1688980957
transform 1 0 8280 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_90
timestamp 1688980957
transform 1 0 9384 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_96
timestamp 1688980957
transform 1 0 9936 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 1688980957
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 1688980957
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_121
timestamp 1688980957
transform 1 0 12236 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 1688980957
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 1688980957
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 1688980957
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 1688980957
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 1688980957
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 1688980957
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 1688980957
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 1688980957
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 1688980957
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 1688980957
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 1688980957
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 1688980957
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 1688980957
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 1688980957
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 1688980957
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_361
timestamp 1688980957
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_373
timestamp 1688980957
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_385
timestamp 1688980957
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 1688980957
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_405
timestamp 1688980957
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_417
timestamp 1688980957
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_429
timestamp 1688980957
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_441
timestamp 1688980957
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_447
timestamp 1688980957
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_449
timestamp 1688980957
transform 1 0 42412 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_457
timestamp 1688980957
transform 1 0 43148 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_466
timestamp 1688980957
transform 1 0 43976 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_493
timestamp 1688980957
transform 1 0 46460 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_497
timestamp 1688980957
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_503
timestamp 1688980957
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_505
timestamp 1688980957
transform 1 0 47564 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_536
timestamp 1688980957
transform 1 0 50416 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_543
timestamp 1688980957
transform 1 0 51060 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_547
timestamp 1688980957
transform 1 0 51428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_559
timestamp 1688980957
transform 1 0 52532 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_604
timestamp 1688980957
transform 1 0 56672 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_614
timestamp 1688980957
transform 1 0 57592 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_11
timestamp 1688980957
transform 1 0 2116 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_16
timestamp 1688980957
transform 1 0 2576 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_91
timestamp 1688980957
transform 1 0 9476 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_94
timestamp 1688980957
transform 1 0 9752 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_102
timestamp 1688980957
transform 1 0 10488 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_110
timestamp 1688980957
transform 1 0 11224 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_117
timestamp 1688980957
transform 1 0 11868 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 1688980957
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 1688980957
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 1688980957
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 1688980957
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 1688980957
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 1688980957
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 1688980957
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 1688980957
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 1688980957
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 1688980957
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 1688980957
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 1688980957
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 1688980957
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 1688980957
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 1688980957
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 1688980957
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 1688980957
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 1688980957
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_389
timestamp 1688980957
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_401
timestamp 1688980957
transform 1 0 37996 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_413
timestamp 1688980957
transform 1 0 39100 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_419
timestamp 1688980957
transform 1 0 39652 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_421
timestamp 1688980957
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_456
timestamp 1688980957
transform 1 0 43056 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_460
timestamp 1688980957
transform 1 0 43424 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_472
timestamp 1688980957
transform 1 0 44528 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_493
timestamp 1688980957
transform 1 0 46460 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_499
timestamp 1688980957
transform 1 0 47012 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_506
timestamp 1688980957
transform 1 0 47656 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_512
timestamp 1688980957
transform 1 0 48208 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_519
timestamp 1688980957
transform 1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_525
timestamp 1688980957
transform 1 0 49404 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_529
timestamp 1688980957
transform 1 0 49772 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_533
timestamp 1688980957
transform 1 0 50140 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_541
timestamp 1688980957
transform 1 0 50876 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_556
timestamp 1688980957
transform 1 0 52256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_569
timestamp 1688980957
transform 1 0 53452 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_593
timestamp 1688980957
transform 1 0 55660 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_610
timestamp 1688980957
transform 1 0 57224 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_34
timestamp 1688980957
transform 1 0 4232 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_40
timestamp 1688980957
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_52
timestamp 1688980957
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_73
timestamp 1688980957
transform 1 0 7820 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_80
timestamp 1688980957
transform 1 0 8464 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_84
timestamp 1688980957
transform 1 0 8832 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_119
timestamp 1688980957
transform 1 0 12052 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_130
timestamp 1688980957
transform 1 0 13064 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_142
timestamp 1688980957
transform 1 0 14168 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_154
timestamp 1688980957
transform 1 0 15272 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_166
timestamp 1688980957
transform 1 0 16376 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 1688980957
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1688980957
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1688980957
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 1688980957
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 1688980957
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 1688980957
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 1688980957
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 1688980957
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 1688980957
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 1688980957
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 1688980957
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 1688980957
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 1688980957
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 1688980957
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 1688980957
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_373
timestamp 1688980957
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 1688980957
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 1688980957
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_405
timestamp 1688980957
transform 1 0 38364 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_413
timestamp 1688980957
transform 1 0 39100 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_417
timestamp 1688980957
transform 1 0 39468 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_421
timestamp 1688980957
transform 1 0 39836 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_425
timestamp 1688980957
transform 1 0 40204 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_429
timestamp 1688980957
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_441
timestamp 1688980957
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_447
timestamp 1688980957
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_457
timestamp 1688980957
transform 1 0 43148 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_469
timestamp 1688980957
transform 1 0 44252 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_481
timestamp 1688980957
transform 1 0 45356 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_511
timestamp 1688980957
transform 1 0 48116 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_541
timestamp 1688980957
transform 1 0 50876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_553
timestamp 1688980957
transform 1 0 51980 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_559
timestamp 1688980957
transform 1 0 52532 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_561
timestamp 1688980957
transform 1 0 52716 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_572
timestamp 1688980957
transform 1 0 53728 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_584
timestamp 1688980957
transform 1 0 54832 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_590
timestamp 1688980957
transform 1 0 55384 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_602
timestamp 1688980957
transform 1 0 56488 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_613
timestamp 1688980957
transform 1 0 57500 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_617
timestamp 1688980957
transform 1 0 57868 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_32
timestamp 1688980957
transform 1 0 4048 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_59
timestamp 1688980957
transform 1 0 6532 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_64
timestamp 1688980957
transform 1 0 6992 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_69
timestamp 1688980957
transform 1 0 7452 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_73
timestamp 1688980957
transform 1 0 7820 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_79
timestamp 1688980957
transform 1 0 8372 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_93
timestamp 1688980957
transform 1 0 9660 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_99
timestamp 1688980957
transform 1 0 10212 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_111
timestamp 1688980957
transform 1 0 11316 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_119
timestamp 1688980957
transform 1 0 12052 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_124
timestamp 1688980957
transform 1 0 12512 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_129
timestamp 1688980957
transform 1 0 12972 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_137
timestamp 1688980957
transform 1 0 13708 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 1688980957
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 1688980957
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 1688980957
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 1688980957
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 1688980957
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 1688980957
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 1688980957
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 1688980957
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 1688980957
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 1688980957
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 1688980957
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 1688980957
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 1688980957
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 1688980957
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 1688980957
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 1688980957
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_377
timestamp 1688980957
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_389
timestamp 1688980957
transform 1 0 36892 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_415
timestamp 1688980957
transform 1 0 39284 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_444
timestamp 1688980957
transform 1 0 41952 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_449
timestamp 1688980957
transform 1 0 42412 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_453
timestamp 1688980957
transform 1 0 42780 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_465
timestamp 1688980957
transform 1 0 43884 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_473
timestamp 1688980957
transform 1 0 44620 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_500
timestamp 1688980957
transform 1 0 47104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_504
timestamp 1688980957
transform 1 0 47472 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_511
timestamp 1688980957
transform 1 0 48116 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_531
timestamp 1688980957
transform 1 0 49956 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_564
timestamp 1688980957
transform 1 0 52992 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_568
timestamp 1688980957
transform 1 0 53360 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_572
timestamp 1688980957
transform 1 0 53728 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_584
timestamp 1688980957
transform 1 0 54832 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_595
timestamp 1688980957
transform 1 0 55844 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_599
timestamp 1688980957
transform 1 0 56212 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_617
timestamp 1688980957
transform 1 0 57868 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_624
timestamp 1688980957
transform 1 0 58512 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_25
timestamp 1688980957
transform 1 0 3404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_92
timestamp 1688980957
transform 1 0 9568 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_104
timestamp 1688980957
transform 1 0 10672 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_108
timestamp 1688980957
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_117
timestamp 1688980957
transform 1 0 11868 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_122
timestamp 1688980957
transform 1 0 12328 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_145
timestamp 1688980957
transform 1 0 14444 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_157
timestamp 1688980957
transform 1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_165
timestamp 1688980957
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 1688980957
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 1688980957
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 1688980957
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 1688980957
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 1688980957
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 1688980957
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 1688980957
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 1688980957
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 1688980957
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1688980957
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1688980957
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 1688980957
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_361
timestamp 1688980957
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_373
timestamp 1688980957
transform 1 0 35420 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_391
timestamp 1688980957
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_393
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_409
timestamp 1688980957
transform 1 0 38732 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_421
timestamp 1688980957
transform 1 0 39836 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_429
timestamp 1688980957
transform 1 0 40572 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_438
timestamp 1688980957
transform 1 0 41400 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_447
timestamp 1688980957
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_472
timestamp 1688980957
transform 1 0 44528 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_484
timestamp 1688980957
transform 1 0 45632 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_495
timestamp 1688980957
transform 1 0 46644 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_503
timestamp 1688980957
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_505
timestamp 1688980957
transform 1 0 47564 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_512
timestamp 1688980957
transform 1 0 48208 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_520
timestamp 1688980957
transform 1 0 48944 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_540
timestamp 1688980957
transform 1 0 50784 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_552
timestamp 1688980957
transform 1 0 51888 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_564
timestamp 1688980957
transform 1 0 52992 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_572
timestamp 1688980957
transform 1 0 53728 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_588
timestamp 1688980957
transform 1 0 55200 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_596
timestamp 1688980957
transform 1 0 55936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_615
timestamp 1688980957
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_37
timestamp 1688980957
transform 1 0 4508 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_42
timestamp 1688980957
transform 1 0 4968 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_54
timestamp 1688980957
transform 1 0 6072 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_60
timestamp 1688980957
transform 1 0 6624 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_72
timestamp 1688980957
transform 1 0 7728 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_76
timestamp 1688980957
transform 1 0 8096 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_81
timestamp 1688980957
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_93
timestamp 1688980957
transform 1 0 9660 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_127
timestamp 1688980957
transform 1 0 12788 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_145
timestamp 1688980957
transform 1 0 14444 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_157
timestamp 1688980957
transform 1 0 15548 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_169
timestamp 1688980957
transform 1 0 16652 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_181
timestamp 1688980957
transform 1 0 17756 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_193
timestamp 1688980957
transform 1 0 18860 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 1688980957
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 1688980957
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 1688980957
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 1688980957
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 1688980957
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 1688980957
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1688980957
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 1688980957
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 1688980957
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 1688980957
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 1688980957
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 1688980957
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 1688980957
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_424
timestamp 1688980957
transform 1 0 40112 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_436
timestamp 1688980957
transform 1 0 41216 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_457
timestamp 1688980957
transform 1 0 43148 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_461
timestamp 1688980957
transform 1 0 43516 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_465
timestamp 1688980957
transform 1 0 43884 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_474
timestamp 1688980957
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_485
timestamp 1688980957
transform 1 0 45724 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_493
timestamp 1688980957
transform 1 0 46460 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_504
timestamp 1688980957
transform 1 0 47472 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_508
timestamp 1688980957
transform 1 0 47840 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_512
timestamp 1688980957
transform 1 0 48208 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_526
timestamp 1688980957
transform 1 0 49496 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_530
timestamp 1688980957
transform 1 0 49864 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_533
timestamp 1688980957
transform 1 0 50140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_537
timestamp 1688980957
transform 1 0 50508 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_541
timestamp 1688980957
transform 1 0 50876 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_551
timestamp 1688980957
transform 1 0 51796 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_559
timestamp 1688980957
transform 1 0 52532 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_565
timestamp 1688980957
transform 1 0 53084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_577
timestamp 1688980957
transform 1 0 54188 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_581
timestamp 1688980957
transform 1 0 54556 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_585
timestamp 1688980957
transform 1 0 54924 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_600
timestamp 1688980957
transform 1 0 56304 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_609
timestamp 1688980957
transform 1 0 57132 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_623
timestamp 1688980957
transform 1 0 58420 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_19
timestamp 1688980957
transform 1 0 2852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_30
timestamp 1688980957
transform 1 0 3864 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_34
timestamp 1688980957
transform 1 0 4232 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_46
timestamp 1688980957
transform 1 0 5336 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_54
timestamp 1688980957
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 1688980957
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_97
timestamp 1688980957
transform 1 0 10028 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_100
timestamp 1688980957
transform 1 0 10304 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_122
timestamp 1688980957
transform 1 0 12328 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_127
timestamp 1688980957
transform 1 0 12788 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_147
timestamp 1688980957
transform 1 0 14628 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_159
timestamp 1688980957
transform 1 0 15732 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 1688980957
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 1688980957
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 1688980957
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 1688980957
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 1688980957
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 1688980957
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 1688980957
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 1688980957
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 1688980957
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 1688980957
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 1688980957
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 1688980957
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_385
timestamp 1688980957
transform 1 0 36524 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_389
timestamp 1688980957
transform 1 0 36892 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_399
timestamp 1688980957
transform 1 0 37812 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_413
timestamp 1688980957
transform 1 0 39100 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_419
timestamp 1688980957
transform 1 0 39652 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_423
timestamp 1688980957
transform 1 0 40020 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_433
timestamp 1688980957
transform 1 0 40940 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_438
timestamp 1688980957
transform 1 0 41400 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_442
timestamp 1688980957
transform 1 0 41768 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_446
timestamp 1688980957
transform 1 0 42136 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_449
timestamp 1688980957
transform 1 0 42412 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_474
timestamp 1688980957
transform 1 0 44712 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_483
timestamp 1688980957
transform 1 0 45540 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_505
timestamp 1688980957
transform 1 0 47564 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_537
timestamp 1688980957
transform 1 0 50508 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_555
timestamp 1688980957
transform 1 0 52164 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_559
timestamp 1688980957
transform 1 0 52532 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_570
timestamp 1688980957
transform 1 0 53544 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_574
timestamp 1688980957
transform 1 0 53912 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_602
timestamp 1688980957
transform 1 0 56488 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_610
timestamp 1688980957
transform 1 0 57224 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_623
timestamp 1688980957
transform 1 0 58420 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_11
timestamp 1688980957
transform 1 0 2116 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_17
timestamp 1688980957
transform 1 0 2668 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_26
timestamp 1688980957
transform 1 0 3496 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_35
timestamp 1688980957
transform 1 0 4324 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_46
timestamp 1688980957
transform 1 0 5336 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_71
timestamp 1688980957
transform 1 0 7636 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_77
timestamp 1688980957
transform 1 0 8188 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_91
timestamp 1688980957
transform 1 0 9476 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_101
timestamp 1688980957
transform 1 0 10396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_113
timestamp 1688980957
transform 1 0 11500 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_121
timestamp 1688980957
transform 1 0 12236 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_125
timestamp 1688980957
transform 1 0 12604 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_136
timestamp 1688980957
transform 1 0 13616 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 1688980957
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 1688980957
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 1688980957
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 1688980957
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 1688980957
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 1688980957
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 1688980957
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 1688980957
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 1688980957
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 1688980957
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 1688980957
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 1688980957
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 1688980957
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 1688980957
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_377
timestamp 1688980957
transform 1 0 35788 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_385
timestamp 1688980957
transform 1 0 36524 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_403
timestamp 1688980957
transform 1 0 38180 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_412
timestamp 1688980957
transform 1 0 39008 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_416
timestamp 1688980957
transform 1 0 39376 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_424
timestamp 1688980957
transform 1 0 40112 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_428
timestamp 1688980957
transform 1 0 40480 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_449
timestamp 1688980957
transform 1 0 42412 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_470
timestamp 1688980957
transform 1 0 44344 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_474
timestamp 1688980957
transform 1 0 44712 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_503
timestamp 1688980957
transform 1 0 47380 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_512
timestamp 1688980957
transform 1 0 48208 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_525
timestamp 1688980957
transform 1 0 49404 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_531
timestamp 1688980957
transform 1 0 49956 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_533
timestamp 1688980957
transform 1 0 50140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_549
timestamp 1688980957
transform 1 0 51612 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_561
timestamp 1688980957
transform 1 0 52716 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_575
timestamp 1688980957
transform 1 0 54004 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_580
timestamp 1688980957
transform 1 0 54464 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_584
timestamp 1688980957
transform 1 0 54832 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_597
timestamp 1688980957
transform 1 0 56028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_613
timestamp 1688980957
transform 1 0 57500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_623
timestamp 1688980957
transform 1 0 58420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_31
timestamp 1688980957
transform 1 0 3956 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_48
timestamp 1688980957
transform 1 0 5520 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_65
timestamp 1688980957
transform 1 0 7084 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_70
timestamp 1688980957
transform 1 0 7544 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_84
timestamp 1688980957
transform 1 0 8832 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_92
timestamp 1688980957
transform 1 0 9568 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_98
timestamp 1688980957
transform 1 0 10120 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_106
timestamp 1688980957
transform 1 0 10856 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 1688980957
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 1688980957
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 1688980957
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 1688980957
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 1688980957
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 1688980957
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_311
timestamp 1688980957
transform 1 0 29716 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_332
timestamp 1688980957
transform 1 0 31648 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 1688980957
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 1688980957
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_390
timestamp 1688980957
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_396
timestamp 1688980957
transform 1 0 37536 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_401
timestamp 1688980957
transform 1 0 37996 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_405
timestamp 1688980957
transform 1 0 38364 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_411
timestamp 1688980957
transform 1 0 38916 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_415
timestamp 1688980957
transform 1 0 39284 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_419
timestamp 1688980957
transform 1 0 39652 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_423
timestamp 1688980957
transform 1 0 40020 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_435
timestamp 1688980957
transform 1 0 41124 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_438
timestamp 1688980957
transform 1 0 41400 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_443
timestamp 1688980957
transform 1 0 41860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_447
timestamp 1688980957
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_449
timestamp 1688980957
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_461
timestamp 1688980957
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_473
timestamp 1688980957
transform 1 0 44620 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_479
timestamp 1688980957
transform 1 0 45172 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_483
timestamp 1688980957
transform 1 0 45540 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_493
timestamp 1688980957
transform 1 0 46460 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_499
timestamp 1688980957
transform 1 0 47012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_503
timestamp 1688980957
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_505
timestamp 1688980957
transform 1 0 47564 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_513
timestamp 1688980957
transform 1 0 48300 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_517
timestamp 1688980957
transform 1 0 48668 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_521
timestamp 1688980957
transform 1 0 49036 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_542
timestamp 1688980957
transform 1 0 50968 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_559
timestamp 1688980957
transform 1 0 52532 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_572
timestamp 1688980957
transform 1 0 53728 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_580
timestamp 1688980957
transform 1 0 54464 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_584
timestamp 1688980957
transform 1 0 54832 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_588
timestamp 1688980957
transform 1 0 55200 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_600
timestamp 1688980957
transform 1 0 56304 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_606
timestamp 1688980957
transform 1 0 56856 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_611
timestamp 1688980957
transform 1 0 57316 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_615
timestamp 1688980957
transform 1 0 57684 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_623
timestamp 1688980957
transform 1 0 58420 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_32
timestamp 1688980957
transform 1 0 4048 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_53
timestamp 1688980957
transform 1 0 5980 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_58
timestamp 1688980957
transform 1 0 6440 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_63
timestamp 1688980957
transform 1 0 6900 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_75
timestamp 1688980957
transform 1 0 8004 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_79
timestamp 1688980957
transform 1 0 8372 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 1688980957
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_93
timestamp 1688980957
transform 1 0 9660 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_99
timestamp 1688980957
transform 1 0 10212 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_111
timestamp 1688980957
transform 1 0 11316 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_119
timestamp 1688980957
transform 1 0 12052 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_145
timestamp 1688980957
transform 1 0 14444 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_157
timestamp 1688980957
transform 1 0 15548 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_169
timestamp 1688980957
transform 1 0 16652 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_181
timestamp 1688980957
transform 1 0 17756 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_193
timestamp 1688980957
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 1688980957
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 1688980957
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 1688980957
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 1688980957
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 1688980957
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 1688980957
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 1688980957
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 1688980957
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 1688980957
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 1688980957
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 1688980957
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 1688980957
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_365
timestamp 1688980957
transform 1 0 34684 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_414
timestamp 1688980957
transform 1 0 39192 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_418
timestamp 1688980957
transform 1 0 39560 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_421
timestamp 1688980957
transform 1 0 39836 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_425
timestamp 1688980957
transform 1 0 40204 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_430
timestamp 1688980957
transform 1 0 40664 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_442
timestamp 1688980957
transform 1 0 41768 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_446
timestamp 1688980957
transform 1 0 42136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_450
timestamp 1688980957
transform 1 0 42504 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_454
timestamp 1688980957
transform 1 0 42872 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_459
timestamp 1688980957
transform 1 0 43332 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_471
timestamp 1688980957
transform 1 0 44436 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_483
timestamp 1688980957
transform 1 0 45540 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_495
timestamp 1688980957
transform 1 0 46644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_510
timestamp 1688980957
transform 1 0 48024 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_553
timestamp 1688980957
transform 1 0 51980 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_583
timestamp 1688980957
transform 1 0 54740 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_624
timestamp 1688980957
transform 1 0 58512 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_9
timestamp 1688980957
transform 1 0 1932 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_22
timestamp 1688980957
transform 1 0 3128 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_34
timestamp 1688980957
transform 1 0 4232 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_43
timestamp 1688980957
transform 1 0 5060 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_61
timestamp 1688980957
transform 1 0 6716 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_86
timestamp 1688980957
transform 1 0 9016 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_94
timestamp 1688980957
transform 1 0 9752 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_105
timestamp 1688980957
transform 1 0 10764 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_120
timestamp 1688980957
transform 1 0 12144 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_125
timestamp 1688980957
transform 1 0 12604 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_129
timestamp 1688980957
transform 1 0 12972 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_141
timestamp 1688980957
transform 1 0 14076 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_153
timestamp 1688980957
transform 1 0 15180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_165
timestamp 1688980957
transform 1 0 16284 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 1688980957
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 1688980957
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 1688980957
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 1688980957
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 1688980957
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 1688980957
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 1688980957
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 1688980957
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 1688980957
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 1688980957
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 1688980957
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 1688980957
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 1688980957
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 1688980957
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_373
timestamp 1688980957
transform 1 0 35420 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_381
timestamp 1688980957
transform 1 0 36156 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_390
timestamp 1688980957
transform 1 0 36984 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_397
timestamp 1688980957
transform 1 0 37628 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_403
timestamp 1688980957
transform 1 0 38180 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_412
timestamp 1688980957
transform 1 0 39008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_418
timestamp 1688980957
transform 1 0 39560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_446
timestamp 1688980957
transform 1 0 42136 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_452
timestamp 1688980957
transform 1 0 42688 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_468
timestamp 1688980957
transform 1 0 44160 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_478
timestamp 1688980957
transform 1 0 45080 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_495
timestamp 1688980957
transform 1 0 46644 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_499
timestamp 1688980957
transform 1 0 47012 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_503
timestamp 1688980957
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_505
timestamp 1688980957
transform 1 0 47564 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_515
timestamp 1688980957
transform 1 0 48484 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_519
timestamp 1688980957
transform 1 0 48852 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_523
timestamp 1688980957
transform 1 0 49220 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_551
timestamp 1688980957
transform 1 0 51796 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_559
timestamp 1688980957
transform 1 0 52532 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_561
timestamp 1688980957
transform 1 0 52716 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_572
timestamp 1688980957
transform 1 0 53728 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_582
timestamp 1688980957
transform 1 0 54648 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_598
timestamp 1688980957
transform 1 0 56120 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_615
timestamp 1688980957
transform 1 0 57684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_26
timestamp 1688980957
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_51
timestamp 1688980957
transform 1 0 5796 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_55
timestamp 1688980957
transform 1 0 6164 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_61
timestamp 1688980957
transform 1 0 6716 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_72
timestamp 1688980957
transform 1 0 7728 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_76
timestamp 1688980957
transform 1 0 8096 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_89
timestamp 1688980957
transform 1 0 9292 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_105
timestamp 1688980957
transform 1 0 10764 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_128
timestamp 1688980957
transform 1 0 12880 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_132
timestamp 1688980957
transform 1 0 13248 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_136
timestamp 1688980957
transform 1 0 13616 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_157
timestamp 1688980957
transform 1 0 15548 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_169
timestamp 1688980957
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_181
timestamp 1688980957
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_193
timestamp 1688980957
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 1688980957
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 1688980957
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_266
timestamp 1688980957
transform 1 0 25576 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_270
timestamp 1688980957
transform 1 0 25944 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_282
timestamp 1688980957
transform 1 0 27048 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_294
timestamp 1688980957
transform 1 0 28152 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_306
timestamp 1688980957
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 1688980957
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 1688980957
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 1688980957
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_357
timestamp 1688980957
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 1688980957
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1688980957
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_389
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_397
timestamp 1688980957
transform 1 0 37628 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_404
timestamp 1688980957
transform 1 0 38272 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_412
timestamp 1688980957
transform 1 0 39008 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_416
timestamp 1688980957
transform 1 0 39376 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_428
timestamp 1688980957
transform 1 0 40480 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_440
timestamp 1688980957
transform 1 0 41584 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_448
timestamp 1688980957
transform 1 0 42320 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_456
timestamp 1688980957
transform 1 0 43056 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_463
timestamp 1688980957
transform 1 0 43700 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_467
timestamp 1688980957
transform 1 0 44068 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_491
timestamp 1688980957
transform 1 0 46276 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_495
timestamp 1688980957
transform 1 0 46644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_503
timestamp 1688980957
transform 1 0 47380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_507
timestamp 1688980957
transform 1 0 47748 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_518
timestamp 1688980957
transform 1 0 48760 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_522
timestamp 1688980957
transform 1 0 49128 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_526
timestamp 1688980957
transform 1 0 49496 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_536
timestamp 1688980957
transform 1 0 50416 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_540
timestamp 1688980957
transform 1 0 50784 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_560
timestamp 1688980957
transform 1 0 52624 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_564
timestamp 1688980957
transform 1 0 52992 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_568
timestamp 1688980957
transform 1 0 53360 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_587
timestamp 1688980957
transform 1 0 55108 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_592
timestamp 1688980957
transform 1 0 55568 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_615
timestamp 1688980957
transform 1 0 57684 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_33
timestamp 1688980957
transform 1 0 4140 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_39
timestamp 1688980957
transform 1 0 4692 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_43
timestamp 1688980957
transform 1 0 5060 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_47
timestamp 1688980957
transform 1 0 5428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_63
timestamp 1688980957
transform 1 0 6900 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_93
timestamp 1688980957
transform 1 0 9660 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_101
timestamp 1688980957
transform 1 0 10396 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_107
timestamp 1688980957
transform 1 0 10948 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 1688980957
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_131
timestamp 1688980957
transform 1 0 13156 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_135
timestamp 1688980957
transform 1 0 13524 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_147
timestamp 1688980957
transform 1 0 14628 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_159
timestamp 1688980957
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 1688980957
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 1688980957
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 1688980957
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 1688980957
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 1688980957
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 1688980957
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 1688980957
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 1688980957
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_361
timestamp 1688980957
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_373
timestamp 1688980957
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_385
timestamp 1688980957
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 1688980957
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_393
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_401
timestamp 1688980957
transform 1 0 37996 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_428
timestamp 1688980957
transform 1 0 40480 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_433
timestamp 1688980957
transform 1 0 40940 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_438
timestamp 1688980957
transform 1 0 41400 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_442
timestamp 1688980957
transform 1 0 41768 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_449
timestamp 1688980957
transform 1 0 42412 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_457
timestamp 1688980957
transform 1 0 43148 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_464
timestamp 1688980957
transform 1 0 43792 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_468
timestamp 1688980957
transform 1 0 44160 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_472
timestamp 1688980957
transform 1 0 44528 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_530
timestamp 1688980957
transform 1 0 49864 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_534
timestamp 1688980957
transform 1 0 50232 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_546
timestamp 1688980957
transform 1 0 51336 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_597
timestamp 1688980957
transform 1 0 56028 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_614
timestamp 1688980957
transform 1 0 57592 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_26
timestamp 1688980957
transform 1 0 3496 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_36
timestamp 1688980957
transform 1 0 4416 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_41
timestamp 1688980957
transform 1 0 4876 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_45
timestamp 1688980957
transform 1 0 5244 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_75
timestamp 1688980957
transform 1 0 8004 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_93
timestamp 1688980957
transform 1 0 9660 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_98
timestamp 1688980957
transform 1 0 10120 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_104
timestamp 1688980957
transform 1 0 10672 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_115
timestamp 1688980957
transform 1 0 11684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_127
timestamp 1688980957
transform 1 0 12788 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_131
timestamp 1688980957
transform 1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 1688980957
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 1688980957
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 1688980957
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 1688980957
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 1688980957
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 1688980957
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 1688980957
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 1688980957
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 1688980957
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 1688980957
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 1688980957
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 1688980957
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 1688980957
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 1688980957
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 1688980957
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 1688980957
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 1688980957
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_377
timestamp 1688980957
transform 1 0 35788 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_410
timestamp 1688980957
transform 1 0 38824 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_414
timestamp 1688980957
transform 1 0 39192 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_418
timestamp 1688980957
transform 1 0 39560 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_421
timestamp 1688980957
transform 1 0 39836 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_429
timestamp 1688980957
transform 1 0 40572 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_451
timestamp 1688980957
transform 1 0 42596 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_477
timestamp 1688980957
transform 1 0 44988 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_504
timestamp 1688980957
transform 1 0 47472 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_508
timestamp 1688980957
transform 1 0 47840 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_539
timestamp 1688980957
transform 1 0 50692 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_547
timestamp 1688980957
transform 1 0 51428 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_558
timestamp 1688980957
transform 1 0 52440 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_569
timestamp 1688980957
transform 1 0 53452 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_581
timestamp 1688980957
transform 1 0 54556 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_587
timestamp 1688980957
transform 1 0 55108 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_589
timestamp 1688980957
transform 1 0 55292 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_601
timestamp 1688980957
transform 1 0 56396 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_607
timestamp 1688980957
transform 1 0 56948 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_610
timestamp 1688980957
transform 1 0 57224 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_616
timestamp 1688980957
transform 1 0 57776 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_623
timestamp 1688980957
transform 1 0 58420 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_31
timestamp 1688980957
transform 1 0 3956 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_52
timestamp 1688980957
transform 1 0 5888 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_62
timestamp 1688980957
transform 1 0 6808 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_74
timestamp 1688980957
transform 1 0 7912 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_82
timestamp 1688980957
transform 1 0 8648 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_110
timestamp 1688980957
transform 1 0 11224 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_130
timestamp 1688980957
transform 1 0 13064 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_134
timestamp 1688980957
transform 1 0 13432 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_146
timestamp 1688980957
transform 1 0 14536 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_158
timestamp 1688980957
transform 1 0 15640 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_166
timestamp 1688980957
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 1688980957
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 1688980957
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 1688980957
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 1688980957
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 1688980957
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 1688980957
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 1688980957
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 1688980957
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 1688980957
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 1688980957
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 1688980957
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 1688980957
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 1688980957
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_361
timestamp 1688980957
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_373
timestamp 1688980957
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_385
timestamp 1688980957
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 1688980957
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_393
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_420
timestamp 1688980957
transform 1 0 39744 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_457
timestamp 1688980957
transform 1 0 43148 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_462
timestamp 1688980957
transform 1 0 43608 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_515
timestamp 1688980957
transform 1 0 48484 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_532
timestamp 1688980957
transform 1 0 50048 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_540
timestamp 1688980957
transform 1 0 50784 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_548
timestamp 1688980957
transform 1 0 51520 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_552
timestamp 1688980957
transform 1 0 51888 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_556
timestamp 1688980957
transform 1 0 52256 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_561
timestamp 1688980957
transform 1 0 52716 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_565
timestamp 1688980957
transform 1 0 53084 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_573
timestamp 1688980957
transform 1 0 53820 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_581
timestamp 1688980957
transform 1 0 54556 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_603
timestamp 1688980957
transform 1 0 56580 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_613
timestamp 1688980957
transform 1 0 57500 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_617
timestamp 1688980957
transform 1 0 57868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_623
timestamp 1688980957
transform 1 0 58420 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_19
timestamp 1688980957
transform 1 0 2852 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_40
timestamp 1688980957
transform 1 0 4784 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_52
timestamp 1688980957
transform 1 0 5888 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_55
timestamp 1688980957
transform 1 0 6164 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_66
timestamp 1688980957
transform 1 0 7176 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_74
timestamp 1688980957
transform 1 0 7912 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_91
timestamp 1688980957
transform 1 0 9476 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_95
timestamp 1688980957
transform 1 0 9844 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_106
timestamp 1688980957
transform 1 0 10856 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_114
timestamp 1688980957
transform 1 0 11592 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_125
timestamp 1688980957
transform 1 0 12604 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_137
timestamp 1688980957
transform 1 0 13708 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_157
timestamp 1688980957
transform 1 0 15548 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_161
timestamp 1688980957
transform 1 0 15916 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_173
timestamp 1688980957
transform 1 0 17020 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_185
timestamp 1688980957
transform 1 0 18124 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_193
timestamp 1688980957
transform 1 0 18860 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 1688980957
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 1688980957
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 1688980957
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 1688980957
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 1688980957
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 1688980957
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 1688980957
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 1688980957
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 1688980957
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 1688980957
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 1688980957
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 1688980957
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 1688980957
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_377
timestamp 1688980957
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_389
timestamp 1688980957
transform 1 0 36892 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_414
timestamp 1688980957
transform 1 0 39192 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_421
timestamp 1688980957
transform 1 0 39836 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_425
timestamp 1688980957
transform 1 0 40204 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_437
timestamp 1688980957
transform 1 0 41308 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_450
timestamp 1688980957
transform 1 0 42504 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_460
timestamp 1688980957
transform 1 0 43424 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_468
timestamp 1688980957
transform 1 0 44160 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_500
timestamp 1688980957
transform 1 0 47104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_524
timestamp 1688980957
transform 1 0 49312 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_559
timestamp 1688980957
transform 1 0 52532 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_563
timestamp 1688980957
transform 1 0 52900 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_573
timestamp 1688980957
transform 1 0 53820 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_577
timestamp 1688980957
transform 1 0 54188 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_605
timestamp 1688980957
transform 1 0 56764 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_610
timestamp 1688980957
transform 1 0 57224 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_29
timestamp 1688980957
transform 1 0 3772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_53
timestamp 1688980957
transform 1 0 5980 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_73
timestamp 1688980957
transform 1 0 7820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_85
timestamp 1688980957
transform 1 0 8924 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_97
timestamp 1688980957
transform 1 0 10028 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_109
timestamp 1688980957
transform 1 0 11132 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_129
timestamp 1688980957
transform 1 0 12972 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_141
timestamp 1688980957
transform 1 0 14076 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_153
timestamp 1688980957
transform 1 0 15180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_165
timestamp 1688980957
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 1688980957
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 1688980957
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 1688980957
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 1688980957
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 1688980957
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 1688980957
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 1688980957
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 1688980957
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 1688980957
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 1688980957
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 1688980957
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_361
timestamp 1688980957
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 1688980957
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 1688980957
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 1688980957
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_405
timestamp 1688980957
transform 1 0 38364 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_411
timestamp 1688980957
transform 1 0 38916 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_417
timestamp 1688980957
transform 1 0 39468 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_421
timestamp 1688980957
transform 1 0 39836 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_425
timestamp 1688980957
transform 1 0 40204 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_469
timestamp 1688980957
transform 1 0 44252 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_477
timestamp 1688980957
transform 1 0 44988 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_485
timestamp 1688980957
transform 1 0 45724 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_489
timestamp 1688980957
transform 1 0 46092 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_501
timestamp 1688980957
transform 1 0 47196 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_505
timestamp 1688980957
transform 1 0 47564 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_516
timestamp 1688980957
transform 1 0 48576 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_540
timestamp 1688980957
transform 1 0 50784 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_558
timestamp 1688980957
transform 1 0 52440 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_561
timestamp 1688980957
transform 1 0 52716 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_566
timestamp 1688980957
transform 1 0 53176 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_570
timestamp 1688980957
transform 1 0 53544 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_581
timestamp 1688980957
transform 1 0 54556 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_586
timestamp 1688980957
transform 1 0 55016 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_596
timestamp 1688980957
transform 1 0 55936 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_608
timestamp 1688980957
transform 1 0 57040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_612
timestamp 1688980957
transform 1 0 57408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_623
timestamp 1688980957
transform 1 0 58420 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_43
timestamp 1688980957
transform 1 0 5060 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_47
timestamp 1688980957
transform 1 0 5428 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_53
timestamp 1688980957
transform 1 0 5980 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_57
timestamp 1688980957
transform 1 0 6348 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_61
timestamp 1688980957
transform 1 0 6716 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_67
timestamp 1688980957
transform 1 0 7268 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_71
timestamp 1688980957
transform 1 0 7636 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_79
timestamp 1688980957
transform 1 0 8372 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_91
timestamp 1688980957
transform 1 0 9476 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_121
timestamp 1688980957
transform 1 0 12236 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_125
timestamp 1688980957
transform 1 0 12604 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_137
timestamp 1688980957
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_157
timestamp 1688980957
transform 1 0 15548 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_178
timestamp 1688980957
transform 1 0 17480 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_182
timestamp 1688980957
transform 1 0 17848 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_194
timestamp 1688980957
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 1688980957
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 1688980957
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 1688980957
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 1688980957
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 1688980957
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 1688980957
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 1688980957
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 1688980957
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 1688980957
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 1688980957
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 1688980957
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 1688980957
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 1688980957
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 1688980957
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 1688980957
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 1688980957
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_401
timestamp 1688980957
transform 1 0 37996 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_410
timestamp 1688980957
transform 1 0 38824 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_418
timestamp 1688980957
transform 1 0 39560 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_425
timestamp 1688980957
transform 1 0 40204 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_448
timestamp 1688980957
transform 1 0 42320 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_454
timestamp 1688980957
transform 1 0 42872 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_458
timestamp 1688980957
transform 1 0 43240 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_462
timestamp 1688980957
transform 1 0 43608 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_474
timestamp 1688980957
transform 1 0 44712 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_477
timestamp 1688980957
transform 1 0 44988 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_481
timestamp 1688980957
transform 1 0 45356 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_486
timestamp 1688980957
transform 1 0 45816 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_490
timestamp 1688980957
transform 1 0 46184 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_494
timestamp 1688980957
transform 1 0 46552 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_531
timestamp 1688980957
transform 1 0 49956 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_533
timestamp 1688980957
transform 1 0 50140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_545
timestamp 1688980957
transform 1 0 51244 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_549
timestamp 1688980957
transform 1 0 51612 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_561
timestamp 1688980957
transform 1 0 52716 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_570
timestamp 1688980957
transform 1 0 53544 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_580
timestamp 1688980957
transform 1 0 54464 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_589
timestamp 1688980957
transform 1 0 55292 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_601
timestamp 1688980957
transform 1 0 56396 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_614
timestamp 1688980957
transform 1 0 57592 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_623
timestamp 1688980957
transform 1 0 58420 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_19
timestamp 1688980957
transform 1 0 2852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_36
timestamp 1688980957
transform 1 0 4416 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_40
timestamp 1688980957
transform 1 0 4784 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_46
timestamp 1688980957
transform 1 0 5336 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_50
timestamp 1688980957
transform 1 0 5704 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_61
timestamp 1688980957
transform 1 0 6716 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_67
timestamp 1688980957
transform 1 0 7268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_79
timestamp 1688980957
transform 1 0 8372 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_86
timestamp 1688980957
transform 1 0 9016 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_90
timestamp 1688980957
transform 1 0 9384 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_94
timestamp 1688980957
transform 1 0 9752 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_106
timestamp 1688980957
transform 1 0 10856 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 1688980957
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 1688980957
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1688980957
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1688980957
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 1688980957
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 1688980957
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 1688980957
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 1688980957
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 1688980957
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 1688980957
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 1688980957
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 1688980957
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 1688980957
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 1688980957
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 1688980957
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 1688980957
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_385
timestamp 1688980957
transform 1 0 36524 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_401
timestamp 1688980957
transform 1 0 37996 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_427
timestamp 1688980957
transform 1 0 40388 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_442
timestamp 1688980957
transform 1 0 41768 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_449
timestamp 1688980957
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_461
timestamp 1688980957
transform 1 0 43516 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_492
timestamp 1688980957
transform 1 0 46368 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_500
timestamp 1688980957
transform 1 0 47104 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_505
timestamp 1688980957
transform 1 0 47564 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_514
timestamp 1688980957
transform 1 0 48392 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_523
timestamp 1688980957
transform 1 0 49220 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_535
timestamp 1688980957
transform 1 0 50324 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_559
timestamp 1688980957
transform 1 0 52532 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_561
timestamp 1688980957
transform 1 0 52716 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_566
timestamp 1688980957
transform 1 0 53176 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_578
timestamp 1688980957
transform 1 0 54280 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_586
timestamp 1688980957
transform 1 0 55016 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_596
timestamp 1688980957
transform 1 0 55936 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_614
timestamp 1688980957
transform 1 0 57592 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_37
timestamp 1688980957
transform 1 0 4508 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_43
timestamp 1688980957
transform 1 0 5060 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_76
timestamp 1688980957
transform 1 0 8096 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_80
timestamp 1688980957
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_118
timestamp 1688980957
transform 1 0 11960 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_130
timestamp 1688980957
transform 1 0 13064 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_138
timestamp 1688980957
transform 1 0 13800 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 1688980957
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 1688980957
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 1688980957
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 1688980957
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 1688980957
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 1688980957
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 1688980957
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 1688980957
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 1688980957
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 1688980957
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 1688980957
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 1688980957
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 1688980957
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 1688980957
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 1688980957
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_377
timestamp 1688980957
transform 1 0 35788 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_381
timestamp 1688980957
transform 1 0 36156 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_441
timestamp 1688980957
transform 1 0 41676 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_451
timestamp 1688980957
transform 1 0 42596 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_467
timestamp 1688980957
transform 1 0 44068 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_472
timestamp 1688980957
transform 1 0 44528 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_477
timestamp 1688980957
transform 1 0 44988 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_481
timestamp 1688980957
transform 1 0 45356 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_505
timestamp 1688980957
transform 1 0 47564 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_517
timestamp 1688980957
transform 1 0 48668 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_522
timestamp 1688980957
transform 1 0 49128 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_527
timestamp 1688980957
transform 1 0 49588 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_533
timestamp 1688980957
transform 1 0 50140 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_537
timestamp 1688980957
transform 1 0 50508 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_558
timestamp 1688980957
transform 1 0 52440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_575
timestamp 1688980957
transform 1 0 54004 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_583
timestamp 1688980957
transform 1 0 54740 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_621
timestamp 1688980957
transform 1 0 58236 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_61
timestamp 1688980957
transform 1 0 6716 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_73
timestamp 1688980957
transform 1 0 7820 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_100
timestamp 1688980957
transform 1 0 10304 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_104
timestamp 1688980957
transform 1 0 10672 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 1688980957
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 1688980957
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 1688980957
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 1688980957
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 1688980957
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 1688980957
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 1688980957
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 1688980957
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 1688980957
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 1688980957
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 1688980957
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 1688980957
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 1688980957
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 1688980957
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 1688980957
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 1688980957
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 1688980957
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 1688980957
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 1688980957
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 1688980957
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_401
timestamp 1688980957
transform 1 0 37996 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_406
timestamp 1688980957
transform 1 0 38456 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_418
timestamp 1688980957
transform 1 0 39560 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_426
timestamp 1688980957
transform 1 0 40296 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_440
timestamp 1688980957
transform 1 0 41584 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_457
timestamp 1688980957
transform 1 0 43148 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_481
timestamp 1688980957
transform 1 0 45356 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_515
timestamp 1688980957
transform 1 0 48484 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_522
timestamp 1688980957
transform 1 0 49128 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_534
timestamp 1688980957
transform 1 0 50232 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_546
timestamp 1688980957
transform 1 0 51336 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_558
timestamp 1688980957
transform 1 0 52440 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_561
timestamp 1688980957
transform 1 0 52716 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_581
timestamp 1688980957
transform 1 0 54556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_585
timestamp 1688980957
transform 1 0 54924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_594
timestamp 1688980957
transform 1 0 55752 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_606
timestamp 1688980957
transform 1 0 56856 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_614
timestamp 1688980957
transform 1 0 57592 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_617
timestamp 1688980957
transform 1 0 57868 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_623
timestamp 1688980957
transform 1 0 58420 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_37
timestamp 1688980957
transform 1 0 4508 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_42
timestamp 1688980957
transform 1 0 4968 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_52
timestamp 1688980957
transform 1 0 5888 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_62
timestamp 1688980957
transform 1 0 6808 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_66
timestamp 1688980957
transform 1 0 7176 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_73
timestamp 1688980957
transform 1 0 7820 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_81
timestamp 1688980957
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 1688980957
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 1688980957
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 1688980957
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 1688980957
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 1688980957
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 1688980957
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 1688980957
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 1688980957
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 1688980957
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 1688980957
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 1688980957
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 1688980957
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 1688980957
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 1688980957
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_401
timestamp 1688980957
transform 1 0 37996 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_413
timestamp 1688980957
transform 1 0 39100 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_419
timestamp 1688980957
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_421
timestamp 1688980957
transform 1 0 39836 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_425
timestamp 1688980957
transform 1 0 40204 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_474
timestamp 1688980957
transform 1 0 44712 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_488
timestamp 1688980957
transform 1 0 46000 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_492
timestamp 1688980957
transform 1 0 46368 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_504
timestamp 1688980957
transform 1 0 47472 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_533
timestamp 1688980957
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_547
timestamp 1688980957
transform 1 0 51428 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_559
timestamp 1688980957
transform 1 0 52532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_571
timestamp 1688980957
transform 1 0 53636 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_583
timestamp 1688980957
transform 1 0 54740 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_587
timestamp 1688980957
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_589
timestamp 1688980957
transform 1 0 55292 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_597
timestamp 1688980957
transform 1 0 56028 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_606
timestamp 1688980957
transform 1 0 56856 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_613
timestamp 1688980957
transform 1 0 57500 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_621
timestamp 1688980957
transform 1 0 58236 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_21
timestamp 1688980957
transform 1 0 3036 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_50
timestamp 1688980957
transform 1 0 5704 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_60
timestamp 1688980957
transform 1 0 6624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_83
timestamp 1688980957
transform 1 0 8740 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_97
timestamp 1688980957
transform 1 0 10028 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_101
timestamp 1688980957
transform 1 0 10396 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 1688980957
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 1688980957
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 1688980957
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 1688980957
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 1688980957
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 1688980957
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 1688980957
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 1688980957
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 1688980957
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 1688980957
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 1688980957
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 1688980957
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 1688980957
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 1688980957
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 1688980957
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 1688980957
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 1688980957
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 1688980957
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 1688980957
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_393
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_405
timestamp 1688980957
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_417
timestamp 1688980957
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_429
timestamp 1688980957
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_441
timestamp 1688980957
transform 1 0 41676 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_471
timestamp 1688980957
transform 1 0 44436 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_501
timestamp 1688980957
transform 1 0 47196 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_528
timestamp 1688980957
transform 1 0 49680 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_532
timestamp 1688980957
transform 1 0 50048 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_556
timestamp 1688980957
transform 1 0 52256 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_561
timestamp 1688980957
transform 1 0 52716 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_573
timestamp 1688980957
transform 1 0 53820 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_585
timestamp 1688980957
transform 1 0 54924 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_595
timestamp 1688980957
transform 1 0 55844 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_603
timestamp 1688980957
transform 1 0 56580 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_620
timestamp 1688980957
transform 1 0 58144 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_26
timestamp 1688980957
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_37
timestamp 1688980957
transform 1 0 4508 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_43
timestamp 1688980957
transform 1 0 5060 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_65
timestamp 1688980957
transform 1 0 7084 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_69
timestamp 1688980957
transform 1 0 7452 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_81
timestamp 1688980957
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_105
timestamp 1688980957
transform 1 0 10764 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_117
timestamp 1688980957
transform 1 0 11868 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_129
timestamp 1688980957
transform 1 0 12972 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_137
timestamp 1688980957
transform 1 0 13708 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1688980957
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 1688980957
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 1688980957
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 1688980957
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 1688980957
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 1688980957
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 1688980957
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 1688980957
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 1688980957
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 1688980957
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 1688980957
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 1688980957
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 1688980957
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 1688980957
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 1688980957
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_401
timestamp 1688980957
transform 1 0 37996 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_413
timestamp 1688980957
transform 1 0 39100 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_419
timestamp 1688980957
transform 1 0 39652 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_421
timestamp 1688980957
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_433
timestamp 1688980957
transform 1 0 40940 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_439
timestamp 1688980957
transform 1 0 41492 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_471
timestamp 1688980957
transform 1 0 44436 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_475
timestamp 1688980957
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_477
timestamp 1688980957
transform 1 0 44988 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_481
timestamp 1688980957
transform 1 0 45356 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_485
timestamp 1688980957
transform 1 0 45724 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_491
timestamp 1688980957
transform 1 0 46276 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_494
timestamp 1688980957
transform 1 0 46552 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_506
timestamp 1688980957
transform 1 0 47656 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_518
timestamp 1688980957
transform 1 0 48760 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_530
timestamp 1688980957
transform 1 0 49864 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_541
timestamp 1688980957
transform 1 0 50876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_553
timestamp 1688980957
transform 1 0 51980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_565
timestamp 1688980957
transform 1 0 53084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_577
timestamp 1688980957
transform 1 0 54188 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_585
timestamp 1688980957
transform 1 0 54924 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_589
timestamp 1688980957
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_601
timestamp 1688980957
transform 1 0 56396 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_609
timestamp 1688980957
transform 1 0 57132 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_613
timestamp 1688980957
transform 1 0 57500 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_623
timestamp 1688980957
transform 1 0 58420 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_31
timestamp 1688980957
transform 1 0 3956 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_35
timestamp 1688980957
transform 1 0 4324 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_40
timestamp 1688980957
transform 1 0 4784 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_52
timestamp 1688980957
transform 1 0 5888 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 1688980957
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 1688980957
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 1688980957
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 1688980957
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 1688980957
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 1688980957
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 1688980957
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 1688980957
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 1688980957
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 1688980957
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 1688980957
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 1688980957
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1688980957
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_405
timestamp 1688980957
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_417
timestamp 1688980957
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_429
timestamp 1688980957
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_441
timestamp 1688980957
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_447
timestamp 1688980957
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_449
timestamp 1688980957
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_461
timestamp 1688980957
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_473
timestamp 1688980957
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_485
timestamp 1688980957
transform 1 0 45724 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_497
timestamp 1688980957
transform 1 0 46828 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_503
timestamp 1688980957
transform 1 0 47380 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_505
timestamp 1688980957
transform 1 0 47564 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_517
timestamp 1688980957
transform 1 0 48668 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_547
timestamp 1688980957
transform 1 0 51428 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_551
timestamp 1688980957
transform 1 0 51796 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_555
timestamp 1688980957
transform 1 0 52164 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_559
timestamp 1688980957
transform 1 0 52532 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_561
timestamp 1688980957
transform 1 0 52716 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_573
timestamp 1688980957
transform 1 0 53820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_585
timestamp 1688980957
transform 1 0 54924 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_596
timestamp 1688980957
transform 1 0 55936 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_607
timestamp 1688980957
transform 1 0 56948 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_617
timestamp 1688980957
transform 1 0 57868 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_621
timestamp 1688980957
transform 1 0 58236 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_11
timestamp 1688980957
transform 1 0 2116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_22
timestamp 1688980957
transform 1 0 3128 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_32
timestamp 1688980957
transform 1 0 4048 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_38
timestamp 1688980957
transform 1 0 4600 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_58
timestamp 1688980957
transform 1 0 6440 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_70
timestamp 1688980957
transform 1 0 7544 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 1688980957
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 1688980957
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 1688980957
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 1688980957
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 1688980957
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 1688980957
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 1688980957
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 1688980957
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 1688980957
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 1688980957
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 1688980957
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 1688980957
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 1688980957
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 1688980957
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 1688980957
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1688980957
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1688980957
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_401
timestamp 1688980957
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_413
timestamp 1688980957
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_419
timestamp 1688980957
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_421
timestamp 1688980957
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_433
timestamp 1688980957
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_445
timestamp 1688980957
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_457
timestamp 1688980957
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_469
timestamp 1688980957
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_475
timestamp 1688980957
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_477
timestamp 1688980957
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_489
timestamp 1688980957
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_501
timestamp 1688980957
transform 1 0 47196 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_513
timestamp 1688980957
transform 1 0 48300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_525
timestamp 1688980957
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_531
timestamp 1688980957
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_533
timestamp 1688980957
transform 1 0 50140 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_545
timestamp 1688980957
transform 1 0 51244 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_557
timestamp 1688980957
transform 1 0 52348 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_569
timestamp 1688980957
transform 1 0 53452 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_581
timestamp 1688980957
transform 1 0 54556 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_587
timestamp 1688980957
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_589
timestamp 1688980957
transform 1 0 55292 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_601
timestamp 1688980957
transform 1 0 56396 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_605
timestamp 1688980957
transform 1 0 56764 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_621
timestamp 1688980957
transform 1 0 58236 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_31
timestamp 1688980957
transform 1 0 3956 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_86
timestamp 1688980957
transform 1 0 9016 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_90
timestamp 1688980957
transform 1 0 9384 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_102
timestamp 1688980957
transform 1 0 10488 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_110
timestamp 1688980957
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1688980957
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 1688980957
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 1688980957
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 1688980957
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 1688980957
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 1688980957
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 1688980957
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 1688980957
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 1688980957
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 1688980957
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 1688980957
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 1688980957
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 1688980957
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 1688980957
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_405
timestamp 1688980957
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_417
timestamp 1688980957
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_429
timestamp 1688980957
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_441
timestamp 1688980957
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_447
timestamp 1688980957
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_449
timestamp 1688980957
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_461
timestamp 1688980957
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_473
timestamp 1688980957
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_485
timestamp 1688980957
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_497
timestamp 1688980957
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_503
timestamp 1688980957
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_505
timestamp 1688980957
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_517
timestamp 1688980957
transform 1 0 48668 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_529
timestamp 1688980957
transform 1 0 49772 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_541
timestamp 1688980957
transform 1 0 50876 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_553
timestamp 1688980957
transform 1 0 51980 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_559
timestamp 1688980957
transform 1 0 52532 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_561
timestamp 1688980957
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_573
timestamp 1688980957
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_585
timestamp 1688980957
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_597
timestamp 1688980957
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_609
timestamp 1688980957
transform 1 0 57132 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_613
timestamp 1688980957
transform 1 0 57500 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_624
timestamp 1688980957
transform 1 0 58512 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_26
timestamp 1688980957
transform 1 0 3496 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_33
timestamp 1688980957
transform 1 0 4140 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_45
timestamp 1688980957
transform 1 0 5244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_57
timestamp 1688980957
transform 1 0 6348 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_74
timestamp 1688980957
transform 1 0 7912 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_79
timestamp 1688980957
transform 1 0 8372 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 1688980957
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 1688980957
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1688980957
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 1688980957
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 1688980957
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 1688980957
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 1688980957
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 1688980957
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 1688980957
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 1688980957
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1688980957
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 1688980957
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 1688980957
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 1688980957
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 1688980957
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 1688980957
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 1688980957
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1688980957
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_401
timestamp 1688980957
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_413
timestamp 1688980957
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_419
timestamp 1688980957
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_421
timestamp 1688980957
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_433
timestamp 1688980957
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_445
timestamp 1688980957
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_457
timestamp 1688980957
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_469
timestamp 1688980957
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_475
timestamp 1688980957
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_477
timestamp 1688980957
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_489
timestamp 1688980957
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_501
timestamp 1688980957
transform 1 0 47196 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_513
timestamp 1688980957
transform 1 0 48300 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_525
timestamp 1688980957
transform 1 0 49404 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_531
timestamp 1688980957
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_533
timestamp 1688980957
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_545
timestamp 1688980957
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_557
timestamp 1688980957
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_569
timestamp 1688980957
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_581
timestamp 1688980957
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_587
timestamp 1688980957
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_589
timestamp 1688980957
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_601
timestamp 1688980957
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_617
timestamp 1688980957
transform 1 0 57868 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_621
timestamp 1688980957
transform 1 0 58236 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_29
timestamp 1688980957
transform 1 0 3772 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_103
timestamp 1688980957
transform 1 0 10580 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_107
timestamp 1688980957
transform 1 0 10948 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1688980957
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 1688980957
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 1688980957
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 1688980957
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 1688980957
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 1688980957
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 1688980957
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 1688980957
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 1688980957
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 1688980957
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 1688980957
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 1688980957
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1688980957
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1688980957
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 1688980957
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 1688980957
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 1688980957
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 1688980957
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 1688980957
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_405
timestamp 1688980957
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_417
timestamp 1688980957
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_429
timestamp 1688980957
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_441
timestamp 1688980957
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_447
timestamp 1688980957
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_449
timestamp 1688980957
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_461
timestamp 1688980957
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_473
timestamp 1688980957
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_485
timestamp 1688980957
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_497
timestamp 1688980957
transform 1 0 46828 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_503
timestamp 1688980957
transform 1 0 47380 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_505
timestamp 1688980957
transform 1 0 47564 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_517
timestamp 1688980957
transform 1 0 48668 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_529
timestamp 1688980957
transform 1 0 49772 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_541
timestamp 1688980957
transform 1 0 50876 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_553
timestamp 1688980957
transform 1 0 51980 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_559
timestamp 1688980957
transform 1 0 52532 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_561
timestamp 1688980957
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_573
timestamp 1688980957
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_585
timestamp 1688980957
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_597
timestamp 1688980957
transform 1 0 56028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_609
timestamp 1688980957
transform 1 0 57132 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_613
timestamp 1688980957
transform 1 0 57500 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_620
timestamp 1688980957
transform 1 0 58144 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_19
timestamp 1688980957
transform 1 0 2852 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_46
timestamp 1688980957
transform 1 0 5336 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_80
timestamp 1688980957
transform 1 0 8464 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_93
timestamp 1688980957
transform 1 0 9660 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_105
timestamp 1688980957
transform 1 0 10764 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_117
timestamp 1688980957
transform 1 0 11868 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_129
timestamp 1688980957
transform 1 0 12972 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_137
timestamp 1688980957
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_177
timestamp 1688980957
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_189
timestamp 1688980957
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_195
timestamp 1688980957
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 1688980957
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_221
timestamp 1688980957
transform 1 0 21436 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_233
timestamp 1688980957
transform 1 0 22540 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_245
timestamp 1688980957
transform 1 0 23644 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_251
timestamp 1688980957
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 1688980957
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_277
timestamp 1688980957
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_289
timestamp 1688980957
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_301
timestamp 1688980957
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_307
timestamp 1688980957
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 1688980957
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_333
timestamp 1688980957
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_345
timestamp 1688980957
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 1688980957
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1688980957
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1688980957
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_401
timestamp 1688980957
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_413
timestamp 1688980957
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_419
timestamp 1688980957
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_421
timestamp 1688980957
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_433
timestamp 1688980957
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_445
timestamp 1688980957
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_457
timestamp 1688980957
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_469
timestamp 1688980957
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_475
timestamp 1688980957
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_477
timestamp 1688980957
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_489
timestamp 1688980957
transform 1 0 46092 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_501
timestamp 1688980957
transform 1 0 47196 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_513
timestamp 1688980957
transform 1 0 48300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_525
timestamp 1688980957
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_531
timestamp 1688980957
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_533
timestamp 1688980957
transform 1 0 50140 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_545
timestamp 1688980957
transform 1 0 51244 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_557
timestamp 1688980957
transform 1 0 52348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_569
timestamp 1688980957
transform 1 0 53452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_581
timestamp 1688980957
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_587
timestamp 1688980957
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_589
timestamp 1688980957
transform 1 0 55292 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_601
timestamp 1688980957
transform 1 0 56396 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_613
timestamp 1688980957
transform 1 0 57500 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_621
timestamp 1688980957
transform 1 0 58236 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_31
timestamp 1688980957
transform 1 0 3956 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_40
timestamp 1688980957
transform 1 0 4784 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_52
timestamp 1688980957
transform 1 0 5888 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_71
timestamp 1688980957
transform 1 0 7636 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_82
timestamp 1688980957
transform 1 0 8648 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_92
timestamp 1688980957
transform 1 0 9568 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_104
timestamp 1688980957
transform 1 0 10672 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_137
timestamp 1688980957
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 1688980957
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_161
timestamp 1688980957
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 1688980957
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_181
timestamp 1688980957
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_193
timestamp 1688980957
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_205
timestamp 1688980957
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_217
timestamp 1688980957
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 1688980957
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_237
timestamp 1688980957
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_249
timestamp 1688980957
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_261
timestamp 1688980957
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_273
timestamp 1688980957
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_279
timestamp 1688980957
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_281
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_293
timestamp 1688980957
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_305
timestamp 1688980957
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_317
timestamp 1688980957
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_329
timestamp 1688980957
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_335
timestamp 1688980957
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1688980957
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 1688980957
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 1688980957
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 1688980957
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 1688980957
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_393
timestamp 1688980957
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_405
timestamp 1688980957
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_417
timestamp 1688980957
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_429
timestamp 1688980957
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_441
timestamp 1688980957
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_447
timestamp 1688980957
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_449
timestamp 1688980957
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_461
timestamp 1688980957
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_473
timestamp 1688980957
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_485
timestamp 1688980957
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_497
timestamp 1688980957
transform 1 0 46828 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_503
timestamp 1688980957
transform 1 0 47380 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_505
timestamp 1688980957
transform 1 0 47564 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_517
timestamp 1688980957
transform 1 0 48668 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_529
timestamp 1688980957
transform 1 0 49772 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_541
timestamp 1688980957
transform 1 0 50876 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_553
timestamp 1688980957
transform 1 0 51980 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_559
timestamp 1688980957
transform 1 0 52532 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_561
timestamp 1688980957
transform 1 0 52716 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_573
timestamp 1688980957
transform 1 0 53820 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_585
timestamp 1688980957
transform 1 0 54924 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_597
timestamp 1688980957
transform 1 0 56028 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_609
timestamp 1688980957
transform 1 0 57132 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_613
timestamp 1688980957
transform 1 0 57500 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_624
timestamp 1688980957
transform 1 0 58512 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_7
timestamp 1688980957
transform 1 0 1748 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_33
timestamp 1688980957
transform 1 0 4140 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_45
timestamp 1688980957
transform 1 0 5244 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_53
timestamp 1688980957
transform 1 0 5980 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_71
timestamp 1688980957
transform 1 0 7636 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_106
timestamp 1688980957
transform 1 0 10856 0 1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_110
timestamp 1688980957
transform 1 0 11224 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_122
timestamp 1688980957
transform 1 0 12328 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_134
timestamp 1688980957
transform 1 0 13432 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1688980957
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 1688980957
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1688980957
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_209
timestamp 1688980957
transform 1 0 20332 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_221
timestamp 1688980957
transform 1 0 21436 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_233
timestamp 1688980957
transform 1 0 22540 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_245
timestamp 1688980957
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 1688980957
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_253
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_265
timestamp 1688980957
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_277
timestamp 1688980957
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_289
timestamp 1688980957
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_301
timestamp 1688980957
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 1688980957
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_309
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_321
timestamp 1688980957
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_333
timestamp 1688980957
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_345
timestamp 1688980957
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_357
timestamp 1688980957
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1688980957
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_365
timestamp 1688980957
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_377
timestamp 1688980957
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_389
timestamp 1688980957
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_401
timestamp 1688980957
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_413
timestamp 1688980957
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_419
timestamp 1688980957
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_421
timestamp 1688980957
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_433
timestamp 1688980957
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_445
timestamp 1688980957
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_457
timestamp 1688980957
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_469
timestamp 1688980957
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_475
timestamp 1688980957
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_477
timestamp 1688980957
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_489
timestamp 1688980957
transform 1 0 46092 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_501
timestamp 1688980957
transform 1 0 47196 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_513
timestamp 1688980957
transform 1 0 48300 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_525
timestamp 1688980957
transform 1 0 49404 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_531
timestamp 1688980957
transform 1 0 49956 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_533
timestamp 1688980957
transform 1 0 50140 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_545
timestamp 1688980957
transform 1 0 51244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_557
timestamp 1688980957
transform 1 0 52348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_569
timestamp 1688980957
transform 1 0 53452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_581
timestamp 1688980957
transform 1 0 54556 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_587
timestamp 1688980957
transform 1 0 55108 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_589
timestamp 1688980957
transform 1 0 55292 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_601
timestamp 1688980957
transform 1 0 56396 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_623
timestamp 1688980957
transform 1 0 58420 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_49
timestamp 1688980957
transform 1 0 5612 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_55
timestamp 1688980957
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_89
timestamp 1688980957
transform 1 0 9292 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_98
timestamp 1688980957
transform 1 0 10120 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_110
timestamp 1688980957
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_125
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_137
timestamp 1688980957
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_149
timestamp 1688980957
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 1688980957
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1688980957
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_181
timestamp 1688980957
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_193
timestamp 1688980957
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_205
timestamp 1688980957
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_217
timestamp 1688980957
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_223
timestamp 1688980957
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_237
timestamp 1688980957
transform 1 0 22908 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_249
timestamp 1688980957
transform 1 0 24012 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_261
timestamp 1688980957
transform 1 0 25116 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_273
timestamp 1688980957
transform 1 0 26220 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_279
timestamp 1688980957
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_281
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_293
timestamp 1688980957
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_305
timestamp 1688980957
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_317
timestamp 1688980957
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 1688980957
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 1688980957
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_337
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_349
timestamp 1688980957
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_361
timestamp 1688980957
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_373
timestamp 1688980957
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_385
timestamp 1688980957
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_391
timestamp 1688980957
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_393
timestamp 1688980957
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_405
timestamp 1688980957
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_417
timestamp 1688980957
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_429
timestamp 1688980957
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_441
timestamp 1688980957
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_447
timestamp 1688980957
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_449
timestamp 1688980957
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_461
timestamp 1688980957
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_473
timestamp 1688980957
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_485
timestamp 1688980957
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_497
timestamp 1688980957
transform 1 0 46828 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_503
timestamp 1688980957
transform 1 0 47380 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_505
timestamp 1688980957
transform 1 0 47564 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_517
timestamp 1688980957
transform 1 0 48668 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_529
timestamp 1688980957
transform 1 0 49772 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_541
timestamp 1688980957
transform 1 0 50876 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_553
timestamp 1688980957
transform 1 0 51980 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_559
timestamp 1688980957
transform 1 0 52532 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_561
timestamp 1688980957
transform 1 0 52716 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_573
timestamp 1688980957
transform 1 0 53820 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_585
timestamp 1688980957
transform 1 0 54924 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_597
timestamp 1688980957
transform 1 0 56028 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_609
timestamp 1688980957
transform 1 0 57132 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_613
timestamp 1688980957
transform 1 0 57500 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_617
timestamp 1688980957
transform 1 0 57868 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_624
timestamp 1688980957
transform 1 0 58512 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_26
timestamp 1688980957
transform 1 0 3496 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_48
timestamp 1688980957
transform 1 0 5520 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_56
timestamp 1688980957
transform 1 0 6256 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_67
timestamp 1688980957
transform 1 0 7268 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_75
timestamp 1688980957
transform 1 0 8004 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_93
timestamp 1688980957
transform 1 0 9660 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_105
timestamp 1688980957
transform 1 0 10764 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_117
timestamp 1688980957
transform 1 0 11868 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_129
timestamp 1688980957
transform 1 0 12972 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_137
timestamp 1688980957
transform 1 0 13708 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 1688980957
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 1688980957
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_189
timestamp 1688980957
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_195
timestamp 1688980957
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_209
timestamp 1688980957
transform 1 0 20332 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_221
timestamp 1688980957
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_233
timestamp 1688980957
transform 1 0 22540 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_245
timestamp 1688980957
transform 1 0 23644 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_251
timestamp 1688980957
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_253
timestamp 1688980957
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_265
timestamp 1688980957
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_277
timestamp 1688980957
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_289
timestamp 1688980957
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_301
timestamp 1688980957
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_307
timestamp 1688980957
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_309
timestamp 1688980957
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_321
timestamp 1688980957
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_333
timestamp 1688980957
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_345
timestamp 1688980957
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_357
timestamp 1688980957
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_363
timestamp 1688980957
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_365
timestamp 1688980957
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_377
timestamp 1688980957
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_389
timestamp 1688980957
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_401
timestamp 1688980957
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_413
timestamp 1688980957
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_419
timestamp 1688980957
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_421
timestamp 1688980957
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_433
timestamp 1688980957
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_445
timestamp 1688980957
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_457
timestamp 1688980957
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_469
timestamp 1688980957
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_475
timestamp 1688980957
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_477
timestamp 1688980957
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_489
timestamp 1688980957
transform 1 0 46092 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_501
timestamp 1688980957
transform 1 0 47196 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_513
timestamp 1688980957
transform 1 0 48300 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_525
timestamp 1688980957
transform 1 0 49404 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_531
timestamp 1688980957
transform 1 0 49956 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_533
timestamp 1688980957
transform 1 0 50140 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_545
timestamp 1688980957
transform 1 0 51244 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_557
timestamp 1688980957
transform 1 0 52348 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_569
timestamp 1688980957
transform 1 0 53452 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_581
timestamp 1688980957
transform 1 0 54556 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_587
timestamp 1688980957
transform 1 0 55108 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_589
timestamp 1688980957
transform 1 0 55292 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_601
timestamp 1688980957
transform 1 0 56396 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_607
timestamp 1688980957
transform 1 0 56948 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_7
timestamp 1688980957
transform 1 0 1748 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_28
timestamp 1688980957
transform 1 0 3680 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_40
timestamp 1688980957
transform 1 0 4784 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_52
timestamp 1688980957
transform 1 0 5888 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_69
timestamp 1688980957
transform 1 0 7452 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_110
timestamp 1688980957
transform 1 0 11224 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_117
timestamp 1688980957
transform 1 0 11868 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_129
timestamp 1688980957
transform 1 0 12972 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_141
timestamp 1688980957
transform 1 0 14076 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_153
timestamp 1688980957
transform 1 0 15180 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_165
timestamp 1688980957
transform 1 0 16284 0 -1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 1688980957
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_193
timestamp 1688980957
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_205
timestamp 1688980957
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_217
timestamp 1688980957
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_223
timestamp 1688980957
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_225
timestamp 1688980957
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_237
timestamp 1688980957
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_249
timestamp 1688980957
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_261
timestamp 1688980957
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_273
timestamp 1688980957
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_279
timestamp 1688980957
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_281
timestamp 1688980957
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_293
timestamp 1688980957
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_305
timestamp 1688980957
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_317
timestamp 1688980957
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_329
timestamp 1688980957
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_335
timestamp 1688980957
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_337
timestamp 1688980957
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_349
timestamp 1688980957
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_361
timestamp 1688980957
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_373
timestamp 1688980957
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_385
timestamp 1688980957
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_391
timestamp 1688980957
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_393
timestamp 1688980957
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_405
timestamp 1688980957
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_417
timestamp 1688980957
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_429
timestamp 1688980957
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_441
timestamp 1688980957
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_447
timestamp 1688980957
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_449
timestamp 1688980957
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_461
timestamp 1688980957
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_473
timestamp 1688980957
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_485
timestamp 1688980957
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_497
timestamp 1688980957
transform 1 0 46828 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_503
timestamp 1688980957
transform 1 0 47380 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_505
timestamp 1688980957
transform 1 0 47564 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_517
timestamp 1688980957
transform 1 0 48668 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_529
timestamp 1688980957
transform 1 0 49772 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_541
timestamp 1688980957
transform 1 0 50876 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_553
timestamp 1688980957
transform 1 0 51980 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_559
timestamp 1688980957
transform 1 0 52532 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_561
timestamp 1688980957
transform 1 0 52716 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_573
timestamp 1688980957
transform 1 0 53820 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_585
timestamp 1688980957
transform 1 0 54924 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_597
timestamp 1688980957
transform 1 0 56028 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_609
timestamp 1688980957
transform 1 0 57132 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_617
timestamp 1688980957
transform 1 0 57868 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_623
timestamp 1688980957
transform 1 0 58420 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_3
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_15
timestamp 1688980957
transform 1 0 2484 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_25
timestamp 1688980957
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_53
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_65
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 1688980957
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 1688980957
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 1688980957
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 1688980957
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 1688980957
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 1688980957
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_165
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_177
timestamp 1688980957
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_189
timestamp 1688980957
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_195
timestamp 1688980957
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_197
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_209
timestamp 1688980957
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_221
timestamp 1688980957
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_233
timestamp 1688980957
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_245
timestamp 1688980957
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_251
timestamp 1688980957
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_253
timestamp 1688980957
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_265
timestamp 1688980957
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_277
timestamp 1688980957
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_289
timestamp 1688980957
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_301
timestamp 1688980957
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_307
timestamp 1688980957
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_309
timestamp 1688980957
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_321
timestamp 1688980957
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_333
timestamp 1688980957
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_345
timestamp 1688980957
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_357
timestamp 1688980957
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_363
timestamp 1688980957
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_365
timestamp 1688980957
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_377
timestamp 1688980957
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_389
timestamp 1688980957
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_401
timestamp 1688980957
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_413
timestamp 1688980957
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_419
timestamp 1688980957
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_421
timestamp 1688980957
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_433
timestamp 1688980957
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_445
timestamp 1688980957
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_457
timestamp 1688980957
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_469
timestamp 1688980957
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_475
timestamp 1688980957
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_477
timestamp 1688980957
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_489
timestamp 1688980957
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_501
timestamp 1688980957
transform 1 0 47196 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_513
timestamp 1688980957
transform 1 0 48300 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_525
timestamp 1688980957
transform 1 0 49404 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_531
timestamp 1688980957
transform 1 0 49956 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_533
timestamp 1688980957
transform 1 0 50140 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_545
timestamp 1688980957
transform 1 0 51244 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_557
timestamp 1688980957
transform 1 0 52348 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_569
timestamp 1688980957
transform 1 0 53452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_581
timestamp 1688980957
transform 1 0 54556 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_587
timestamp 1688980957
transform 1 0 55108 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_589
timestamp 1688980957
transform 1 0 55292 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_601
timestamp 1688980957
transform 1 0 56396 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_613
timestamp 1688980957
transform 1 0 57500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_623
timestamp 1688980957
transform 1 0 58420 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_19
timestamp 1688980957
transform 1 0 2852 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_31
timestamp 1688980957
transform 1 0 3956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_43
timestamp 1688980957
transform 1 0 5060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1688980957
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 1688980957
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_93
timestamp 1688980957
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_105
timestamp 1688980957
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_111
timestamp 1688980957
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 1688980957
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 1688980957
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 1688980957
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1688980957
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_193
timestamp 1688980957
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_205
timestamp 1688980957
transform 1 0 19964 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_217
timestamp 1688980957
transform 1 0 21068 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_223
timestamp 1688980957
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_225
timestamp 1688980957
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_237
timestamp 1688980957
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_249
timestamp 1688980957
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_261
timestamp 1688980957
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_273
timestamp 1688980957
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_279
timestamp 1688980957
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_281
timestamp 1688980957
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_293
timestamp 1688980957
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_305
timestamp 1688980957
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_317
timestamp 1688980957
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_329
timestamp 1688980957
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_335
timestamp 1688980957
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_337
timestamp 1688980957
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_349
timestamp 1688980957
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_361
timestamp 1688980957
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_373
timestamp 1688980957
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_385
timestamp 1688980957
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_391
timestamp 1688980957
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_393
timestamp 1688980957
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_405
timestamp 1688980957
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_417
timestamp 1688980957
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_429
timestamp 1688980957
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_441
timestamp 1688980957
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_447
timestamp 1688980957
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_449
timestamp 1688980957
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_461
timestamp 1688980957
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_473
timestamp 1688980957
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_485
timestamp 1688980957
transform 1 0 45724 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_497
timestamp 1688980957
transform 1 0 46828 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_503
timestamp 1688980957
transform 1 0 47380 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_505
timestamp 1688980957
transform 1 0 47564 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_517
timestamp 1688980957
transform 1 0 48668 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_529
timestamp 1688980957
transform 1 0 49772 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_541
timestamp 1688980957
transform 1 0 50876 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_553
timestamp 1688980957
transform 1 0 51980 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_559
timestamp 1688980957
transform 1 0 52532 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_561
timestamp 1688980957
transform 1 0 52716 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_573
timestamp 1688980957
transform 1 0 53820 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_585
timestamp 1688980957
transform 1 0 54924 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_597
timestamp 1688980957
transform 1 0 56028 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_609
timestamp 1688980957
transform 1 0 57132 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_615
timestamp 1688980957
transform 1 0 57684 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_624
timestamp 1688980957
transform 1 0 58512 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_15
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_53
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_77
timestamp 1688980957
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_83
timestamp 1688980957
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1688980957
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1688980957
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1688980957
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 1688980957
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 1688980957
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_177
timestamp 1688980957
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_189
timestamp 1688980957
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_195
timestamp 1688980957
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_197
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_209
timestamp 1688980957
transform 1 0 20332 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_221
timestamp 1688980957
transform 1 0 21436 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_233
timestamp 1688980957
transform 1 0 22540 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_245
timestamp 1688980957
transform 1 0 23644 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_251
timestamp 1688980957
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_253
timestamp 1688980957
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_265
timestamp 1688980957
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_277
timestamp 1688980957
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_289
timestamp 1688980957
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_301
timestamp 1688980957
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_307
timestamp 1688980957
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_309
timestamp 1688980957
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_321
timestamp 1688980957
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_333
timestamp 1688980957
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_345
timestamp 1688980957
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_357
timestamp 1688980957
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_363
timestamp 1688980957
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_365
timestamp 1688980957
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_377
timestamp 1688980957
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_389
timestamp 1688980957
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_401
timestamp 1688980957
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_413
timestamp 1688980957
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_419
timestamp 1688980957
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_421
timestamp 1688980957
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_433
timestamp 1688980957
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_445
timestamp 1688980957
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_457
timestamp 1688980957
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_469
timestamp 1688980957
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_475
timestamp 1688980957
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_477
timestamp 1688980957
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_489
timestamp 1688980957
transform 1 0 46092 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_501
timestamp 1688980957
transform 1 0 47196 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_513
timestamp 1688980957
transform 1 0 48300 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_525
timestamp 1688980957
transform 1 0 49404 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_531
timestamp 1688980957
transform 1 0 49956 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_533
timestamp 1688980957
transform 1 0 50140 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_545
timestamp 1688980957
transform 1 0 51244 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_557
timestamp 1688980957
transform 1 0 52348 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_569
timestamp 1688980957
transform 1 0 53452 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_581
timestamp 1688980957
transform 1 0 54556 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_587
timestamp 1688980957
transform 1 0 55108 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_589
timestamp 1688980957
transform 1 0 55292 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_601
timestamp 1688980957
transform 1 0 56396 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_613
timestamp 1688980957
transform 1 0 57500 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_15
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_27
timestamp 1688980957
transform 1 0 3588 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_39
timestamp 1688980957
transform 1 0 4692 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73_51
timestamp 1688980957
transform 1 0 5796 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_55
timestamp 1688980957
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_69
timestamp 1688980957
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_81
timestamp 1688980957
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_93
timestamp 1688980957
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_105
timestamp 1688980957
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_111
timestamp 1688980957
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_149
timestamp 1688980957
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_161
timestamp 1688980957
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 1688980957
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 1688980957
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_193
timestamp 1688980957
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_205
timestamp 1688980957
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_217
timestamp 1688980957
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_223
timestamp 1688980957
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_225
timestamp 1688980957
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_237
timestamp 1688980957
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_249
timestamp 1688980957
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_261
timestamp 1688980957
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_273
timestamp 1688980957
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_279
timestamp 1688980957
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_281
timestamp 1688980957
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_293
timestamp 1688980957
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_305
timestamp 1688980957
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_317
timestamp 1688980957
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_329
timestamp 1688980957
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_335
timestamp 1688980957
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_337
timestamp 1688980957
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_349
timestamp 1688980957
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_361
timestamp 1688980957
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_373
timestamp 1688980957
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_385
timestamp 1688980957
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_391
timestamp 1688980957
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_393
timestamp 1688980957
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_405
timestamp 1688980957
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_417
timestamp 1688980957
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_429
timestamp 1688980957
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_441
timestamp 1688980957
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_447
timestamp 1688980957
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_449
timestamp 1688980957
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_461
timestamp 1688980957
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_473
timestamp 1688980957
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_485
timestamp 1688980957
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_497
timestamp 1688980957
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_503
timestamp 1688980957
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_505
timestamp 1688980957
transform 1 0 47564 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_517
timestamp 1688980957
transform 1 0 48668 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_529
timestamp 1688980957
transform 1 0 49772 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_541
timestamp 1688980957
transform 1 0 50876 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_553
timestamp 1688980957
transform 1 0 51980 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_559
timestamp 1688980957
transform 1 0 52532 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_561
timestamp 1688980957
transform 1 0 52716 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_573
timestamp 1688980957
transform 1 0 53820 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_585
timestamp 1688980957
transform 1 0 54924 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_597
timestamp 1688980957
transform 1 0 56028 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_617
timestamp 1688980957
transform 1 0 57868 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_74_19
timestamp 1688980957
transform 1 0 2852 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_27
timestamp 1688980957
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_41
timestamp 1688980957
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_53
timestamp 1688980957
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_65
timestamp 1688980957
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_77
timestamp 1688980957
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_83
timestamp 1688980957
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_85
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 1688980957
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1688980957
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 1688980957
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 1688980957
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1688980957
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_153
timestamp 1688980957
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_165
timestamp 1688980957
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_177
timestamp 1688980957
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_189
timestamp 1688980957
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_195
timestamp 1688980957
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_197
timestamp 1688980957
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_209
timestamp 1688980957
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_221
timestamp 1688980957
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_233
timestamp 1688980957
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_245
timestamp 1688980957
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_251
timestamp 1688980957
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_253
timestamp 1688980957
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_265
timestamp 1688980957
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_277
timestamp 1688980957
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_289
timestamp 1688980957
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_301
timestamp 1688980957
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_307
timestamp 1688980957
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_309
timestamp 1688980957
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_321
timestamp 1688980957
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_333
timestamp 1688980957
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_345
timestamp 1688980957
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_357
timestamp 1688980957
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_363
timestamp 1688980957
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_365
timestamp 1688980957
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_377
timestamp 1688980957
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_389
timestamp 1688980957
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_401
timestamp 1688980957
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_413
timestamp 1688980957
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_419
timestamp 1688980957
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_421
timestamp 1688980957
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_433
timestamp 1688980957
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_445
timestamp 1688980957
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_457
timestamp 1688980957
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_469
timestamp 1688980957
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_475
timestamp 1688980957
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_477
timestamp 1688980957
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_489
timestamp 1688980957
transform 1 0 46092 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_501
timestamp 1688980957
transform 1 0 47196 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_513
timestamp 1688980957
transform 1 0 48300 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_525
timestamp 1688980957
transform 1 0 49404 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_531
timestamp 1688980957
transform 1 0 49956 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_533
timestamp 1688980957
transform 1 0 50140 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_545
timestamp 1688980957
transform 1 0 51244 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_557
timestamp 1688980957
transform 1 0 52348 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_569
timestamp 1688980957
transform 1 0 53452 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_581
timestamp 1688980957
transform 1 0 54556 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_587
timestamp 1688980957
transform 1 0 55108 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_589
timestamp 1688980957
transform 1 0 55292 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_595
timestamp 1688980957
transform 1 0 55844 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_607
timestamp 1688980957
transform 1 0 56948 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_618
timestamp 1688980957
transform 1 0 57960 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_15
timestamp 1688980957
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_27
timestamp 1688980957
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_39
timestamp 1688980957
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_51
timestamp 1688980957
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_55
timestamp 1688980957
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_69
timestamp 1688980957
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_81
timestamp 1688980957
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_93
timestamp 1688980957
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_105
timestamp 1688980957
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_111
timestamp 1688980957
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 1688980957
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 1688980957
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_161
timestamp 1688980957
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 1688980957
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_169
timestamp 1688980957
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_181
timestamp 1688980957
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_193
timestamp 1688980957
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_205
timestamp 1688980957
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_217
timestamp 1688980957
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_223
timestamp 1688980957
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_225
timestamp 1688980957
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_237
timestamp 1688980957
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_249
timestamp 1688980957
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_261
timestamp 1688980957
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_273
timestamp 1688980957
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_279
timestamp 1688980957
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_281
timestamp 1688980957
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_293
timestamp 1688980957
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_305
timestamp 1688980957
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_317
timestamp 1688980957
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_329
timestamp 1688980957
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_335
timestamp 1688980957
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_337
timestamp 1688980957
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_349
timestamp 1688980957
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_361
timestamp 1688980957
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_373
timestamp 1688980957
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_385
timestamp 1688980957
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_391
timestamp 1688980957
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_393
timestamp 1688980957
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_405
timestamp 1688980957
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_417
timestamp 1688980957
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_429
timestamp 1688980957
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_441
timestamp 1688980957
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_447
timestamp 1688980957
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_449
timestamp 1688980957
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_461
timestamp 1688980957
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_473
timestamp 1688980957
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_485
timestamp 1688980957
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_497
timestamp 1688980957
transform 1 0 46828 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_503
timestamp 1688980957
transform 1 0 47380 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_505
timestamp 1688980957
transform 1 0 47564 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_517
timestamp 1688980957
transform 1 0 48668 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_529
timestamp 1688980957
transform 1 0 49772 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_541
timestamp 1688980957
transform 1 0 50876 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_553
timestamp 1688980957
transform 1 0 51980 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_559
timestamp 1688980957
transform 1 0 52532 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_561
timestamp 1688980957
transform 1 0 52716 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_573
timestamp 1688980957
transform 1 0 53820 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_585
timestamp 1688980957
transform 1 0 54924 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_597
timestamp 1688980957
transform 1 0 56028 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_601
timestamp 1688980957
transform 1 0 56396 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_614
timestamp 1688980957
transform 1 0 57592 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_623
timestamp 1688980957
transform 1 0 58420 0 -1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_3
timestamp 1688980957
transform 1 0 1380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_15
timestamp 1688980957
transform 1 0 2484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_27
timestamp 1688980957
transform 1 0 3588 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_41
timestamp 1688980957
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_53
timestamp 1688980957
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_65
timestamp 1688980957
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_77
timestamp 1688980957
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_83
timestamp 1688980957
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_85
timestamp 1688980957
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_97
timestamp 1688980957
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_109
timestamp 1688980957
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_121
timestamp 1688980957
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_133
timestamp 1688980957
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 1688980957
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_141
timestamp 1688980957
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_153
timestamp 1688980957
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_165
timestamp 1688980957
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_177
timestamp 1688980957
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_189
timestamp 1688980957
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_195
timestamp 1688980957
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_197
timestamp 1688980957
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_209
timestamp 1688980957
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_221
timestamp 1688980957
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_233
timestamp 1688980957
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_245
timestamp 1688980957
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_251
timestamp 1688980957
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_253
timestamp 1688980957
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_265
timestamp 1688980957
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_277
timestamp 1688980957
transform 1 0 26588 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_289
timestamp 1688980957
transform 1 0 27692 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_301
timestamp 1688980957
transform 1 0 28796 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_307
timestamp 1688980957
transform 1 0 29348 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_309
timestamp 1688980957
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_321
timestamp 1688980957
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_333
timestamp 1688980957
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_345
timestamp 1688980957
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_357
timestamp 1688980957
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_363
timestamp 1688980957
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_365
timestamp 1688980957
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_377
timestamp 1688980957
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_389
timestamp 1688980957
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_401
timestamp 1688980957
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_413
timestamp 1688980957
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_419
timestamp 1688980957
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_421
timestamp 1688980957
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_433
timestamp 1688980957
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_445
timestamp 1688980957
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_457
timestamp 1688980957
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_469
timestamp 1688980957
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_475
timestamp 1688980957
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_477
timestamp 1688980957
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_489
timestamp 1688980957
transform 1 0 46092 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_501
timestamp 1688980957
transform 1 0 47196 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_513
timestamp 1688980957
transform 1 0 48300 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_525
timestamp 1688980957
transform 1 0 49404 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_531
timestamp 1688980957
transform 1 0 49956 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_533
timestamp 1688980957
transform 1 0 50140 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_545
timestamp 1688980957
transform 1 0 51244 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_557
timestamp 1688980957
transform 1 0 52348 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_569
timestamp 1688980957
transform 1 0 53452 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_581
timestamp 1688980957
transform 1 0 54556 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_587
timestamp 1688980957
transform 1 0 55108 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_589
timestamp 1688980957
transform 1 0 55292 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_76_601
timestamp 1688980957
transform 1 0 56396 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_613
timestamp 1688980957
transform 1 0 57500 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_623
timestamp 1688980957
transform 1 0 58420 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_19
timestamp 1688980957
transform 1 0 2852 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_31
timestamp 1688980957
transform 1 0 3956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_43
timestamp 1688980957
transform 1 0 5060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1688980957
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_57
timestamp 1688980957
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_69
timestamp 1688980957
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_81
timestamp 1688980957
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_93
timestamp 1688980957
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_105
timestamp 1688980957
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 1688980957
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_113
timestamp 1688980957
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_125
timestamp 1688980957
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_137
timestamp 1688980957
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_149
timestamp 1688980957
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_161
timestamp 1688980957
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_167
timestamp 1688980957
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_169
timestamp 1688980957
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_181
timestamp 1688980957
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_193
timestamp 1688980957
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_205
timestamp 1688980957
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_217
timestamp 1688980957
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_223
timestamp 1688980957
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_225
timestamp 1688980957
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_237
timestamp 1688980957
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_249
timestamp 1688980957
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_261
timestamp 1688980957
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_273
timestamp 1688980957
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_279
timestamp 1688980957
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_281
timestamp 1688980957
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_293
timestamp 1688980957
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_305
timestamp 1688980957
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_317
timestamp 1688980957
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_329
timestamp 1688980957
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_335
timestamp 1688980957
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_337
timestamp 1688980957
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_349
timestamp 1688980957
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_361
timestamp 1688980957
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_373
timestamp 1688980957
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_385
timestamp 1688980957
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_391
timestamp 1688980957
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_393
timestamp 1688980957
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_405
timestamp 1688980957
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_417
timestamp 1688980957
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_429
timestamp 1688980957
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_441
timestamp 1688980957
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_447
timestamp 1688980957
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_449
timestamp 1688980957
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_461
timestamp 1688980957
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_473
timestamp 1688980957
transform 1 0 44620 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_485
timestamp 1688980957
transform 1 0 45724 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_497
timestamp 1688980957
transform 1 0 46828 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_503
timestamp 1688980957
transform 1 0 47380 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_505
timestamp 1688980957
transform 1 0 47564 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_517
timestamp 1688980957
transform 1 0 48668 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_529
timestamp 1688980957
transform 1 0 49772 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_541
timestamp 1688980957
transform 1 0 50876 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_553
timestamp 1688980957
transform 1 0 51980 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_559
timestamp 1688980957
transform 1 0 52532 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_561
timestamp 1688980957
transform 1 0 52716 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_573
timestamp 1688980957
transform 1 0 53820 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_585
timestamp 1688980957
transform 1 0 54924 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_77_597
timestamp 1688980957
transform 1 0 56028 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77_609
timestamp 1688980957
transform 1 0 57132 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_615
timestamp 1688980957
transform 1 0 57684 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_617
timestamp 1688980957
transform 1 0 57868 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_621
timestamp 1688980957
transform 1 0 58236 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_3
timestamp 1688980957
transform 1 0 1380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_15
timestamp 1688980957
transform 1 0 2484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_27
timestamp 1688980957
transform 1 0 3588 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_29
timestamp 1688980957
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_41
timestamp 1688980957
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_53
timestamp 1688980957
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_65
timestamp 1688980957
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_77
timestamp 1688980957
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_83
timestamp 1688980957
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_85
timestamp 1688980957
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_97
timestamp 1688980957
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_109
timestamp 1688980957
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_121
timestamp 1688980957
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_133
timestamp 1688980957
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_139
timestamp 1688980957
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_141
timestamp 1688980957
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_153
timestamp 1688980957
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_165
timestamp 1688980957
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_177
timestamp 1688980957
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_189
timestamp 1688980957
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_195
timestamp 1688980957
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_197
timestamp 1688980957
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_209
timestamp 1688980957
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_221
timestamp 1688980957
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_233
timestamp 1688980957
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_245
timestamp 1688980957
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_251
timestamp 1688980957
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_253
timestamp 1688980957
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_265
timestamp 1688980957
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_277
timestamp 1688980957
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_289
timestamp 1688980957
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_301
timestamp 1688980957
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_307
timestamp 1688980957
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_309
timestamp 1688980957
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_321
timestamp 1688980957
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_333
timestamp 1688980957
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_345
timestamp 1688980957
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_357
timestamp 1688980957
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_363
timestamp 1688980957
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_365
timestamp 1688980957
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_377
timestamp 1688980957
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_389
timestamp 1688980957
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_401
timestamp 1688980957
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_413
timestamp 1688980957
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_419
timestamp 1688980957
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_421
timestamp 1688980957
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_433
timestamp 1688980957
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_445
timestamp 1688980957
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_457
timestamp 1688980957
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_469
timestamp 1688980957
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_475
timestamp 1688980957
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_477
timestamp 1688980957
transform 1 0 44988 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_489
timestamp 1688980957
transform 1 0 46092 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_501
timestamp 1688980957
transform 1 0 47196 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_513
timestamp 1688980957
transform 1 0 48300 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_525
timestamp 1688980957
transform 1 0 49404 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_531
timestamp 1688980957
transform 1 0 49956 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_533
timestamp 1688980957
transform 1 0 50140 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_545
timestamp 1688980957
transform 1 0 51244 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_557
timestamp 1688980957
transform 1 0 52348 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_569
timestamp 1688980957
transform 1 0 53452 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78_581
timestamp 1688980957
transform 1 0 54556 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_587
timestamp 1688980957
transform 1 0 55108 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_589
timestamp 1688980957
transform 1 0 55292 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_78_601
timestamp 1688980957
transform 1 0 56396 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_78_613
timestamp 1688980957
transform 1 0 57500 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78_621
timestamp 1688980957
transform 1 0 58236 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_3
timestamp 1688980957
transform 1 0 1380 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_15
timestamp 1688980957
transform 1 0 2484 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_27
timestamp 1688980957
transform 1 0 3588 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_39
timestamp 1688980957
transform 1 0 4692 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_79_51
timestamp 1688980957
transform 1 0 5796 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_55
timestamp 1688980957
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_57
timestamp 1688980957
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_69
timestamp 1688980957
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_81
timestamp 1688980957
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_93
timestamp 1688980957
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_105
timestamp 1688980957
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_111
timestamp 1688980957
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_113
timestamp 1688980957
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_125
timestamp 1688980957
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_137
timestamp 1688980957
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_149
timestamp 1688980957
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_161
timestamp 1688980957
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_167
timestamp 1688980957
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_169
timestamp 1688980957
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_181
timestamp 1688980957
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_193
timestamp 1688980957
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_205
timestamp 1688980957
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_217
timestamp 1688980957
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_223
timestamp 1688980957
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_225
timestamp 1688980957
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_237
timestamp 1688980957
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_249
timestamp 1688980957
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_261
timestamp 1688980957
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_273
timestamp 1688980957
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_279
timestamp 1688980957
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_281
timestamp 1688980957
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_293
timestamp 1688980957
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_305
timestamp 1688980957
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_317
timestamp 1688980957
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_329
timestamp 1688980957
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_335
timestamp 1688980957
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_337
timestamp 1688980957
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_349
timestamp 1688980957
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_361
timestamp 1688980957
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_373
timestamp 1688980957
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_385
timestamp 1688980957
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_391
timestamp 1688980957
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_393
timestamp 1688980957
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_405
timestamp 1688980957
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_417
timestamp 1688980957
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_429
timestamp 1688980957
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_441
timestamp 1688980957
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_447
timestamp 1688980957
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_449
timestamp 1688980957
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_461
timestamp 1688980957
transform 1 0 43516 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_473
timestamp 1688980957
transform 1 0 44620 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_485
timestamp 1688980957
transform 1 0 45724 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_497
timestamp 1688980957
transform 1 0 46828 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_503
timestamp 1688980957
transform 1 0 47380 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_505
timestamp 1688980957
transform 1 0 47564 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_517
timestamp 1688980957
transform 1 0 48668 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_529
timestamp 1688980957
transform 1 0 49772 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_541
timestamp 1688980957
transform 1 0 50876 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_553
timestamp 1688980957
transform 1 0 51980 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_559
timestamp 1688980957
transform 1 0 52532 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_561
timestamp 1688980957
transform 1 0 52716 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_573
timestamp 1688980957
transform 1 0 53820 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_585
timestamp 1688980957
transform 1 0 54924 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_79_597
timestamp 1688980957
transform 1 0 56028 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_79_609
timestamp 1688980957
transform 1 0 57132 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79_615
timestamp 1688980957
transform 1 0 57684 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_79_617
timestamp 1688980957
transform 1 0 57868 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_19
timestamp 1688980957
transform 1 0 2852 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_27
timestamp 1688980957
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_29
timestamp 1688980957
transform 1 0 3772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_41
timestamp 1688980957
transform 1 0 4876 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_53
timestamp 1688980957
transform 1 0 5980 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_65
timestamp 1688980957
transform 1 0 7084 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_77
timestamp 1688980957
transform 1 0 8188 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_83
timestamp 1688980957
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_85
timestamp 1688980957
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_97
timestamp 1688980957
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_109
timestamp 1688980957
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_121
timestamp 1688980957
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_133
timestamp 1688980957
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_139
timestamp 1688980957
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_141
timestamp 1688980957
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_153
timestamp 1688980957
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_165
timestamp 1688980957
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_177
timestamp 1688980957
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_189
timestamp 1688980957
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_195
timestamp 1688980957
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_197
timestamp 1688980957
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_209
timestamp 1688980957
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_221
timestamp 1688980957
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_233
timestamp 1688980957
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_245
timestamp 1688980957
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_251
timestamp 1688980957
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_253
timestamp 1688980957
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_265
timestamp 1688980957
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_277
timestamp 1688980957
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_289
timestamp 1688980957
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_301
timestamp 1688980957
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_307
timestamp 1688980957
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_309
timestamp 1688980957
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_321
timestamp 1688980957
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_333
timestamp 1688980957
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_345
timestamp 1688980957
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_357
timestamp 1688980957
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_363
timestamp 1688980957
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_365
timestamp 1688980957
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_377
timestamp 1688980957
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_389
timestamp 1688980957
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_401
timestamp 1688980957
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_413
timestamp 1688980957
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_419
timestamp 1688980957
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_421
timestamp 1688980957
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_433
timestamp 1688980957
transform 1 0 40940 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_445
timestamp 1688980957
transform 1 0 42044 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_457
timestamp 1688980957
transform 1 0 43148 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_469
timestamp 1688980957
transform 1 0 44252 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_475
timestamp 1688980957
transform 1 0 44804 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_477
timestamp 1688980957
transform 1 0 44988 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_489
timestamp 1688980957
transform 1 0 46092 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_501
timestamp 1688980957
transform 1 0 47196 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_513
timestamp 1688980957
transform 1 0 48300 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_525
timestamp 1688980957
transform 1 0 49404 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_531
timestamp 1688980957
transform 1 0 49956 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_533
timestamp 1688980957
transform 1 0 50140 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_545
timestamp 1688980957
transform 1 0 51244 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_557
timestamp 1688980957
transform 1 0 52348 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_569
timestamp 1688980957
transform 1 0 53452 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_80_581
timestamp 1688980957
transform 1 0 54556 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_587
timestamp 1688980957
transform 1 0 55108 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_589
timestamp 1688980957
transform 1 0 55292 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_80_601
timestamp 1688980957
transform 1 0 56396 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_80_613
timestamp 1688980957
transform 1 0 57500 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80_621
timestamp 1688980957
transform 1 0 58236 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_3
timestamp 1688980957
transform 1 0 1380 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_15
timestamp 1688980957
transform 1 0 2484 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_27
timestamp 1688980957
transform 1 0 3588 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_39
timestamp 1688980957
transform 1 0 4692 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_51
timestamp 1688980957
transform 1 0 5796 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_55
timestamp 1688980957
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_57
timestamp 1688980957
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_69
timestamp 1688980957
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_81
timestamp 1688980957
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_93
timestamp 1688980957
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_105
timestamp 1688980957
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_111
timestamp 1688980957
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_113
timestamp 1688980957
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_125
timestamp 1688980957
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_137
timestamp 1688980957
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_149
timestamp 1688980957
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_161
timestamp 1688980957
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_167
timestamp 1688980957
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_169
timestamp 1688980957
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_181
timestamp 1688980957
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_193
timestamp 1688980957
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_205
timestamp 1688980957
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_217
timestamp 1688980957
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_223
timestamp 1688980957
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_225
timestamp 1688980957
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_237
timestamp 1688980957
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_249
timestamp 1688980957
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_261
timestamp 1688980957
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_273
timestamp 1688980957
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_279
timestamp 1688980957
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_281
timestamp 1688980957
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_293
timestamp 1688980957
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_305
timestamp 1688980957
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_317
timestamp 1688980957
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_329
timestamp 1688980957
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_335
timestamp 1688980957
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_337
timestamp 1688980957
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_349
timestamp 1688980957
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_361
timestamp 1688980957
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_373
timestamp 1688980957
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_385
timestamp 1688980957
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_391
timestamp 1688980957
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_393
timestamp 1688980957
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_405
timestamp 1688980957
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_417
timestamp 1688980957
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_429
timestamp 1688980957
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_441
timestamp 1688980957
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_447
timestamp 1688980957
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_449
timestamp 1688980957
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_461
timestamp 1688980957
transform 1 0 43516 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_473
timestamp 1688980957
transform 1 0 44620 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_485
timestamp 1688980957
transform 1 0 45724 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_497
timestamp 1688980957
transform 1 0 46828 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_503
timestamp 1688980957
transform 1 0 47380 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_505
timestamp 1688980957
transform 1 0 47564 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_517
timestamp 1688980957
transform 1 0 48668 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_529
timestamp 1688980957
transform 1 0 49772 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_541
timestamp 1688980957
transform 1 0 50876 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_553
timestamp 1688980957
transform 1 0 51980 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_559
timestamp 1688980957
transform 1 0 52532 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_561
timestamp 1688980957
transform 1 0 52716 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_573
timestamp 1688980957
transform 1 0 53820 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_585
timestamp 1688980957
transform 1 0 54924 0 -1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_81_597
timestamp 1688980957
transform 1 0 56028 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_81_609
timestamp 1688980957
transform 1 0 57132 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_615
timestamp 1688980957
transform 1 0 57684 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_81_617
timestamp 1688980957
transform 1 0 57868 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_81_621
timestamp 1688980957
transform 1 0 58236 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_3
timestamp 1688980957
transform 1 0 1380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_15
timestamp 1688980957
transform 1 0 2484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_27
timestamp 1688980957
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_29
timestamp 1688980957
transform 1 0 3772 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_41
timestamp 1688980957
transform 1 0 4876 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_53
timestamp 1688980957
transform 1 0 5980 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_65
timestamp 1688980957
transform 1 0 7084 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_77
timestamp 1688980957
transform 1 0 8188 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_83
timestamp 1688980957
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_85
timestamp 1688980957
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_97
timestamp 1688980957
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_109
timestamp 1688980957
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_121
timestamp 1688980957
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_133
timestamp 1688980957
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_139
timestamp 1688980957
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_141
timestamp 1688980957
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_153
timestamp 1688980957
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_165
timestamp 1688980957
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_177
timestamp 1688980957
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_189
timestamp 1688980957
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_195
timestamp 1688980957
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_197
timestamp 1688980957
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_209
timestamp 1688980957
transform 1 0 20332 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_221
timestamp 1688980957
transform 1 0 21436 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_233
timestamp 1688980957
transform 1 0 22540 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_245
timestamp 1688980957
transform 1 0 23644 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_251
timestamp 1688980957
transform 1 0 24196 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_253
timestamp 1688980957
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_265
timestamp 1688980957
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_277
timestamp 1688980957
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_289
timestamp 1688980957
transform 1 0 27692 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_301
timestamp 1688980957
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_307
timestamp 1688980957
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_309
timestamp 1688980957
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_321
timestamp 1688980957
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_333
timestamp 1688980957
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_345
timestamp 1688980957
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_357
timestamp 1688980957
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_363
timestamp 1688980957
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_365
timestamp 1688980957
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_377
timestamp 1688980957
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_389
timestamp 1688980957
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_401
timestamp 1688980957
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_413
timestamp 1688980957
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_419
timestamp 1688980957
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_421
timestamp 1688980957
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_433
timestamp 1688980957
transform 1 0 40940 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_445
timestamp 1688980957
transform 1 0 42044 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_457
timestamp 1688980957
transform 1 0 43148 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_469
timestamp 1688980957
transform 1 0 44252 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_475
timestamp 1688980957
transform 1 0 44804 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_477
timestamp 1688980957
transform 1 0 44988 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_489
timestamp 1688980957
transform 1 0 46092 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_501
timestamp 1688980957
transform 1 0 47196 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_513
timestamp 1688980957
transform 1 0 48300 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_525
timestamp 1688980957
transform 1 0 49404 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_531
timestamp 1688980957
transform 1 0 49956 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_533
timestamp 1688980957
transform 1 0 50140 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_545
timestamp 1688980957
transform 1 0 51244 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_557
timestamp 1688980957
transform 1 0 52348 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_569
timestamp 1688980957
transform 1 0 53452 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_82_581
timestamp 1688980957
transform 1 0 54556 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_82_587
timestamp 1688980957
transform 1 0 55108 0 1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_589
timestamp 1688980957
transform 1 0 55292 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_601
timestamp 1688980957
transform 1 0 56396 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_82_613
timestamp 1688980957
transform 1 0 57500 0 1 46784
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_19
timestamp 1688980957
transform 1 0 2852 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_31
timestamp 1688980957
transform 1 0 3956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_43
timestamp 1688980957
transform 1 0 5060 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_55
timestamp 1688980957
transform 1 0 6164 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_57
timestamp 1688980957
transform 1 0 6348 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_69
timestamp 1688980957
transform 1 0 7452 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_81
timestamp 1688980957
transform 1 0 8556 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_93
timestamp 1688980957
transform 1 0 9660 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_105
timestamp 1688980957
transform 1 0 10764 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_111
timestamp 1688980957
transform 1 0 11316 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_113
timestamp 1688980957
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_125
timestamp 1688980957
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_137
timestamp 1688980957
transform 1 0 13708 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_149
timestamp 1688980957
transform 1 0 14812 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_161
timestamp 1688980957
transform 1 0 15916 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_167
timestamp 1688980957
transform 1 0 16468 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_169
timestamp 1688980957
transform 1 0 16652 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_181
timestamp 1688980957
transform 1 0 17756 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_193
timestamp 1688980957
transform 1 0 18860 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_205
timestamp 1688980957
transform 1 0 19964 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_217
timestamp 1688980957
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_223
timestamp 1688980957
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_225
timestamp 1688980957
transform 1 0 21804 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_237
timestamp 1688980957
transform 1 0 22908 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_249
timestamp 1688980957
transform 1 0 24012 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_261
timestamp 1688980957
transform 1 0 25116 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_273
timestamp 1688980957
transform 1 0 26220 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_279
timestamp 1688980957
transform 1 0 26772 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_281
timestamp 1688980957
transform 1 0 26956 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_293
timestamp 1688980957
transform 1 0 28060 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_305
timestamp 1688980957
transform 1 0 29164 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_317
timestamp 1688980957
transform 1 0 30268 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_329
timestamp 1688980957
transform 1 0 31372 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_335
timestamp 1688980957
transform 1 0 31924 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_337
timestamp 1688980957
transform 1 0 32108 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_349
timestamp 1688980957
transform 1 0 33212 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_361
timestamp 1688980957
transform 1 0 34316 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_373
timestamp 1688980957
transform 1 0 35420 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_385
timestamp 1688980957
transform 1 0 36524 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_391
timestamp 1688980957
transform 1 0 37076 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_393
timestamp 1688980957
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_405
timestamp 1688980957
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_417
timestamp 1688980957
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_429
timestamp 1688980957
transform 1 0 40572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_441
timestamp 1688980957
transform 1 0 41676 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_447
timestamp 1688980957
transform 1 0 42228 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_449
timestamp 1688980957
transform 1 0 42412 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_461
timestamp 1688980957
transform 1 0 43516 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_473
timestamp 1688980957
transform 1 0 44620 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_485
timestamp 1688980957
transform 1 0 45724 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_497
timestamp 1688980957
transform 1 0 46828 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_503
timestamp 1688980957
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_505
timestamp 1688980957
transform 1 0 47564 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_517
timestamp 1688980957
transform 1 0 48668 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_529
timestamp 1688980957
transform 1 0 49772 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_541
timestamp 1688980957
transform 1 0 50876 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_553
timestamp 1688980957
transform 1 0 51980 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_559
timestamp 1688980957
transform 1 0 52532 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_561
timestamp 1688980957
transform 1 0 52716 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_573
timestamp 1688980957
transform 1 0 53820 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_585
timestamp 1688980957
transform 1 0 54924 0 -1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_83_597
timestamp 1688980957
transform 1 0 56028 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_83_609
timestamp 1688980957
transform 1 0 57132 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_615
timestamp 1688980957
transform 1 0 57684 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_83_617
timestamp 1688980957
transform 1 0 57868 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83_621
timestamp 1688980957
transform 1 0 58236 0 -1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_3
timestamp 1688980957
transform 1 0 1380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_15
timestamp 1688980957
transform 1 0 2484 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_27
timestamp 1688980957
transform 1 0 3588 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_29
timestamp 1688980957
transform 1 0 3772 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_41
timestamp 1688980957
transform 1 0 4876 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_53
timestamp 1688980957
transform 1 0 5980 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_65
timestamp 1688980957
transform 1 0 7084 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_77
timestamp 1688980957
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_83
timestamp 1688980957
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_85
timestamp 1688980957
transform 1 0 8924 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_97
timestamp 1688980957
transform 1 0 10028 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_109
timestamp 1688980957
transform 1 0 11132 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_121
timestamp 1688980957
transform 1 0 12236 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_133
timestamp 1688980957
transform 1 0 13340 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_139
timestamp 1688980957
transform 1 0 13892 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_141
timestamp 1688980957
transform 1 0 14076 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_153
timestamp 1688980957
transform 1 0 15180 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_165
timestamp 1688980957
transform 1 0 16284 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_177
timestamp 1688980957
transform 1 0 17388 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_189
timestamp 1688980957
transform 1 0 18492 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_195
timestamp 1688980957
transform 1 0 19044 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_197
timestamp 1688980957
transform 1 0 19228 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_209
timestamp 1688980957
transform 1 0 20332 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_221
timestamp 1688980957
transform 1 0 21436 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_233
timestamp 1688980957
transform 1 0 22540 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_245
timestamp 1688980957
transform 1 0 23644 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_251
timestamp 1688980957
transform 1 0 24196 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_253
timestamp 1688980957
transform 1 0 24380 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_265
timestamp 1688980957
transform 1 0 25484 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_277
timestamp 1688980957
transform 1 0 26588 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_289
timestamp 1688980957
transform 1 0 27692 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_301
timestamp 1688980957
transform 1 0 28796 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_307
timestamp 1688980957
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_309
timestamp 1688980957
transform 1 0 29532 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_321
timestamp 1688980957
transform 1 0 30636 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_333
timestamp 1688980957
transform 1 0 31740 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_345
timestamp 1688980957
transform 1 0 32844 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_357
timestamp 1688980957
transform 1 0 33948 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_363
timestamp 1688980957
transform 1 0 34500 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_365
timestamp 1688980957
transform 1 0 34684 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_377
timestamp 1688980957
transform 1 0 35788 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_389
timestamp 1688980957
transform 1 0 36892 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_401
timestamp 1688980957
transform 1 0 37996 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_413
timestamp 1688980957
transform 1 0 39100 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_419
timestamp 1688980957
transform 1 0 39652 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_421
timestamp 1688980957
transform 1 0 39836 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_433
timestamp 1688980957
transform 1 0 40940 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_445
timestamp 1688980957
transform 1 0 42044 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_457
timestamp 1688980957
transform 1 0 43148 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_469
timestamp 1688980957
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_475
timestamp 1688980957
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_477
timestamp 1688980957
transform 1 0 44988 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_489
timestamp 1688980957
transform 1 0 46092 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_501
timestamp 1688980957
transform 1 0 47196 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_513
timestamp 1688980957
transform 1 0 48300 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_525
timestamp 1688980957
transform 1 0 49404 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_531
timestamp 1688980957
transform 1 0 49956 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_533
timestamp 1688980957
transform 1 0 50140 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_545
timestamp 1688980957
transform 1 0 51244 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_557
timestamp 1688980957
transform 1 0 52348 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_569
timestamp 1688980957
transform 1 0 53452 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_84_581
timestamp 1688980957
transform 1 0 54556 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_587
timestamp 1688980957
transform 1 0 55108 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_589
timestamp 1688980957
transform 1 0 55292 0 1 47872
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_84_601
timestamp 1688980957
transform 1 0 56396 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_84_613
timestamp 1688980957
transform 1 0 57500 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_84_621
timestamp 1688980957
transform 1 0 58236 0 1 47872
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_3
timestamp 1688980957
transform 1 0 1380 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_15
timestamp 1688980957
transform 1 0 2484 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_27
timestamp 1688980957
transform 1 0 3588 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_39
timestamp 1688980957
transform 1 0 4692 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_85_51
timestamp 1688980957
transform 1 0 5796 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_55
timestamp 1688980957
transform 1 0 6164 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_57
timestamp 1688980957
transform 1 0 6348 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_69
timestamp 1688980957
transform 1 0 7452 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_81
timestamp 1688980957
transform 1 0 8556 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_93
timestamp 1688980957
transform 1 0 9660 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_105
timestamp 1688980957
transform 1 0 10764 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_111
timestamp 1688980957
transform 1 0 11316 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_113
timestamp 1688980957
transform 1 0 11500 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_125
timestamp 1688980957
transform 1 0 12604 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_137
timestamp 1688980957
transform 1 0 13708 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_149
timestamp 1688980957
transform 1 0 14812 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_161
timestamp 1688980957
transform 1 0 15916 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_167
timestamp 1688980957
transform 1 0 16468 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_169
timestamp 1688980957
transform 1 0 16652 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_181
timestamp 1688980957
transform 1 0 17756 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_193
timestamp 1688980957
transform 1 0 18860 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_205
timestamp 1688980957
transform 1 0 19964 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_217
timestamp 1688980957
transform 1 0 21068 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_223
timestamp 1688980957
transform 1 0 21620 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_225
timestamp 1688980957
transform 1 0 21804 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_237
timestamp 1688980957
transform 1 0 22908 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_249
timestamp 1688980957
transform 1 0 24012 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_261
timestamp 1688980957
transform 1 0 25116 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_273
timestamp 1688980957
transform 1 0 26220 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_279
timestamp 1688980957
transform 1 0 26772 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_281
timestamp 1688980957
transform 1 0 26956 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_293
timestamp 1688980957
transform 1 0 28060 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_305
timestamp 1688980957
transform 1 0 29164 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_317
timestamp 1688980957
transform 1 0 30268 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_329
timestamp 1688980957
transform 1 0 31372 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_335
timestamp 1688980957
transform 1 0 31924 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_337
timestamp 1688980957
transform 1 0 32108 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_349
timestamp 1688980957
transform 1 0 33212 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_361
timestamp 1688980957
transform 1 0 34316 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_373
timestamp 1688980957
transform 1 0 35420 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_385
timestamp 1688980957
transform 1 0 36524 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_391
timestamp 1688980957
transform 1 0 37076 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_393
timestamp 1688980957
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_405
timestamp 1688980957
transform 1 0 38364 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_417
timestamp 1688980957
transform 1 0 39468 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_429
timestamp 1688980957
transform 1 0 40572 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_441
timestamp 1688980957
transform 1 0 41676 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_447
timestamp 1688980957
transform 1 0 42228 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_449
timestamp 1688980957
transform 1 0 42412 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_461
timestamp 1688980957
transform 1 0 43516 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_473
timestamp 1688980957
transform 1 0 44620 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_485
timestamp 1688980957
transform 1 0 45724 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_497
timestamp 1688980957
transform 1 0 46828 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_503
timestamp 1688980957
transform 1 0 47380 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_505
timestamp 1688980957
transform 1 0 47564 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_517
timestamp 1688980957
transform 1 0 48668 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_529
timestamp 1688980957
transform 1 0 49772 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_541
timestamp 1688980957
transform 1 0 50876 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_553
timestamp 1688980957
transform 1 0 51980 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_559
timestamp 1688980957
transform 1 0 52532 0 -1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_561
timestamp 1688980957
transform 1 0 52716 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_573
timestamp 1688980957
transform 1 0 53820 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_585
timestamp 1688980957
transform 1 0 54924 0 -1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85_597
timestamp 1688980957
transform 1 0 56028 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85_609
timestamp 1688980957
transform 1 0 57132 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85_615
timestamp 1688980957
transform 1 0 57684 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85_617
timestamp 1688980957
transform 1 0 57868 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_19
timestamp 1688980957
transform 1 0 2852 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_27
timestamp 1688980957
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_29
timestamp 1688980957
transform 1 0 3772 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_41
timestamp 1688980957
transform 1 0 4876 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_53
timestamp 1688980957
transform 1 0 5980 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_65
timestamp 1688980957
transform 1 0 7084 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_77
timestamp 1688980957
transform 1 0 8188 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_83
timestamp 1688980957
transform 1 0 8740 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_85
timestamp 1688980957
transform 1 0 8924 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_97
timestamp 1688980957
transform 1 0 10028 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_109
timestamp 1688980957
transform 1 0 11132 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_121
timestamp 1688980957
transform 1 0 12236 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_133
timestamp 1688980957
transform 1 0 13340 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_139
timestamp 1688980957
transform 1 0 13892 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_141
timestamp 1688980957
transform 1 0 14076 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_153
timestamp 1688980957
transform 1 0 15180 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_165
timestamp 1688980957
transform 1 0 16284 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_177
timestamp 1688980957
transform 1 0 17388 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_189
timestamp 1688980957
transform 1 0 18492 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_195
timestamp 1688980957
transform 1 0 19044 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_197
timestamp 1688980957
transform 1 0 19228 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_209
timestamp 1688980957
transform 1 0 20332 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_221
timestamp 1688980957
transform 1 0 21436 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_233
timestamp 1688980957
transform 1 0 22540 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_245
timestamp 1688980957
transform 1 0 23644 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_251
timestamp 1688980957
transform 1 0 24196 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_253
timestamp 1688980957
transform 1 0 24380 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_265
timestamp 1688980957
transform 1 0 25484 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_277
timestamp 1688980957
transform 1 0 26588 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_289
timestamp 1688980957
transform 1 0 27692 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_301
timestamp 1688980957
transform 1 0 28796 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_307
timestamp 1688980957
transform 1 0 29348 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_309
timestamp 1688980957
transform 1 0 29532 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_321
timestamp 1688980957
transform 1 0 30636 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_333
timestamp 1688980957
transform 1 0 31740 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_345
timestamp 1688980957
transform 1 0 32844 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_357
timestamp 1688980957
transform 1 0 33948 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_363
timestamp 1688980957
transform 1 0 34500 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_365
timestamp 1688980957
transform 1 0 34684 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_377
timestamp 1688980957
transform 1 0 35788 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_389
timestamp 1688980957
transform 1 0 36892 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_401
timestamp 1688980957
transform 1 0 37996 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_413
timestamp 1688980957
transform 1 0 39100 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_419
timestamp 1688980957
transform 1 0 39652 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_421
timestamp 1688980957
transform 1 0 39836 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_433
timestamp 1688980957
transform 1 0 40940 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_445
timestamp 1688980957
transform 1 0 42044 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_457
timestamp 1688980957
transform 1 0 43148 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_469
timestamp 1688980957
transform 1 0 44252 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_475
timestamp 1688980957
transform 1 0 44804 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_477
timestamp 1688980957
transform 1 0 44988 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_489
timestamp 1688980957
transform 1 0 46092 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_501
timestamp 1688980957
transform 1 0 47196 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_513
timestamp 1688980957
transform 1 0 48300 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_525
timestamp 1688980957
transform 1 0 49404 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_531
timestamp 1688980957
transform 1 0 49956 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_533
timestamp 1688980957
transform 1 0 50140 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_545
timestamp 1688980957
transform 1 0 51244 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_557
timestamp 1688980957
transform 1 0 52348 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_569
timestamp 1688980957
transform 1 0 53452 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86_581
timestamp 1688980957
transform 1 0 54556 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_587
timestamp 1688980957
transform 1 0 55108 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_589
timestamp 1688980957
transform 1 0 55292 0 1 48960
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_86_601
timestamp 1688980957
transform 1 0 56396 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_86_613
timestamp 1688980957
transform 1 0 57500 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_86_621
timestamp 1688980957
transform 1 0 58236 0 1 48960
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_3
timestamp 1688980957
transform 1 0 1380 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_15
timestamp 1688980957
transform 1 0 2484 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_27
timestamp 1688980957
transform 1 0 3588 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_39
timestamp 1688980957
transform 1 0 4692 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_51
timestamp 1688980957
transform 1 0 5796 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_55
timestamp 1688980957
transform 1 0 6164 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_57
timestamp 1688980957
transform 1 0 6348 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_69
timestamp 1688980957
transform 1 0 7452 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_81
timestamp 1688980957
transform 1 0 8556 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_93
timestamp 1688980957
transform 1 0 9660 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_105
timestamp 1688980957
transform 1 0 10764 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_111
timestamp 1688980957
transform 1 0 11316 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_113
timestamp 1688980957
transform 1 0 11500 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_125
timestamp 1688980957
transform 1 0 12604 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_137
timestamp 1688980957
transform 1 0 13708 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_149
timestamp 1688980957
transform 1 0 14812 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_161
timestamp 1688980957
transform 1 0 15916 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_167
timestamp 1688980957
transform 1 0 16468 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_169
timestamp 1688980957
transform 1 0 16652 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_181
timestamp 1688980957
transform 1 0 17756 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_193
timestamp 1688980957
transform 1 0 18860 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_205
timestamp 1688980957
transform 1 0 19964 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_217
timestamp 1688980957
transform 1 0 21068 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_223
timestamp 1688980957
transform 1 0 21620 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_225
timestamp 1688980957
transform 1 0 21804 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_237
timestamp 1688980957
transform 1 0 22908 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_249
timestamp 1688980957
transform 1 0 24012 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_261
timestamp 1688980957
transform 1 0 25116 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_273
timestamp 1688980957
transform 1 0 26220 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_279
timestamp 1688980957
transform 1 0 26772 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_281
timestamp 1688980957
transform 1 0 26956 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_293
timestamp 1688980957
transform 1 0 28060 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_305
timestamp 1688980957
transform 1 0 29164 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_317
timestamp 1688980957
transform 1 0 30268 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_329
timestamp 1688980957
transform 1 0 31372 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_335
timestamp 1688980957
transform 1 0 31924 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_337
timestamp 1688980957
transform 1 0 32108 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_349
timestamp 1688980957
transform 1 0 33212 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_361
timestamp 1688980957
transform 1 0 34316 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_373
timestamp 1688980957
transform 1 0 35420 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_385
timestamp 1688980957
transform 1 0 36524 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_391
timestamp 1688980957
transform 1 0 37076 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_393
timestamp 1688980957
transform 1 0 37260 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_405
timestamp 1688980957
transform 1 0 38364 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_417
timestamp 1688980957
transform 1 0 39468 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_429
timestamp 1688980957
transform 1 0 40572 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_441
timestamp 1688980957
transform 1 0 41676 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_447
timestamp 1688980957
transform 1 0 42228 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_449
timestamp 1688980957
transform 1 0 42412 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_461
timestamp 1688980957
transform 1 0 43516 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_473
timestamp 1688980957
transform 1 0 44620 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_485
timestamp 1688980957
transform 1 0 45724 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_497
timestamp 1688980957
transform 1 0 46828 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_503
timestamp 1688980957
transform 1 0 47380 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_505
timestamp 1688980957
transform 1 0 47564 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_517
timestamp 1688980957
transform 1 0 48668 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_529
timestamp 1688980957
transform 1 0 49772 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_541
timestamp 1688980957
transform 1 0 50876 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_553
timestamp 1688980957
transform 1 0 51980 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_559
timestamp 1688980957
transform 1 0 52532 0 -1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_561
timestamp 1688980957
transform 1 0 52716 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_573
timestamp 1688980957
transform 1 0 53820 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_585
timestamp 1688980957
transform 1 0 54924 0 -1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_87_597
timestamp 1688980957
transform 1 0 56028 0 -1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87_609
timestamp 1688980957
transform 1 0 57132 0 -1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_87_615
timestamp 1688980957
transform 1 0 57684 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87_617
timestamp 1688980957
transform 1 0 57868 0 -1 50048
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_3
timestamp 1688980957
transform 1 0 1380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_15
timestamp 1688980957
transform 1 0 2484 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_27
timestamp 1688980957
transform 1 0 3588 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_29
timestamp 1688980957
transform 1 0 3772 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_41
timestamp 1688980957
transform 1 0 4876 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_53
timestamp 1688980957
transform 1 0 5980 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_65
timestamp 1688980957
transform 1 0 7084 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_77
timestamp 1688980957
transform 1 0 8188 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_83
timestamp 1688980957
transform 1 0 8740 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_85
timestamp 1688980957
transform 1 0 8924 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_97
timestamp 1688980957
transform 1 0 10028 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_109
timestamp 1688980957
transform 1 0 11132 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_121
timestamp 1688980957
transform 1 0 12236 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_133
timestamp 1688980957
transform 1 0 13340 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_139
timestamp 1688980957
transform 1 0 13892 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_141
timestamp 1688980957
transform 1 0 14076 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_153
timestamp 1688980957
transform 1 0 15180 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_165
timestamp 1688980957
transform 1 0 16284 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_177
timestamp 1688980957
transform 1 0 17388 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_189
timestamp 1688980957
transform 1 0 18492 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_195
timestamp 1688980957
transform 1 0 19044 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_197
timestamp 1688980957
transform 1 0 19228 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_209
timestamp 1688980957
transform 1 0 20332 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_221
timestamp 1688980957
transform 1 0 21436 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_233
timestamp 1688980957
transform 1 0 22540 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_245
timestamp 1688980957
transform 1 0 23644 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_251
timestamp 1688980957
transform 1 0 24196 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_253
timestamp 1688980957
transform 1 0 24380 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_265
timestamp 1688980957
transform 1 0 25484 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_277
timestamp 1688980957
transform 1 0 26588 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_289
timestamp 1688980957
transform 1 0 27692 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_301
timestamp 1688980957
transform 1 0 28796 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_307
timestamp 1688980957
transform 1 0 29348 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_309
timestamp 1688980957
transform 1 0 29532 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_321
timestamp 1688980957
transform 1 0 30636 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_333
timestamp 1688980957
transform 1 0 31740 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_345
timestamp 1688980957
transform 1 0 32844 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_357
timestamp 1688980957
transform 1 0 33948 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_363
timestamp 1688980957
transform 1 0 34500 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_365
timestamp 1688980957
transform 1 0 34684 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_377
timestamp 1688980957
transform 1 0 35788 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_389
timestamp 1688980957
transform 1 0 36892 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_401
timestamp 1688980957
transform 1 0 37996 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_413
timestamp 1688980957
transform 1 0 39100 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_419
timestamp 1688980957
transform 1 0 39652 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_421
timestamp 1688980957
transform 1 0 39836 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_433
timestamp 1688980957
transform 1 0 40940 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_445
timestamp 1688980957
transform 1 0 42044 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_457
timestamp 1688980957
transform 1 0 43148 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_469
timestamp 1688980957
transform 1 0 44252 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_475
timestamp 1688980957
transform 1 0 44804 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_477
timestamp 1688980957
transform 1 0 44988 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_489
timestamp 1688980957
transform 1 0 46092 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_501
timestamp 1688980957
transform 1 0 47196 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_513
timestamp 1688980957
transform 1 0 48300 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_525
timestamp 1688980957
transform 1 0 49404 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_531
timestamp 1688980957
transform 1 0 49956 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_533
timestamp 1688980957
transform 1 0 50140 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_545
timestamp 1688980957
transform 1 0 51244 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_557
timestamp 1688980957
transform 1 0 52348 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_569
timestamp 1688980957
transform 1 0 53452 0 1 50048
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_88_581
timestamp 1688980957
transform 1 0 54556 0 1 50048
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88_587
timestamp 1688980957
transform 1 0 55108 0 1 50048
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_589
timestamp 1688980957
transform 1 0 55292 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_601
timestamp 1688980957
transform 1 0 56396 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_88_613
timestamp 1688980957
transform 1 0 57500 0 1 50048
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_19
timestamp 1688980957
transform 1 0 2852 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_31
timestamp 1688980957
transform 1 0 3956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_43
timestamp 1688980957
transform 1 0 5060 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_55
timestamp 1688980957
transform 1 0 6164 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_57
timestamp 1688980957
transform 1 0 6348 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_69
timestamp 1688980957
transform 1 0 7452 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_81
timestamp 1688980957
transform 1 0 8556 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_93
timestamp 1688980957
transform 1 0 9660 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_105
timestamp 1688980957
transform 1 0 10764 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_111
timestamp 1688980957
transform 1 0 11316 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_113
timestamp 1688980957
transform 1 0 11500 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_125
timestamp 1688980957
transform 1 0 12604 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_137
timestamp 1688980957
transform 1 0 13708 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_149
timestamp 1688980957
transform 1 0 14812 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_161
timestamp 1688980957
transform 1 0 15916 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_167
timestamp 1688980957
transform 1 0 16468 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_169
timestamp 1688980957
transform 1 0 16652 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_181
timestamp 1688980957
transform 1 0 17756 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_193
timestamp 1688980957
transform 1 0 18860 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_205
timestamp 1688980957
transform 1 0 19964 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_217
timestamp 1688980957
transform 1 0 21068 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_223
timestamp 1688980957
transform 1 0 21620 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_225
timestamp 1688980957
transform 1 0 21804 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_237
timestamp 1688980957
transform 1 0 22908 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_249
timestamp 1688980957
transform 1 0 24012 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_261
timestamp 1688980957
transform 1 0 25116 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_273
timestamp 1688980957
transform 1 0 26220 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_279
timestamp 1688980957
transform 1 0 26772 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_281
timestamp 1688980957
transform 1 0 26956 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_293
timestamp 1688980957
transform 1 0 28060 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_305
timestamp 1688980957
transform 1 0 29164 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_317
timestamp 1688980957
transform 1 0 30268 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_329
timestamp 1688980957
transform 1 0 31372 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_335
timestamp 1688980957
transform 1 0 31924 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_337
timestamp 1688980957
transform 1 0 32108 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_349
timestamp 1688980957
transform 1 0 33212 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_361
timestamp 1688980957
transform 1 0 34316 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_373
timestamp 1688980957
transform 1 0 35420 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_385
timestamp 1688980957
transform 1 0 36524 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_391
timestamp 1688980957
transform 1 0 37076 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_393
timestamp 1688980957
transform 1 0 37260 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_405
timestamp 1688980957
transform 1 0 38364 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_417
timestamp 1688980957
transform 1 0 39468 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_429
timestamp 1688980957
transform 1 0 40572 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_441
timestamp 1688980957
transform 1 0 41676 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_447
timestamp 1688980957
transform 1 0 42228 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_449
timestamp 1688980957
transform 1 0 42412 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_461
timestamp 1688980957
transform 1 0 43516 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_473
timestamp 1688980957
transform 1 0 44620 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_485
timestamp 1688980957
transform 1 0 45724 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_497
timestamp 1688980957
transform 1 0 46828 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_503
timestamp 1688980957
transform 1 0 47380 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_505
timestamp 1688980957
transform 1 0 47564 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_517
timestamp 1688980957
transform 1 0 48668 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_529
timestamp 1688980957
transform 1 0 49772 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_541
timestamp 1688980957
transform 1 0 50876 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_553
timestamp 1688980957
transform 1 0 51980 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_559
timestamp 1688980957
transform 1 0 52532 0 -1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_561
timestamp 1688980957
transform 1 0 52716 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_573
timestamp 1688980957
transform 1 0 53820 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_585
timestamp 1688980957
transform 1 0 54924 0 -1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_89_597
timestamp 1688980957
transform 1 0 56028 0 -1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_89_609
timestamp 1688980957
transform 1 0 57132 0 -1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89_615
timestamp 1688980957
transform 1 0 57684 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_89_617
timestamp 1688980957
transform 1 0 57868 0 -1 51136
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_3
timestamp 1688980957
transform 1 0 1380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_15
timestamp 1688980957
transform 1 0 2484 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_27
timestamp 1688980957
transform 1 0 3588 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_29
timestamp 1688980957
transform 1 0 3772 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_41
timestamp 1688980957
transform 1 0 4876 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_53
timestamp 1688980957
transform 1 0 5980 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_65
timestamp 1688980957
transform 1 0 7084 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_77
timestamp 1688980957
transform 1 0 8188 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_83
timestamp 1688980957
transform 1 0 8740 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_85
timestamp 1688980957
transform 1 0 8924 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_97
timestamp 1688980957
transform 1 0 10028 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_109
timestamp 1688980957
transform 1 0 11132 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_121
timestamp 1688980957
transform 1 0 12236 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_133
timestamp 1688980957
transform 1 0 13340 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_139
timestamp 1688980957
transform 1 0 13892 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_141
timestamp 1688980957
transform 1 0 14076 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_153
timestamp 1688980957
transform 1 0 15180 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_165
timestamp 1688980957
transform 1 0 16284 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_177
timestamp 1688980957
transform 1 0 17388 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_189
timestamp 1688980957
transform 1 0 18492 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_195
timestamp 1688980957
transform 1 0 19044 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_197
timestamp 1688980957
transform 1 0 19228 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_209
timestamp 1688980957
transform 1 0 20332 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_221
timestamp 1688980957
transform 1 0 21436 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_233
timestamp 1688980957
transform 1 0 22540 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_245
timestamp 1688980957
transform 1 0 23644 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_251
timestamp 1688980957
transform 1 0 24196 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_253
timestamp 1688980957
transform 1 0 24380 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_265
timestamp 1688980957
transform 1 0 25484 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_277
timestamp 1688980957
transform 1 0 26588 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_289
timestamp 1688980957
transform 1 0 27692 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_301
timestamp 1688980957
transform 1 0 28796 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_307
timestamp 1688980957
transform 1 0 29348 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_309
timestamp 1688980957
transform 1 0 29532 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_321
timestamp 1688980957
transform 1 0 30636 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_333
timestamp 1688980957
transform 1 0 31740 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_345
timestamp 1688980957
transform 1 0 32844 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_357
timestamp 1688980957
transform 1 0 33948 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_363
timestamp 1688980957
transform 1 0 34500 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_365
timestamp 1688980957
transform 1 0 34684 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_377
timestamp 1688980957
transform 1 0 35788 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_389
timestamp 1688980957
transform 1 0 36892 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_401
timestamp 1688980957
transform 1 0 37996 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_413
timestamp 1688980957
transform 1 0 39100 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_419
timestamp 1688980957
transform 1 0 39652 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_421
timestamp 1688980957
transform 1 0 39836 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_433
timestamp 1688980957
transform 1 0 40940 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_445
timestamp 1688980957
transform 1 0 42044 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_457
timestamp 1688980957
transform 1 0 43148 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_469
timestamp 1688980957
transform 1 0 44252 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_475
timestamp 1688980957
transform 1 0 44804 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_477
timestamp 1688980957
transform 1 0 44988 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_489
timestamp 1688980957
transform 1 0 46092 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_501
timestamp 1688980957
transform 1 0 47196 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_513
timestamp 1688980957
transform 1 0 48300 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_525
timestamp 1688980957
transform 1 0 49404 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_531
timestamp 1688980957
transform 1 0 49956 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_533
timestamp 1688980957
transform 1 0 50140 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_545
timestamp 1688980957
transform 1 0 51244 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_557
timestamp 1688980957
transform 1 0 52348 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_569
timestamp 1688980957
transform 1 0 53452 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_581
timestamp 1688980957
transform 1 0 54556 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_90_587
timestamp 1688980957
transform 1 0 55108 0 1 51136
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_589
timestamp 1688980957
transform 1 0 55292 0 1 51136
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_90_601
timestamp 1688980957
transform 1 0 56396 0 1 51136
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_90_613
timestamp 1688980957
transform 1 0 57500 0 1 51136
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_3
timestamp 1688980957
transform 1 0 1380 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_15
timestamp 1688980957
transform 1 0 2484 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_27
timestamp 1688980957
transform 1 0 3588 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_39
timestamp 1688980957
transform 1 0 4692 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_91_51
timestamp 1688980957
transform 1 0 5796 0 -1 52224
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_55
timestamp 1688980957
transform 1 0 6164 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_57
timestamp 1688980957
transform 1 0 6348 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_69
timestamp 1688980957
transform 1 0 7452 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_81
timestamp 1688980957
transform 1 0 8556 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_93
timestamp 1688980957
transform 1 0 9660 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_105
timestamp 1688980957
transform 1 0 10764 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_111
timestamp 1688980957
transform 1 0 11316 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_113
timestamp 1688980957
transform 1 0 11500 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_125
timestamp 1688980957
transform 1 0 12604 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_137
timestamp 1688980957
transform 1 0 13708 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_149
timestamp 1688980957
transform 1 0 14812 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_161
timestamp 1688980957
transform 1 0 15916 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_167
timestamp 1688980957
transform 1 0 16468 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_169
timestamp 1688980957
transform 1 0 16652 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_181
timestamp 1688980957
transform 1 0 17756 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_193
timestamp 1688980957
transform 1 0 18860 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_205
timestamp 1688980957
transform 1 0 19964 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_217
timestamp 1688980957
transform 1 0 21068 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_223
timestamp 1688980957
transform 1 0 21620 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_225
timestamp 1688980957
transform 1 0 21804 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_237
timestamp 1688980957
transform 1 0 22908 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_249
timestamp 1688980957
transform 1 0 24012 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_261
timestamp 1688980957
transform 1 0 25116 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_273
timestamp 1688980957
transform 1 0 26220 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_279
timestamp 1688980957
transform 1 0 26772 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_281
timestamp 1688980957
transform 1 0 26956 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_293
timestamp 1688980957
transform 1 0 28060 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_305
timestamp 1688980957
transform 1 0 29164 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_317
timestamp 1688980957
transform 1 0 30268 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_329
timestamp 1688980957
transform 1 0 31372 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_335
timestamp 1688980957
transform 1 0 31924 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_337
timestamp 1688980957
transform 1 0 32108 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_349
timestamp 1688980957
transform 1 0 33212 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_361
timestamp 1688980957
transform 1 0 34316 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_373
timestamp 1688980957
transform 1 0 35420 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_385
timestamp 1688980957
transform 1 0 36524 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_391
timestamp 1688980957
transform 1 0 37076 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_393
timestamp 1688980957
transform 1 0 37260 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_405
timestamp 1688980957
transform 1 0 38364 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_417
timestamp 1688980957
transform 1 0 39468 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_429
timestamp 1688980957
transform 1 0 40572 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_441
timestamp 1688980957
transform 1 0 41676 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_447
timestamp 1688980957
transform 1 0 42228 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_449
timestamp 1688980957
transform 1 0 42412 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_461
timestamp 1688980957
transform 1 0 43516 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_473
timestamp 1688980957
transform 1 0 44620 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_485
timestamp 1688980957
transform 1 0 45724 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_497
timestamp 1688980957
transform 1 0 46828 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_503
timestamp 1688980957
transform 1 0 47380 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_505
timestamp 1688980957
transform 1 0 47564 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_517
timestamp 1688980957
transform 1 0 48668 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_529
timestamp 1688980957
transform 1 0 49772 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_541
timestamp 1688980957
transform 1 0 50876 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_553
timestamp 1688980957
transform 1 0 51980 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_559
timestamp 1688980957
transform 1 0 52532 0 -1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_561
timestamp 1688980957
transform 1 0 52716 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_573
timestamp 1688980957
transform 1 0 53820 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_585
timestamp 1688980957
transform 1 0 54924 0 -1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_91_597
timestamp 1688980957
transform 1 0 56028 0 -1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_91_609
timestamp 1688980957
transform 1 0 57132 0 -1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91_615
timestamp 1688980957
transform 1 0 57684 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_91_617
timestamp 1688980957
transform 1 0 57868 0 -1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_92_19
timestamp 1688980957
transform 1 0 2852 0 1 52224
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_27
timestamp 1688980957
transform 1 0 3588 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_29
timestamp 1688980957
transform 1 0 3772 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_41
timestamp 1688980957
transform 1 0 4876 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_53
timestamp 1688980957
transform 1 0 5980 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_65
timestamp 1688980957
transform 1 0 7084 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_77
timestamp 1688980957
transform 1 0 8188 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_83
timestamp 1688980957
transform 1 0 8740 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_85
timestamp 1688980957
transform 1 0 8924 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_97
timestamp 1688980957
transform 1 0 10028 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_109
timestamp 1688980957
transform 1 0 11132 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_121
timestamp 1688980957
transform 1 0 12236 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_133
timestamp 1688980957
transform 1 0 13340 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_139
timestamp 1688980957
transform 1 0 13892 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_141
timestamp 1688980957
transform 1 0 14076 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_153
timestamp 1688980957
transform 1 0 15180 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_165
timestamp 1688980957
transform 1 0 16284 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_177
timestamp 1688980957
transform 1 0 17388 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_189
timestamp 1688980957
transform 1 0 18492 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_195
timestamp 1688980957
transform 1 0 19044 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_197
timestamp 1688980957
transform 1 0 19228 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_209
timestamp 1688980957
transform 1 0 20332 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_221
timestamp 1688980957
transform 1 0 21436 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_233
timestamp 1688980957
transform 1 0 22540 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_245
timestamp 1688980957
transform 1 0 23644 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_251
timestamp 1688980957
transform 1 0 24196 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_253
timestamp 1688980957
transform 1 0 24380 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_265
timestamp 1688980957
transform 1 0 25484 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_277
timestamp 1688980957
transform 1 0 26588 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_289
timestamp 1688980957
transform 1 0 27692 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_301
timestamp 1688980957
transform 1 0 28796 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_307
timestamp 1688980957
transform 1 0 29348 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_309
timestamp 1688980957
transform 1 0 29532 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_321
timestamp 1688980957
transform 1 0 30636 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_333
timestamp 1688980957
transform 1 0 31740 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_345
timestamp 1688980957
transform 1 0 32844 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_357
timestamp 1688980957
transform 1 0 33948 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_363
timestamp 1688980957
transform 1 0 34500 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_365
timestamp 1688980957
transform 1 0 34684 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_377
timestamp 1688980957
transform 1 0 35788 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_389
timestamp 1688980957
transform 1 0 36892 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_401
timestamp 1688980957
transform 1 0 37996 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_413
timestamp 1688980957
transform 1 0 39100 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_419
timestamp 1688980957
transform 1 0 39652 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_421
timestamp 1688980957
transform 1 0 39836 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_433
timestamp 1688980957
transform 1 0 40940 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_445
timestamp 1688980957
transform 1 0 42044 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_457
timestamp 1688980957
transform 1 0 43148 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_469
timestamp 1688980957
transform 1 0 44252 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_475
timestamp 1688980957
transform 1 0 44804 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_477
timestamp 1688980957
transform 1 0 44988 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_489
timestamp 1688980957
transform 1 0 46092 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_501
timestamp 1688980957
transform 1 0 47196 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_513
timestamp 1688980957
transform 1 0 48300 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_525
timestamp 1688980957
transform 1 0 49404 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_531
timestamp 1688980957
transform 1 0 49956 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_533
timestamp 1688980957
transform 1 0 50140 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_545
timestamp 1688980957
transform 1 0 51244 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_557
timestamp 1688980957
transform 1 0 52348 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_569
timestamp 1688980957
transform 1 0 53452 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_581
timestamp 1688980957
transform 1 0 54556 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92_587
timestamp 1688980957
transform 1 0 55108 0 1 52224
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_589
timestamp 1688980957
transform 1 0 55292 0 1 52224
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_92_601
timestamp 1688980957
transform 1 0 56396 0 1 52224
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_92_613
timestamp 1688980957
transform 1 0 57500 0 1 52224
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_3
timestamp 1688980957
transform 1 0 1380 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_15
timestamp 1688980957
transform 1 0 2484 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_27
timestamp 1688980957
transform 1 0 3588 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_39
timestamp 1688980957
transform 1 0 4692 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_51
timestamp 1688980957
transform 1 0 5796 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_55
timestamp 1688980957
transform 1 0 6164 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_57
timestamp 1688980957
transform 1 0 6348 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_69
timestamp 1688980957
transform 1 0 7452 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_81
timestamp 1688980957
transform 1 0 8556 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_93
timestamp 1688980957
transform 1 0 9660 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_105
timestamp 1688980957
transform 1 0 10764 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_111
timestamp 1688980957
transform 1 0 11316 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_113
timestamp 1688980957
transform 1 0 11500 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_125
timestamp 1688980957
transform 1 0 12604 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_137
timestamp 1688980957
transform 1 0 13708 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_149
timestamp 1688980957
transform 1 0 14812 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_161
timestamp 1688980957
transform 1 0 15916 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_167
timestamp 1688980957
transform 1 0 16468 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_169
timestamp 1688980957
transform 1 0 16652 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_181
timestamp 1688980957
transform 1 0 17756 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_193
timestamp 1688980957
transform 1 0 18860 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_205
timestamp 1688980957
transform 1 0 19964 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_217
timestamp 1688980957
transform 1 0 21068 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_223
timestamp 1688980957
transform 1 0 21620 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_225
timestamp 1688980957
transform 1 0 21804 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_237
timestamp 1688980957
transform 1 0 22908 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_249
timestamp 1688980957
transform 1 0 24012 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_261
timestamp 1688980957
transform 1 0 25116 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_273
timestamp 1688980957
transform 1 0 26220 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_279
timestamp 1688980957
transform 1 0 26772 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_281
timestamp 1688980957
transform 1 0 26956 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_293
timestamp 1688980957
transform 1 0 28060 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_305
timestamp 1688980957
transform 1 0 29164 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_317
timestamp 1688980957
transform 1 0 30268 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_329
timestamp 1688980957
transform 1 0 31372 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_335
timestamp 1688980957
transform 1 0 31924 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_337
timestamp 1688980957
transform 1 0 32108 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_349
timestamp 1688980957
transform 1 0 33212 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_361
timestamp 1688980957
transform 1 0 34316 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_373
timestamp 1688980957
transform 1 0 35420 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_385
timestamp 1688980957
transform 1 0 36524 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_391
timestamp 1688980957
transform 1 0 37076 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_393
timestamp 1688980957
transform 1 0 37260 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_405
timestamp 1688980957
transform 1 0 38364 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_417
timestamp 1688980957
transform 1 0 39468 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_429
timestamp 1688980957
transform 1 0 40572 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_441
timestamp 1688980957
transform 1 0 41676 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_447
timestamp 1688980957
transform 1 0 42228 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_449
timestamp 1688980957
transform 1 0 42412 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_461
timestamp 1688980957
transform 1 0 43516 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_473
timestamp 1688980957
transform 1 0 44620 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_485
timestamp 1688980957
transform 1 0 45724 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_497
timestamp 1688980957
transform 1 0 46828 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_503
timestamp 1688980957
transform 1 0 47380 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_505
timestamp 1688980957
transform 1 0 47564 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_517
timestamp 1688980957
transform 1 0 48668 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_529
timestamp 1688980957
transform 1 0 49772 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_541
timestamp 1688980957
transform 1 0 50876 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_553
timestamp 1688980957
transform 1 0 51980 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_559
timestamp 1688980957
transform 1 0 52532 0 -1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_561
timestamp 1688980957
transform 1 0 52716 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_573
timestamp 1688980957
transform 1 0 53820 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_585
timestamp 1688980957
transform 1 0 54924 0 -1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_93_597
timestamp 1688980957
transform 1 0 56028 0 -1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_93_609
timestamp 1688980957
transform 1 0 57132 0 -1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93_615
timestamp 1688980957
transform 1 0 57684 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_93_617
timestamp 1688980957
transform 1 0 57868 0 -1 53312
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_3
timestamp 1688980957
transform 1 0 1380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_15
timestamp 1688980957
transform 1 0 2484 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_27
timestamp 1688980957
transform 1 0 3588 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_29
timestamp 1688980957
transform 1 0 3772 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_41
timestamp 1688980957
transform 1 0 4876 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_53
timestamp 1688980957
transform 1 0 5980 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_65
timestamp 1688980957
transform 1 0 7084 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_77
timestamp 1688980957
transform 1 0 8188 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_83
timestamp 1688980957
transform 1 0 8740 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_85
timestamp 1688980957
transform 1 0 8924 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_97
timestamp 1688980957
transform 1 0 10028 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_109
timestamp 1688980957
transform 1 0 11132 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_121
timestamp 1688980957
transform 1 0 12236 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_133
timestamp 1688980957
transform 1 0 13340 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_139
timestamp 1688980957
transform 1 0 13892 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_141
timestamp 1688980957
transform 1 0 14076 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_153
timestamp 1688980957
transform 1 0 15180 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_165
timestamp 1688980957
transform 1 0 16284 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_177
timestamp 1688980957
transform 1 0 17388 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_189
timestamp 1688980957
transform 1 0 18492 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_195
timestamp 1688980957
transform 1 0 19044 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_197
timestamp 1688980957
transform 1 0 19228 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_209
timestamp 1688980957
transform 1 0 20332 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_221
timestamp 1688980957
transform 1 0 21436 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_233
timestamp 1688980957
transform 1 0 22540 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_245
timestamp 1688980957
transform 1 0 23644 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_251
timestamp 1688980957
transform 1 0 24196 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_253
timestamp 1688980957
transform 1 0 24380 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_265
timestamp 1688980957
transform 1 0 25484 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_277
timestamp 1688980957
transform 1 0 26588 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_289
timestamp 1688980957
transform 1 0 27692 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_301
timestamp 1688980957
transform 1 0 28796 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_307
timestamp 1688980957
transform 1 0 29348 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_309
timestamp 1688980957
transform 1 0 29532 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_321
timestamp 1688980957
transform 1 0 30636 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_333
timestamp 1688980957
transform 1 0 31740 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_345
timestamp 1688980957
transform 1 0 32844 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_357
timestamp 1688980957
transform 1 0 33948 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_363
timestamp 1688980957
transform 1 0 34500 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_365
timestamp 1688980957
transform 1 0 34684 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_377
timestamp 1688980957
transform 1 0 35788 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_389
timestamp 1688980957
transform 1 0 36892 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_401
timestamp 1688980957
transform 1 0 37996 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_413
timestamp 1688980957
transform 1 0 39100 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_419
timestamp 1688980957
transform 1 0 39652 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_421
timestamp 1688980957
transform 1 0 39836 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_433
timestamp 1688980957
transform 1 0 40940 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_445
timestamp 1688980957
transform 1 0 42044 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_457
timestamp 1688980957
transform 1 0 43148 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_469
timestamp 1688980957
transform 1 0 44252 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_475
timestamp 1688980957
transform 1 0 44804 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_477
timestamp 1688980957
transform 1 0 44988 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_489
timestamp 1688980957
transform 1 0 46092 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_501
timestamp 1688980957
transform 1 0 47196 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_513
timestamp 1688980957
transform 1 0 48300 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_525
timestamp 1688980957
transform 1 0 49404 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_531
timestamp 1688980957
transform 1 0 49956 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_533
timestamp 1688980957
transform 1 0 50140 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_545
timestamp 1688980957
transform 1 0 51244 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_557
timestamp 1688980957
transform 1 0 52348 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_569
timestamp 1688980957
transform 1 0 53452 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94_581
timestamp 1688980957
transform 1 0 54556 0 1 53312
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_94_587
timestamp 1688980957
transform 1 0 55108 0 1 53312
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_589
timestamp 1688980957
transform 1 0 55292 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_601
timestamp 1688980957
transform 1 0 56396 0 1 53312
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_94_613
timestamp 1688980957
transform 1 0 57500 0 1 53312
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_95_19
timestamp 1688980957
transform 1 0 2852 0 -1 54400
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_23
timestamp 1688980957
transform 1 0 3220 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_35
timestamp 1688980957
transform 1 0 4324 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_47
timestamp 1688980957
transform 1 0 5428 0 -1 54400
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_55
timestamp 1688980957
transform 1 0 6164 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_57
timestamp 1688980957
transform 1 0 6348 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_69
timestamp 1688980957
transform 1 0 7452 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_81
timestamp 1688980957
transform 1 0 8556 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_93
timestamp 1688980957
transform 1 0 9660 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_105
timestamp 1688980957
transform 1 0 10764 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_111
timestamp 1688980957
transform 1 0 11316 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_113
timestamp 1688980957
transform 1 0 11500 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_125
timestamp 1688980957
transform 1 0 12604 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_137
timestamp 1688980957
transform 1 0 13708 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_149
timestamp 1688980957
transform 1 0 14812 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_161
timestamp 1688980957
transform 1 0 15916 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_167
timestamp 1688980957
transform 1 0 16468 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_169
timestamp 1688980957
transform 1 0 16652 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_181
timestamp 1688980957
transform 1 0 17756 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_193
timestamp 1688980957
transform 1 0 18860 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_205
timestamp 1688980957
transform 1 0 19964 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_217
timestamp 1688980957
transform 1 0 21068 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_223
timestamp 1688980957
transform 1 0 21620 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_225
timestamp 1688980957
transform 1 0 21804 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_237
timestamp 1688980957
transform 1 0 22908 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_249
timestamp 1688980957
transform 1 0 24012 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_261
timestamp 1688980957
transform 1 0 25116 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_273
timestamp 1688980957
transform 1 0 26220 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_279
timestamp 1688980957
transform 1 0 26772 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_281
timestamp 1688980957
transform 1 0 26956 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_293
timestamp 1688980957
transform 1 0 28060 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_305
timestamp 1688980957
transform 1 0 29164 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_317
timestamp 1688980957
transform 1 0 30268 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_329
timestamp 1688980957
transform 1 0 31372 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_335
timestamp 1688980957
transform 1 0 31924 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_337
timestamp 1688980957
transform 1 0 32108 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_349
timestamp 1688980957
transform 1 0 33212 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_361
timestamp 1688980957
transform 1 0 34316 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_373
timestamp 1688980957
transform 1 0 35420 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_385
timestamp 1688980957
transform 1 0 36524 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_391
timestamp 1688980957
transform 1 0 37076 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_393
timestamp 1688980957
transform 1 0 37260 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_405
timestamp 1688980957
transform 1 0 38364 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_417
timestamp 1688980957
transform 1 0 39468 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_429
timestamp 1688980957
transform 1 0 40572 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_441
timestamp 1688980957
transform 1 0 41676 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_447
timestamp 1688980957
transform 1 0 42228 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_449
timestamp 1688980957
transform 1 0 42412 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_461
timestamp 1688980957
transform 1 0 43516 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_473
timestamp 1688980957
transform 1 0 44620 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_485
timestamp 1688980957
transform 1 0 45724 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_497
timestamp 1688980957
transform 1 0 46828 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_503
timestamp 1688980957
transform 1 0 47380 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_505
timestamp 1688980957
transform 1 0 47564 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_517
timestamp 1688980957
transform 1 0 48668 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_529
timestamp 1688980957
transform 1 0 49772 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_541
timestamp 1688980957
transform 1 0 50876 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_553
timestamp 1688980957
transform 1 0 51980 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_559
timestamp 1688980957
transform 1 0 52532 0 -1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_561
timestamp 1688980957
transform 1 0 52716 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_573
timestamp 1688980957
transform 1 0 53820 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_585
timestamp 1688980957
transform 1 0 54924 0 -1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_95_597
timestamp 1688980957
transform 1 0 56028 0 -1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_95_609
timestamp 1688980957
transform 1 0 57132 0 -1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_95_615
timestamp 1688980957
transform 1 0 57684 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_95_617
timestamp 1688980957
transform 1 0 57868 0 -1 54400
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_3
timestamp 1688980957
transform 1 0 1380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_15
timestamp 1688980957
transform 1 0 2484 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_27
timestamp 1688980957
transform 1 0 3588 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_29
timestamp 1688980957
transform 1 0 3772 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_41
timestamp 1688980957
transform 1 0 4876 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_53
timestamp 1688980957
transform 1 0 5980 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_65
timestamp 1688980957
transform 1 0 7084 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_77
timestamp 1688980957
transform 1 0 8188 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_83
timestamp 1688980957
transform 1 0 8740 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_85
timestamp 1688980957
transform 1 0 8924 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_97
timestamp 1688980957
transform 1 0 10028 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_109
timestamp 1688980957
transform 1 0 11132 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_121
timestamp 1688980957
transform 1 0 12236 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_133
timestamp 1688980957
transform 1 0 13340 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_139
timestamp 1688980957
transform 1 0 13892 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_141
timestamp 1688980957
transform 1 0 14076 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_153
timestamp 1688980957
transform 1 0 15180 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_165
timestamp 1688980957
transform 1 0 16284 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_177
timestamp 1688980957
transform 1 0 17388 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_189
timestamp 1688980957
transform 1 0 18492 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_195
timestamp 1688980957
transform 1 0 19044 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_197
timestamp 1688980957
transform 1 0 19228 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_209
timestamp 1688980957
transform 1 0 20332 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_221
timestamp 1688980957
transform 1 0 21436 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_233
timestamp 1688980957
transform 1 0 22540 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_245
timestamp 1688980957
transform 1 0 23644 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_251
timestamp 1688980957
transform 1 0 24196 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_253
timestamp 1688980957
transform 1 0 24380 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_265
timestamp 1688980957
transform 1 0 25484 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_277
timestamp 1688980957
transform 1 0 26588 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_289
timestamp 1688980957
transform 1 0 27692 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_301
timestamp 1688980957
transform 1 0 28796 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_307
timestamp 1688980957
transform 1 0 29348 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_309
timestamp 1688980957
transform 1 0 29532 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_321
timestamp 1688980957
transform 1 0 30636 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_333
timestamp 1688980957
transform 1 0 31740 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_345
timestamp 1688980957
transform 1 0 32844 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_357
timestamp 1688980957
transform 1 0 33948 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_363
timestamp 1688980957
transform 1 0 34500 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_365
timestamp 1688980957
transform 1 0 34684 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_377
timestamp 1688980957
transform 1 0 35788 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_389
timestamp 1688980957
transform 1 0 36892 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_401
timestamp 1688980957
transform 1 0 37996 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_413
timestamp 1688980957
transform 1 0 39100 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_419
timestamp 1688980957
transform 1 0 39652 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_421
timestamp 1688980957
transform 1 0 39836 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_433
timestamp 1688980957
transform 1 0 40940 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_445
timestamp 1688980957
transform 1 0 42044 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_457
timestamp 1688980957
transform 1 0 43148 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_469
timestamp 1688980957
transform 1 0 44252 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_475
timestamp 1688980957
transform 1 0 44804 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_477
timestamp 1688980957
transform 1 0 44988 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_489
timestamp 1688980957
transform 1 0 46092 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_501
timestamp 1688980957
transform 1 0 47196 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_513
timestamp 1688980957
transform 1 0 48300 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_525
timestamp 1688980957
transform 1 0 49404 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_531
timestamp 1688980957
transform 1 0 49956 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_533
timestamp 1688980957
transform 1 0 50140 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_545
timestamp 1688980957
transform 1 0 51244 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_557
timestamp 1688980957
transform 1 0 52348 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_569
timestamp 1688980957
transform 1 0 53452 0 1 54400
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_96_581
timestamp 1688980957
transform 1 0 54556 0 1 54400
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_96_587
timestamp 1688980957
transform 1 0 55108 0 1 54400
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_589
timestamp 1688980957
transform 1 0 55292 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_601
timestamp 1688980957
transform 1 0 56396 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_96_613
timestamp 1688980957
transform 1 0 57500 0 1 54400
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_3
timestamp 1688980957
transform 1 0 1380 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_15
timestamp 1688980957
transform 1 0 2484 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_27
timestamp 1688980957
transform 1 0 3588 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_39
timestamp 1688980957
transform 1 0 4692 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97_51
timestamp 1688980957
transform 1 0 5796 0 -1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_55
timestamp 1688980957
transform 1 0 6164 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_57
timestamp 1688980957
transform 1 0 6348 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_69
timestamp 1688980957
transform 1 0 7452 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_81
timestamp 1688980957
transform 1 0 8556 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_93
timestamp 1688980957
transform 1 0 9660 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_105
timestamp 1688980957
transform 1 0 10764 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_111
timestamp 1688980957
transform 1 0 11316 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_113
timestamp 1688980957
transform 1 0 11500 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_125
timestamp 1688980957
transform 1 0 12604 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_137
timestamp 1688980957
transform 1 0 13708 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_149
timestamp 1688980957
transform 1 0 14812 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_161
timestamp 1688980957
transform 1 0 15916 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_167
timestamp 1688980957
transform 1 0 16468 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_169
timestamp 1688980957
transform 1 0 16652 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_181
timestamp 1688980957
transform 1 0 17756 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_193
timestamp 1688980957
transform 1 0 18860 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_205
timestamp 1688980957
transform 1 0 19964 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_217
timestamp 1688980957
transform 1 0 21068 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_223
timestamp 1688980957
transform 1 0 21620 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_225
timestamp 1688980957
transform 1 0 21804 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_237
timestamp 1688980957
transform 1 0 22908 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_249
timestamp 1688980957
transform 1 0 24012 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_261
timestamp 1688980957
transform 1 0 25116 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_273
timestamp 1688980957
transform 1 0 26220 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_279
timestamp 1688980957
transform 1 0 26772 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_281
timestamp 1688980957
transform 1 0 26956 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_293
timestamp 1688980957
transform 1 0 28060 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_305
timestamp 1688980957
transform 1 0 29164 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_317
timestamp 1688980957
transform 1 0 30268 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_329
timestamp 1688980957
transform 1 0 31372 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_335
timestamp 1688980957
transform 1 0 31924 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_337
timestamp 1688980957
transform 1 0 32108 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_349
timestamp 1688980957
transform 1 0 33212 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_361
timestamp 1688980957
transform 1 0 34316 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_373
timestamp 1688980957
transform 1 0 35420 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_385
timestamp 1688980957
transform 1 0 36524 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_391
timestamp 1688980957
transform 1 0 37076 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_393
timestamp 1688980957
transform 1 0 37260 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_405
timestamp 1688980957
transform 1 0 38364 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_417
timestamp 1688980957
transform 1 0 39468 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_429
timestamp 1688980957
transform 1 0 40572 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_441
timestamp 1688980957
transform 1 0 41676 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_447
timestamp 1688980957
transform 1 0 42228 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_449
timestamp 1688980957
transform 1 0 42412 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_461
timestamp 1688980957
transform 1 0 43516 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_473
timestamp 1688980957
transform 1 0 44620 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_485
timestamp 1688980957
transform 1 0 45724 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_497
timestamp 1688980957
transform 1 0 46828 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_503
timestamp 1688980957
transform 1 0 47380 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_505
timestamp 1688980957
transform 1 0 47564 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_517
timestamp 1688980957
transform 1 0 48668 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_529
timestamp 1688980957
transform 1 0 49772 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_541
timestamp 1688980957
transform 1 0 50876 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_553
timestamp 1688980957
transform 1 0 51980 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_559
timestamp 1688980957
transform 1 0 52532 0 -1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_561
timestamp 1688980957
transform 1 0 52716 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_573
timestamp 1688980957
transform 1 0 53820 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_585
timestamp 1688980957
transform 1 0 54924 0 -1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97_597
timestamp 1688980957
transform 1 0 56028 0 -1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_97_609
timestamp 1688980957
transform 1 0 57132 0 -1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_97_615
timestamp 1688980957
transform 1 0 57684 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_97_617
timestamp 1688980957
transform 1 0 57868 0 -1 55488
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98_19
timestamp 1688980957
transform 1 0 2852 0 1 55488
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_98_23
timestamp 1688980957
transform 1 0 3220 0 1 55488
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_27
timestamp 1688980957
transform 1 0 3588 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_29
timestamp 1688980957
transform 1 0 3772 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_41
timestamp 1688980957
transform 1 0 4876 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_53
timestamp 1688980957
transform 1 0 5980 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_65
timestamp 1688980957
transform 1 0 7084 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_77
timestamp 1688980957
transform 1 0 8188 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_83
timestamp 1688980957
transform 1 0 8740 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_85
timestamp 1688980957
transform 1 0 8924 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_97
timestamp 1688980957
transform 1 0 10028 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_109
timestamp 1688980957
transform 1 0 11132 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_121
timestamp 1688980957
transform 1 0 12236 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_133
timestamp 1688980957
transform 1 0 13340 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_139
timestamp 1688980957
transform 1 0 13892 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_141
timestamp 1688980957
transform 1 0 14076 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_153
timestamp 1688980957
transform 1 0 15180 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_165
timestamp 1688980957
transform 1 0 16284 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_177
timestamp 1688980957
transform 1 0 17388 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_189
timestamp 1688980957
transform 1 0 18492 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_195
timestamp 1688980957
transform 1 0 19044 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_197
timestamp 1688980957
transform 1 0 19228 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_209
timestamp 1688980957
transform 1 0 20332 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_221
timestamp 1688980957
transform 1 0 21436 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_233
timestamp 1688980957
transform 1 0 22540 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_245
timestamp 1688980957
transform 1 0 23644 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_251
timestamp 1688980957
transform 1 0 24196 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_253
timestamp 1688980957
transform 1 0 24380 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_265
timestamp 1688980957
transform 1 0 25484 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_277
timestamp 1688980957
transform 1 0 26588 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_289
timestamp 1688980957
transform 1 0 27692 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_301
timestamp 1688980957
transform 1 0 28796 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_307
timestamp 1688980957
transform 1 0 29348 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_309
timestamp 1688980957
transform 1 0 29532 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_321
timestamp 1688980957
transform 1 0 30636 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_333
timestamp 1688980957
transform 1 0 31740 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_345
timestamp 1688980957
transform 1 0 32844 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_357
timestamp 1688980957
transform 1 0 33948 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_363
timestamp 1688980957
transform 1 0 34500 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_365
timestamp 1688980957
transform 1 0 34684 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_377
timestamp 1688980957
transform 1 0 35788 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_389
timestamp 1688980957
transform 1 0 36892 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_401
timestamp 1688980957
transform 1 0 37996 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_413
timestamp 1688980957
transform 1 0 39100 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_419
timestamp 1688980957
transform 1 0 39652 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_421
timestamp 1688980957
transform 1 0 39836 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_433
timestamp 1688980957
transform 1 0 40940 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_445
timestamp 1688980957
transform 1 0 42044 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_457
timestamp 1688980957
transform 1 0 43148 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_469
timestamp 1688980957
transform 1 0 44252 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_475
timestamp 1688980957
transform 1 0 44804 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_477
timestamp 1688980957
transform 1 0 44988 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_489
timestamp 1688980957
transform 1 0 46092 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_501
timestamp 1688980957
transform 1 0 47196 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_513
timestamp 1688980957
transform 1 0 48300 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_525
timestamp 1688980957
transform 1 0 49404 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_531
timestamp 1688980957
transform 1 0 49956 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_533
timestamp 1688980957
transform 1 0 50140 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_545
timestamp 1688980957
transform 1 0 51244 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_557
timestamp 1688980957
transform 1 0 52348 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_569
timestamp 1688980957
transform 1 0 53452 0 1 55488
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98_581
timestamp 1688980957
transform 1 0 54556 0 1 55488
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_98_587
timestamp 1688980957
transform 1 0 55108 0 1 55488
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_589
timestamp 1688980957
transform 1 0 55292 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_601
timestamp 1688980957
transform 1 0 56396 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_98_613
timestamp 1688980957
transform 1 0 57500 0 1 55488
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_3
timestamp 1688980957
transform 1 0 1380 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_15
timestamp 1688980957
transform 1 0 2484 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_27
timestamp 1688980957
transform 1 0 3588 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_39
timestamp 1688980957
transform 1 0 4692 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_99_51
timestamp 1688980957
transform 1 0 5796 0 -1 56576
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_55
timestamp 1688980957
transform 1 0 6164 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_57
timestamp 1688980957
transform 1 0 6348 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_69
timestamp 1688980957
transform 1 0 7452 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_81
timestamp 1688980957
transform 1 0 8556 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_93
timestamp 1688980957
transform 1 0 9660 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_105
timestamp 1688980957
transform 1 0 10764 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_111
timestamp 1688980957
transform 1 0 11316 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_113
timestamp 1688980957
transform 1 0 11500 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_125
timestamp 1688980957
transform 1 0 12604 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_137
timestamp 1688980957
transform 1 0 13708 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_149
timestamp 1688980957
transform 1 0 14812 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_161
timestamp 1688980957
transform 1 0 15916 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_167
timestamp 1688980957
transform 1 0 16468 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_169
timestamp 1688980957
transform 1 0 16652 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_181
timestamp 1688980957
transform 1 0 17756 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_193
timestamp 1688980957
transform 1 0 18860 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_205
timestamp 1688980957
transform 1 0 19964 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_217
timestamp 1688980957
transform 1 0 21068 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_223
timestamp 1688980957
transform 1 0 21620 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_225
timestamp 1688980957
transform 1 0 21804 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_237
timestamp 1688980957
transform 1 0 22908 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_249
timestamp 1688980957
transform 1 0 24012 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_261
timestamp 1688980957
transform 1 0 25116 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_273
timestamp 1688980957
transform 1 0 26220 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_279
timestamp 1688980957
transform 1 0 26772 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_281
timestamp 1688980957
transform 1 0 26956 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_293
timestamp 1688980957
transform 1 0 28060 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_305
timestamp 1688980957
transform 1 0 29164 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_317
timestamp 1688980957
transform 1 0 30268 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_329
timestamp 1688980957
transform 1 0 31372 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_335
timestamp 1688980957
transform 1 0 31924 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_337
timestamp 1688980957
transform 1 0 32108 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_349
timestamp 1688980957
transform 1 0 33212 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_361
timestamp 1688980957
transform 1 0 34316 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_373
timestamp 1688980957
transform 1 0 35420 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_385
timestamp 1688980957
transform 1 0 36524 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_391
timestamp 1688980957
transform 1 0 37076 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_393
timestamp 1688980957
transform 1 0 37260 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_405
timestamp 1688980957
transform 1 0 38364 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_417
timestamp 1688980957
transform 1 0 39468 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_429
timestamp 1688980957
transform 1 0 40572 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_441
timestamp 1688980957
transform 1 0 41676 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_447
timestamp 1688980957
transform 1 0 42228 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_449
timestamp 1688980957
transform 1 0 42412 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_461
timestamp 1688980957
transform 1 0 43516 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_473
timestamp 1688980957
transform 1 0 44620 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_485
timestamp 1688980957
transform 1 0 45724 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_497
timestamp 1688980957
transform 1 0 46828 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_503
timestamp 1688980957
transform 1 0 47380 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_505
timestamp 1688980957
transform 1 0 47564 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_517
timestamp 1688980957
transform 1 0 48668 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_529
timestamp 1688980957
transform 1 0 49772 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_541
timestamp 1688980957
transform 1 0 50876 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_553
timestamp 1688980957
transform 1 0 51980 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_559
timestamp 1688980957
transform 1 0 52532 0 -1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_561
timestamp 1688980957
transform 1 0 52716 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_573
timestamp 1688980957
transform 1 0 53820 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_585
timestamp 1688980957
transform 1 0 54924 0 -1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_99_597
timestamp 1688980957
transform 1 0 56028 0 -1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_99_609
timestamp 1688980957
transform 1 0 57132 0 -1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_99_615
timestamp 1688980957
transform 1 0 57684 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_99_617
timestamp 1688980957
transform 1 0 57868 0 -1 56576
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_3
timestamp 1688980957
transform 1 0 1380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_15
timestamp 1688980957
transform 1 0 2484 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_27
timestamp 1688980957
transform 1 0 3588 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_29
timestamp 1688980957
transform 1 0 3772 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_41
timestamp 1688980957
transform 1 0 4876 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_53
timestamp 1688980957
transform 1 0 5980 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_65
timestamp 1688980957
transform 1 0 7084 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_77
timestamp 1688980957
transform 1 0 8188 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_83
timestamp 1688980957
transform 1 0 8740 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_85
timestamp 1688980957
transform 1 0 8924 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_97
timestamp 1688980957
transform 1 0 10028 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_109
timestamp 1688980957
transform 1 0 11132 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_121
timestamp 1688980957
transform 1 0 12236 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_133
timestamp 1688980957
transform 1 0 13340 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_139
timestamp 1688980957
transform 1 0 13892 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_141
timestamp 1688980957
transform 1 0 14076 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_153
timestamp 1688980957
transform 1 0 15180 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_165
timestamp 1688980957
transform 1 0 16284 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_177
timestamp 1688980957
transform 1 0 17388 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_189
timestamp 1688980957
transform 1 0 18492 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_195
timestamp 1688980957
transform 1 0 19044 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_197
timestamp 1688980957
transform 1 0 19228 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_209
timestamp 1688980957
transform 1 0 20332 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_221
timestamp 1688980957
transform 1 0 21436 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_233
timestamp 1688980957
transform 1 0 22540 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_245
timestamp 1688980957
transform 1 0 23644 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_251
timestamp 1688980957
transform 1 0 24196 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_253
timestamp 1688980957
transform 1 0 24380 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_265
timestamp 1688980957
transform 1 0 25484 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_277
timestamp 1688980957
transform 1 0 26588 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_289
timestamp 1688980957
transform 1 0 27692 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_301
timestamp 1688980957
transform 1 0 28796 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_307
timestamp 1688980957
transform 1 0 29348 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_309
timestamp 1688980957
transform 1 0 29532 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_321
timestamp 1688980957
transform 1 0 30636 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_333
timestamp 1688980957
transform 1 0 31740 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_345
timestamp 1688980957
transform 1 0 32844 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_357
timestamp 1688980957
transform 1 0 33948 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_363
timestamp 1688980957
transform 1 0 34500 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_365
timestamp 1688980957
transform 1 0 34684 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_377
timestamp 1688980957
transform 1 0 35788 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_389
timestamp 1688980957
transform 1 0 36892 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_401
timestamp 1688980957
transform 1 0 37996 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_413
timestamp 1688980957
transform 1 0 39100 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_419
timestamp 1688980957
transform 1 0 39652 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_421
timestamp 1688980957
transform 1 0 39836 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_433
timestamp 1688980957
transform 1 0 40940 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_445
timestamp 1688980957
transform 1 0 42044 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_457
timestamp 1688980957
transform 1 0 43148 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_469
timestamp 1688980957
transform 1 0 44252 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_475
timestamp 1688980957
transform 1 0 44804 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_477
timestamp 1688980957
transform 1 0 44988 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_489
timestamp 1688980957
transform 1 0 46092 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_501
timestamp 1688980957
transform 1 0 47196 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_513
timestamp 1688980957
transform 1 0 48300 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_525
timestamp 1688980957
transform 1 0 49404 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_531
timestamp 1688980957
transform 1 0 49956 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_533
timestamp 1688980957
transform 1 0 50140 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_545
timestamp 1688980957
transform 1 0 51244 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_557
timestamp 1688980957
transform 1 0 52348 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_569
timestamp 1688980957
transform 1 0 53452 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_100_581
timestamp 1688980957
transform 1 0 54556 0 1 56576
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100_587
timestamp 1688980957
transform 1 0 55108 0 1 56576
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_589
timestamp 1688980957
transform 1 0 55292 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_601
timestamp 1688980957
transform 1 0 56396 0 1 56576
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_100_613
timestamp 1688980957
transform 1 0 57500 0 1 56576
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_101_19
timestamp 1688980957
transform 1 0 2852 0 -1 57664
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_23
timestamp 1688980957
transform 1 0 3220 0 -1 57664
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_101_27
timestamp 1688980957
transform 1 0 3588 0 -1 57664
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_29
timestamp 1688980957
transform 1 0 3772 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_41
timestamp 1688980957
transform 1 0 4876 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_53
timestamp 1688980957
transform 1 0 5980 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_57
timestamp 1688980957
transform 1 0 6348 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_69
timestamp 1688980957
transform 1 0 7452 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_81
timestamp 1688980957
transform 1 0 8556 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_85
timestamp 1688980957
transform 1 0 8924 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_97
timestamp 1688980957
transform 1 0 10028 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_109
timestamp 1688980957
transform 1 0 11132 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_113
timestamp 1688980957
transform 1 0 11500 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_125
timestamp 1688980957
transform 1 0 12604 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_137
timestamp 1688980957
transform 1 0 13708 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_141
timestamp 1688980957
transform 1 0 14076 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_153
timestamp 1688980957
transform 1 0 15180 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_165
timestamp 1688980957
transform 1 0 16284 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_169
timestamp 1688980957
transform 1 0 16652 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_181
timestamp 1688980957
transform 1 0 17756 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_193
timestamp 1688980957
transform 1 0 18860 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_197
timestamp 1688980957
transform 1 0 19228 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_209
timestamp 1688980957
transform 1 0 20332 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_221
timestamp 1688980957
transform 1 0 21436 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_225
timestamp 1688980957
transform 1 0 21804 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_237
timestamp 1688980957
transform 1 0 22908 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_249
timestamp 1688980957
transform 1 0 24012 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_253
timestamp 1688980957
transform 1 0 24380 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_265
timestamp 1688980957
transform 1 0 25484 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_277
timestamp 1688980957
transform 1 0 26588 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_281
timestamp 1688980957
transform 1 0 26956 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_293
timestamp 1688980957
transform 1 0 28060 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_305
timestamp 1688980957
transform 1 0 29164 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_309
timestamp 1688980957
transform 1 0 29532 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_321
timestamp 1688980957
transform 1 0 30636 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_333
timestamp 1688980957
transform 1 0 31740 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_337
timestamp 1688980957
transform 1 0 32108 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_349
timestamp 1688980957
transform 1 0 33212 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_361
timestamp 1688980957
transform 1 0 34316 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_365
timestamp 1688980957
transform 1 0 34684 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_377
timestamp 1688980957
transform 1 0 35788 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_389
timestamp 1688980957
transform 1 0 36892 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_393
timestamp 1688980957
transform 1 0 37260 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_405
timestamp 1688980957
transform 1 0 38364 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_417
timestamp 1688980957
transform 1 0 39468 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_421
timestamp 1688980957
transform 1 0 39836 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_433
timestamp 1688980957
transform 1 0 40940 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_445
timestamp 1688980957
transform 1 0 42044 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_449
timestamp 1688980957
transform 1 0 42412 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_461
timestamp 1688980957
transform 1 0 43516 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_473
timestamp 1688980957
transform 1 0 44620 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_488
timestamp 1688980957
transform 1 0 46000 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101_500
timestamp 1688980957
transform 1 0 47104 0 -1 57664
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_505
timestamp 1688980957
transform 1 0 47564 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_517
timestamp 1688980957
transform 1 0 48668 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_529
timestamp 1688980957
transform 1 0 49772 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_533
timestamp 1688980957
transform 1 0 50140 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_545
timestamp 1688980957
transform 1 0 51244 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_557
timestamp 1688980957
transform 1 0 52348 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_561
timestamp 1688980957
transform 1 0 52716 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_573
timestamp 1688980957
transform 1 0 53820 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_585
timestamp 1688980957
transform 1 0 54924 0 -1 57664
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_589
timestamp 1688980957
transform 1 0 55292 0 -1 57664
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_101_601
timestamp 1688980957
transform 1 0 56396 0 -1 57664
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101_613
timestamp 1688980957
transform 1 0 57500 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_101_617
timestamp 1688980957
transform 1 0 57868 0 -1 57664
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 49220 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform -1 0 48576 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 48484 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform 1 0 51612 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 51060 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform 1 0 51060 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 51796 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 47932 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 48024 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 54556 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform -1 0 53820 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform -1 0 48944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 48208 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 49220 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1688980957
transform -1 0 48484 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1688980957
transform -1 0 53636 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1688980957
transform 1 0 52164 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1688980957
transform -1 0 58604 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1688980957
transform -1 0 58604 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1688980957
transform 1 0 54924 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1688980957
transform -1 0 54832 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1688980957
transform -1 0 58604 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1688980957
transform -1 0 57500 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1688980957
transform 1 0 54004 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1688980957
transform -1 0 54740 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1688980957
transform -1 0 58604 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1688980957
transform -1 0 57408 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1688980957
transform 1 0 57868 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1688980957
transform -1 0 57592 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1688980957
transform 1 0 55936 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1688980957
transform -1 0 56672 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1688980957
transform -1 0 55936 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1688980957
transform 1 0 55200 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1688980957
transform -1 0 58604 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1688980957
transform -1 0 57592 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1688980957
transform 1 0 49680 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1688980957
transform -1 0 49864 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1688980957
transform 1 0 56764 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1688980957
transform -1 0 56304 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1688980957
transform -1 0 58604 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1688980957
transform -1 0 57684 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1688980957
transform 1 0 56580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1688980957
transform -1 0 57316 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1688980957
transform 1 0 57040 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1688980957
transform -1 0 58604 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1688980957
transform -1 0 56212 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1688980957
transform -1 0 56212 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1688980957
transform -1 0 56212 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1688980957
transform -1 0 56028 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1688980957
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1688980957
transform -1 0 57500 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1688980957
transform 1 0 51428 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1688980957
transform -1 0 51612 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1688980957
transform -1 0 55936 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1688980957
transform -1 0 55752 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1688980957
transform -1 0 54280 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1688980957
transform -1 0 53452 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1688980957
transform -1 0 56120 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1688980957
transform -1 0 56028 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1688980957
transform -1 0 56028 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1688980957
transform -1 0 56028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1688980957
transform -1 0 53452 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1688980957
transform -1 0 52348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1688980957
transform 1 0 52716 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold65
timestamp 1688980957
transform -1 0 53452 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold66
timestamp 1688980957
transform 1 0 55292 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold67
timestamp 1688980957
transform -1 0 55752 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold68
timestamp 1688980957
transform 1 0 38364 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold69
timestamp 1688980957
transform -1 0 39836 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold70
timestamp 1688980957
transform -1 0 39192 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold71
timestamp 1688980957
transform -1 0 47196 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold72
timestamp 1688980957
transform -1 0 46736 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold73
timestamp 1688980957
transform 1 0 46736 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold74
timestamp 1688980957
transform 1 0 47932 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold75
timestamp 1688980957
transform -1 0 49312 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold76
timestamp 1688980957
transform 1 0 49220 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold77
timestamp 1688980957
transform 1 0 37260 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold78
timestamp 1688980957
transform -1 0 36984 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold79
timestamp 1688980957
transform -1 0 36432 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold80
timestamp 1688980957
transform -1 0 39560 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold81
timestamp 1688980957
transform -1 0 39192 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold82
timestamp 1688980957
transform -1 0 38456 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold83
timestamp 1688980957
transform -1 0 40388 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold84
timestamp 1688980957
transform 1 0 40572 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold85
timestamp 1688980957
transform 1 0 46276 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold86
timestamp 1688980957
transform -1 0 48300 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold87
timestamp 1688980957
transform -1 0 48300 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold88
timestamp 1688980957
transform -1 0 49864 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold89
timestamp 1688980957
transform -1 0 48760 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold90
timestamp 1688980957
transform -1 0 49036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold91 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 42780 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold92
timestamp 1688980957
transform -1 0 44252 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold93
timestamp 1688980957
transform -1 0 43148 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold94
timestamp 1688980957
transform 1 0 47564 0 -1 32640
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold95
timestamp 1688980957
transform 1 0 46000 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold96
timestamp 1688980957
transform 1 0 44988 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold97
timestamp 1688980957
transform -1 0 45724 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold98
timestamp 1688980957
transform 1 0 45724 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold99
timestamp 1688980957
transform -1 0 38456 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold100
timestamp 1688980957
transform -1 0 37720 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold101
timestamp 1688980957
transform -1 0 36432 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold102
timestamp 1688980957
transform -1 0 8648 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold103
timestamp 1688980957
transform -1 0 8280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold104
timestamp 1688980957
transform 1 0 6808 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold105
timestamp 1688980957
transform 1 0 46828 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold106
timestamp 1688980957
transform -1 0 46644 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold107
timestamp 1688980957
transform -1 0 46276 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold108
timestamp 1688980957
transform -1 0 4416 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold109
timestamp 1688980957
transform -1 0 4508 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold110
timestamp 1688980957
transform -1 0 3680 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold111
timestamp 1688980957
transform 1 0 49404 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold112
timestamp 1688980957
transform -1 0 48852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold113
timestamp 1688980957
transform 1 0 2668 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold114
timestamp 1688980957
transform -1 0 4508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold115
timestamp 1688980957
transform -1 0 3864 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold116
timestamp 1688980957
transform 1 0 2668 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold117
timestamp 1688980957
transform -1 0 4508 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold118
timestamp 1688980957
transform -1 0 3864 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold119
timestamp 1688980957
transform -1 0 45724 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold120
timestamp 1688980957
transform 1 0 45264 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold121
timestamp 1688980957
transform 1 0 2392 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold122
timestamp 1688980957
transform -1 0 4508 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold123
timestamp 1688980957
transform -1 0 3956 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold124
timestamp 1688980957
transform 1 0 2668 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold125
timestamp 1688980957
transform -1 0 4508 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold126
timestamp 1688980957
transform -1 0 3864 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold127
timestamp 1688980957
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold128
timestamp 1688980957
transform -1 0 3956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold129
timestamp 1688980957
transform 1 0 2760 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold130
timestamp 1688980957
transform 1 0 7544 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold131
timestamp 1688980957
transform -1 0 8832 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold132
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold133
timestamp 1688980957
transform 1 0 43424 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold134
timestamp 1688980957
transform -1 0 43148 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold135
timestamp 1688980957
transform 1 0 3220 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold136
timestamp 1688980957
transform -1 0 4508 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold137
timestamp 1688980957
transform -1 0 3680 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold138
timestamp 1688980957
transform 1 0 2852 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold139
timestamp 1688980957
transform -1 0 3956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold140
timestamp 1688980957
transform 1 0 2668 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold141
timestamp 1688980957
transform 1 0 2852 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold142
timestamp 1688980957
transform -1 0 3956 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold143
timestamp 1688980957
transform 1 0 2668 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold144
timestamp 1688980957
transform 1 0 3220 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold145
timestamp 1688980957
transform -1 0 3588 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold146
timestamp 1688980957
transform 1 0 2024 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold147
timestamp 1688980957
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold148
timestamp 1688980957
transform -1 0 3956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold149
timestamp 1688980957
transform 1 0 2668 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold150
timestamp 1688980957
transform 1 0 2852 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold151
timestamp 1688980957
transform -1 0 3772 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold152
timestamp 1688980957
transform 1 0 2300 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold153
timestamp 1688980957
transform 1 0 10120 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold154
timestamp 1688980957
transform -1 0 10764 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold155
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold156
timestamp 1688980957
transform -1 0 48300 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold157
timestamp 1688980957
transform -1 0 49312 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold158
timestamp 1688980957
transform -1 0 48024 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold159
timestamp 1688980957
transform 1 0 6532 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold160
timestamp 1688980957
transform -1 0 6900 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold161
timestamp 1688980957
transform 1 0 6900 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold162
timestamp 1688980957
transform -1 0 7084 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold163
timestamp 1688980957
transform -1 0 6256 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold164
timestamp 1688980957
transform 1 0 4784 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold165
timestamp 1688980957
transform -1 0 6440 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold166
timestamp 1688980957
transform -1 0 5428 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold167
timestamp 1688980957
transform 1 0 4508 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold168
timestamp 1688980957
transform 1 0 2208 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold169
timestamp 1688980957
transform -1 0 3680 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold170
timestamp 1688980957
transform 1 0 2668 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold171
timestamp 1688980957
transform 1 0 10212 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold172
timestamp 1688980957
transform -1 0 10856 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold173
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold174
timestamp 1688980957
transform 1 0 2852 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold175
timestamp 1688980957
transform -1 0 3680 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold176
timestamp 1688980957
transform 1 0 2208 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold177
timestamp 1688980957
transform -1 0 40204 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold178
timestamp 1688980957
transform 1 0 41308 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold179
timestamp 1688980957
transform -1 0 43148 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold180
timestamp 1688980957
transform -1 0 9568 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold181
timestamp 1688980957
transform -1 0 8832 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold182
timestamp 1688980957
transform 1 0 9384 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold183
timestamp 1688980957
transform -1 0 4600 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold184
timestamp 1688980957
transform -1 0 4784 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold185
timestamp 1688980957
transform 1 0 4600 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold186
timestamp 1688980957
transform -1 0 7912 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold187
timestamp 1688980957
transform -1 0 8648 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold188
timestamp 1688980957
transform 1 0 7636 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold189
timestamp 1688980957
transform 1 0 7176 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold190
timestamp 1688980957
transform -1 0 8464 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold191
timestamp 1688980957
transform -1 0 9016 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold192
timestamp 1688980957
transform -1 0 6256 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold193
timestamp 1688980957
transform -1 0 5520 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold194
timestamp 1688980957
transform 1 0 5244 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold195
timestamp 1688980957
transform 1 0 2852 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold196
timestamp 1688980957
transform -1 0 4232 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold197
timestamp 1688980957
transform 1 0 2760 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold198
timestamp 1688980957
transform 1 0 6624 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold199
timestamp 1688980957
transform -1 0 8188 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold200
timestamp 1688980957
transform 1 0 6992 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold201
timestamp 1688980957
transform 1 0 10120 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold202
timestamp 1688980957
transform -1 0 11224 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold203
timestamp 1688980957
transform -1 0 11592 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold204
timestamp 1688980957
transform 1 0 8280 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold205
timestamp 1688980957
transform -1 0 9752 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold206
timestamp 1688980957
transform 1 0 9384 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold207
timestamp 1688980957
transform -1 0 5520 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold208
timestamp 1688980957
transform -1 0 4784 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold209
timestamp 1688980957
transform 1 0 4508 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold210
timestamp 1688980957
transform 1 0 51152 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold211
timestamp 1688980957
transform 1 0 50140 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold212
timestamp 1688980957
transform 1 0 47840 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold213
timestamp 1688980957
transform 1 0 48484 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold214
timestamp 1688980957
transform -1 0 48484 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold215
timestamp 1688980957
transform -1 0 9660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold216
timestamp 1688980957
transform -1 0 8464 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold217
timestamp 1688980957
transform 1 0 9292 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold218
timestamp 1688980957
transform 1 0 38456 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold219
timestamp 1688980957
transform -1 0 38456 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold220
timestamp 1688980957
transform -1 0 50876 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold221
timestamp 1688980957
transform -1 0 49404 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold222
timestamp 1688980957
transform 1 0 48760 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  hold223
timestamp 1688980957
transform -1 0 49956 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold224
timestamp 1688980957
transform -1 0 49956 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold225
timestamp 1688980957
transform 1 0 50140 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold226
timestamp 1688980957
transform 1 0 43240 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold227
timestamp 1688980957
transform -1 0 43148 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold228
timestamp 1688980957
transform 1 0 42044 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold229
timestamp 1688980957
transform 1 0 43976 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  hold230 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 46276 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold231
timestamp 1688980957
transform -1 0 45724 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold232
timestamp 1688980957
transform -1 0 43516 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold233
timestamp 1688980957
transform 1 0 50140 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold234
timestamp 1688980957
transform -1 0 43148 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold235
timestamp 1688980957
transform -1 0 41768 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold236 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 43608 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold237
timestamp 1688980957
transform -1 0 44344 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold238
timestamp 1688980957
transform -1 0 42872 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold239
timestamp 1688980957
transform -1 0 50876 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold240
timestamp 1688980957
transform -1 0 42504 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold241
timestamp 1688980957
transform -1 0 42228 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold242
timestamp 1688980957
transform -1 0 50048 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold243
timestamp 1688980957
transform 1 0 44620 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_8  input1
timestamp 1688980957
transform 1 0 44988 0 -1 57664
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1688980957
transform -1 0 32844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input5
timestamp 1688980957
transform 1 0 42412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input6
timestamp 1688980957
transform 1 0 52716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform -1 0 58604 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform -1 0 58604 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1688980957
transform -1 0 58604 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform -1 0 58604 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform -1 0 57776 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform -1 0 58604 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform -1 0 58604 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 57500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform -1 0 58328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 58328 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 58052 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform -1 0 58604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 58328 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 57868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform -1 0 58144 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform -1 0 58144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 58236 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform -1 0 58052 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 58328 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 57500 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform -1 0 58144 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform -1 0 58144 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform -1 0 58604 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 58328 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 58328 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 58328 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 58328 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 58328 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 58328 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 58328 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 58328 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform -1 0 57592 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 57224 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform -1 0 58604 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform -1 0 57776 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 58328 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform -1 0 58328 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform -1 0 58604 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 58052 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 58328 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 58328 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 58328 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform 1 0 58328 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 58328 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input51
timestamp 1688980957
transform -1 0 58604 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input52
timestamp 1688980957
transform -1 0 58604 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input53
timestamp 1688980957
transform -1 0 58604 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1688980957
transform -1 0 58604 0 -1 50048
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input55
timestamp 1688980957
transform -1 0 58604 0 1 51136
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input56
timestamp 1688980957
transform -1 0 58604 0 1 52224
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input57
timestamp 1688980957
transform -1 0 58604 0 -1 53312
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1688980957
transform -1 0 58144 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1688980957
transform -1 0 58144 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1688980957
transform 1 0 57868 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform -1 0 58604 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1688980957
transform -1 0 58604 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output63 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 3680 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output64
timestamp 1688980957
transform -1 0 8832 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output65
timestamp 1688980957
transform -1 0 28980 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output66
timestamp 1688980957
transform -1 0 38916 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output67
timestamp 1688980957
transform 1 0 47564 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output68
timestamp 1688980957
transform 1 0 56304 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output69
timestamp 1688980957
transform -1 0 2852 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output70
timestamp 1688980957
transform -1 0 2852 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output71
timestamp 1688980957
transform -1 0 2852 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output72
timestamp 1688980957
transform -1 0 2852 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output73
timestamp 1688980957
transform -1 0 2852 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output74
timestamp 1688980957
transform -1 0 2852 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output75
timestamp 1688980957
transform -1 0 2852 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output76
timestamp 1688980957
transform -1 0 2852 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output77
timestamp 1688980957
transform -1 0 2852 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output78
timestamp 1688980957
transform -1 0 2852 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output79
timestamp 1688980957
transform -1 0 2852 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output80
timestamp 1688980957
transform -1 0 2852 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output81
timestamp 1688980957
transform -1 0 2852 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output82
timestamp 1688980957
transform -1 0 2852 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output83
timestamp 1688980957
transform -1 0 2852 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output84
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output85
timestamp 1688980957
transform -1 0 2852 0 1 42432
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output86
timestamp 1688980957
transform -1 0 2852 0 -1 44608
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output87
timestamp 1688980957
transform -1 0 2852 0 1 45696
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output88
timestamp 1688980957
transform -1 0 2852 0 -1 47872
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output89
timestamp 1688980957
transform -1 0 2852 0 1 48960
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output90
timestamp 1688980957
transform -1 0 2852 0 -1 51136
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output91
timestamp 1688980957
transform -1 0 2852 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output92
timestamp 1688980957
transform -1 0 2852 0 1 52224
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output93
timestamp 1688980957
transform -1 0 2852 0 -1 54400
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output94
timestamp 1688980957
transform -1 0 2852 0 1 55488
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output95
timestamp 1688980957
transform -1 0 2852 0 -1 57664
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output96
timestamp 1688980957
transform -1 0 2852 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output97
timestamp 1688980957
transform -1 0 2852 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output98
timestamp 1688980957
transform -1 0 2852 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output99
timestamp 1688980957
transform -1 0 2852 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output100
timestamp 1688980957
transform -1 0 2852 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output101
timestamp 1688980957
transform -1 0 2852 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output102
timestamp 1688980957
transform -1 0 2852 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 58880 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 58880 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 58880 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 58880 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 58880 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 58880 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 58880 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 58880 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 58880 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 58880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 58880 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 58880 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 58880 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1688980957
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1688980957
transform -1 0 58880 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1688980957
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1688980957
transform -1 0 58880 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1688980957
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1688980957
transform -1 0 58880 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1688980957
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1688980957
transform -1 0 58880 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1688980957
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1688980957
transform -1 0 58880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1688980957
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1688980957
transform -1 0 58880 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1688980957
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1688980957
transform -1 0 58880 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1688980957
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1688980957
transform -1 0 58880 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1688980957
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1688980957
transform -1 0 58880 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1688980957
transform 1 0 1104 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1688980957
transform -1 0 58880 0 -1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1688980957
transform 1 0 1104 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1688980957
transform -1 0 58880 0 1 50048
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1688980957
transform 1 0 1104 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1688980957
transform -1 0 58880 0 -1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1688980957
transform 1 0 1104 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1688980957
transform -1 0 58880 0 1 51136
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1688980957
transform 1 0 1104 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1688980957
transform -1 0 58880 0 -1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1688980957
transform 1 0 1104 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1688980957
transform -1 0 58880 0 1 52224
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1688980957
transform 1 0 1104 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1688980957
transform -1 0 58880 0 -1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1688980957
transform 1 0 1104 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1688980957
transform -1 0 58880 0 1 53312
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1688980957
transform 1 0 1104 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1688980957
transform -1 0 58880 0 -1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1688980957
transform 1 0 1104 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1688980957
transform -1 0 58880 0 1 54400
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1688980957
transform 1 0 1104 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1688980957
transform -1 0 58880 0 -1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1688980957
transform 1 0 1104 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1688980957
transform -1 0 58880 0 1 55488
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1688980957
transform 1 0 1104 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1688980957
transform -1 0 58880 0 -1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1688980957
transform 1 0 1104 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1688980957
transform -1 0 58880 0 1 56576
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1688980957
transform 1 0 1104 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1688980957
transform -1 0 58880 0 -1 57664
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  spi_mem_m_108 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17848 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1688980957
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1688980957
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1688980957
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1688980957
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1688980957
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1688980957
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1688980957
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1688980957
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1688980957
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1688980957
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1688980957
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1688980957
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1688980957
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1688980957
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1688980957
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1688980957
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1688980957
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1688980957
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1688980957
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1688980957
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1688980957
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1688980957
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1688980957
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1688980957
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1688980957
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1688980957
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1688980957
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1688980957
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1688980957
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1688980957
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1688980957
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1688980957
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1688980957
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1688980957
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1688980957
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1688980957
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1688980957
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1688980957
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1688980957
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1688980957
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1688980957
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1688980957
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1688980957
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1688980957
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1688980957
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1688980957
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1688980957
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1688980957
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1688980957
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1688980957
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1688980957
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1688980957
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1688980957
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1688980957
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1688980957
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1688980957
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1688980957
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1688980957
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1688980957
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1688980957
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1688980957
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1688980957
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1688980957
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1688980957
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1688980957
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1688980957
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1688980957
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1688980957
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1688980957
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1688980957
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1688980957
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1688980957
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1688980957
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1688980957
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1688980957
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1688980957
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1688980957
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1688980957
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1688980957
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1688980957
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1688980957
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1688980957
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1688980957
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1688980957
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1688980957
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1688980957
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1688980957
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1688980957
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1688980957
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1688980957
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1688980957
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1688980957
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1688980957
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1688980957
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1688980957
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1688980957
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1688980957
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1688980957
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1688980957
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1688980957
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1688980957
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1688980957
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1688980957
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1688980957
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1688980957
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1688980957
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1688980957
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1688980957
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1688980957
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1688980957
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1688980957
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1688980957
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1688980957
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1688980957
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1688980957
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1688980957
transform 1 0 52624 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1688980957
transform 1 0 57776 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1688980957
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1688980957
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1688980957
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1688980957
transform 1 0 50048 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1688980957
transform 1 0 55200 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1688980957
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1688980957
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1688980957
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1688980957
transform 1 0 52624 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1688980957
transform 1 0 57776 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1688980957
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1688980957
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1688980957
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1688980957
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1688980957
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1688980957
transform 1 0 50048 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1688980957
transform 1 0 55200 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_975
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_976
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_977
timestamp 1688980957
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_978
timestamp 1688980957
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_979
timestamp 1688980957
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_980
timestamp 1688980957
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_981
timestamp 1688980957
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_982
timestamp 1688980957
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_983
timestamp 1688980957
transform 1 0 52624 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_984
timestamp 1688980957
transform 1 0 57776 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_985
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_986
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_987
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_988
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_989
timestamp 1688980957
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_990
timestamp 1688980957
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_991
timestamp 1688980957
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_992
timestamp 1688980957
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_993
timestamp 1688980957
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_994
timestamp 1688980957
transform 1 0 50048 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_995
timestamp 1688980957
transform 1 0 55200 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_996
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_997
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_998
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_999
timestamp 1688980957
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1000
timestamp 1688980957
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1001
timestamp 1688980957
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1002
timestamp 1688980957
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1003
timestamp 1688980957
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1004
timestamp 1688980957
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1005
timestamp 1688980957
transform 1 0 52624 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1006
timestamp 1688980957
transform 1 0 57776 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1007
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1008
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1009
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1010
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1011
timestamp 1688980957
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1012
timestamp 1688980957
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1013
timestamp 1688980957
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1014
timestamp 1688980957
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1015
timestamp 1688980957
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1016
timestamp 1688980957
transform 1 0 50048 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1017
timestamp 1688980957
transform 1 0 55200 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1018
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1019
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1020
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1021
timestamp 1688980957
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1022
timestamp 1688980957
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1023
timestamp 1688980957
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1024
timestamp 1688980957
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1025
timestamp 1688980957
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1026
timestamp 1688980957
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1027
timestamp 1688980957
transform 1 0 52624 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1028
timestamp 1688980957
transform 1 0 57776 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1029
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1030
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1031
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1032
timestamp 1688980957
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1033
timestamp 1688980957
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1034
timestamp 1688980957
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1035
timestamp 1688980957
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1036
timestamp 1688980957
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1037
timestamp 1688980957
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1038
timestamp 1688980957
transform 1 0 50048 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1039
timestamp 1688980957
transform 1 0 55200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1040
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1041
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1042
timestamp 1688980957
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1043
timestamp 1688980957
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1044
timestamp 1688980957
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1045
timestamp 1688980957
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1046
timestamp 1688980957
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1047
timestamp 1688980957
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1048
timestamp 1688980957
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1049
timestamp 1688980957
transform 1 0 52624 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1050
timestamp 1688980957
transform 1 0 57776 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1051
timestamp 1688980957
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1052
timestamp 1688980957
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1053
timestamp 1688980957
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1054
timestamp 1688980957
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1055
timestamp 1688980957
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1056
timestamp 1688980957
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1057
timestamp 1688980957
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1058
timestamp 1688980957
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1059
timestamp 1688980957
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1060
timestamp 1688980957
transform 1 0 50048 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1061
timestamp 1688980957
transform 1 0 55200 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1062
timestamp 1688980957
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1063
timestamp 1688980957
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1064
timestamp 1688980957
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1065
timestamp 1688980957
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1066
timestamp 1688980957
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1067
timestamp 1688980957
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1068
timestamp 1688980957
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1069
timestamp 1688980957
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1070
timestamp 1688980957
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1071
timestamp 1688980957
transform 1 0 52624 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1072
timestamp 1688980957
transform 1 0 57776 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1073
timestamp 1688980957
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1074
timestamp 1688980957
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1075
timestamp 1688980957
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1076
timestamp 1688980957
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1077
timestamp 1688980957
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1078
timestamp 1688980957
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1079
timestamp 1688980957
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1080
timestamp 1688980957
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1081
timestamp 1688980957
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1082
timestamp 1688980957
transform 1 0 50048 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1083
timestamp 1688980957
transform 1 0 55200 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1084
timestamp 1688980957
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1085
timestamp 1688980957
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1086
timestamp 1688980957
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1087
timestamp 1688980957
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1088
timestamp 1688980957
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1089
timestamp 1688980957
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1090
timestamp 1688980957
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1091
timestamp 1688980957
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1092
timestamp 1688980957
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1093
timestamp 1688980957
transform 1 0 52624 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1094
timestamp 1688980957
transform 1 0 57776 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1095
timestamp 1688980957
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1096
timestamp 1688980957
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1097
timestamp 1688980957
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1098
timestamp 1688980957
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1099
timestamp 1688980957
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1100
timestamp 1688980957
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1101
timestamp 1688980957
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1102
timestamp 1688980957
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1103
timestamp 1688980957
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1104
timestamp 1688980957
transform 1 0 50048 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1105
timestamp 1688980957
transform 1 0 55200 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1106
timestamp 1688980957
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1107
timestamp 1688980957
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1108
timestamp 1688980957
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1109
timestamp 1688980957
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1110
timestamp 1688980957
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1111
timestamp 1688980957
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1112
timestamp 1688980957
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1113
timestamp 1688980957
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1114
timestamp 1688980957
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1115
timestamp 1688980957
transform 1 0 52624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1116
timestamp 1688980957
transform 1 0 57776 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1117
timestamp 1688980957
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1118
timestamp 1688980957
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1119
timestamp 1688980957
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1120
timestamp 1688980957
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1121
timestamp 1688980957
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1122
timestamp 1688980957
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1123
timestamp 1688980957
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1124
timestamp 1688980957
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1125
timestamp 1688980957
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1126
timestamp 1688980957
transform 1 0 50048 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1127
timestamp 1688980957
transform 1 0 55200 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1128
timestamp 1688980957
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1129
timestamp 1688980957
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1130
timestamp 1688980957
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1131
timestamp 1688980957
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1132
timestamp 1688980957
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1133
timestamp 1688980957
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1134
timestamp 1688980957
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1135
timestamp 1688980957
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1136
timestamp 1688980957
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1137
timestamp 1688980957
transform 1 0 52624 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1138
timestamp 1688980957
transform 1 0 57776 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1139
timestamp 1688980957
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1140
timestamp 1688980957
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1141
timestamp 1688980957
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1142
timestamp 1688980957
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1143
timestamp 1688980957
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1144
timestamp 1688980957
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1145
timestamp 1688980957
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1146
timestamp 1688980957
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1147
timestamp 1688980957
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1148
timestamp 1688980957
transform 1 0 50048 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1149
timestamp 1688980957
transform 1 0 55200 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1150
timestamp 1688980957
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1151
timestamp 1688980957
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1152
timestamp 1688980957
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1153
timestamp 1688980957
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1154
timestamp 1688980957
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1155
timestamp 1688980957
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1156
timestamp 1688980957
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1157
timestamp 1688980957
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1158
timestamp 1688980957
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1159
timestamp 1688980957
transform 1 0 52624 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1160
timestamp 1688980957
transform 1 0 57776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1161
timestamp 1688980957
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1162
timestamp 1688980957
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1163
timestamp 1688980957
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1164
timestamp 1688980957
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1165
timestamp 1688980957
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1166
timestamp 1688980957
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1167
timestamp 1688980957
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1168
timestamp 1688980957
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1169
timestamp 1688980957
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1170
timestamp 1688980957
transform 1 0 50048 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1171
timestamp 1688980957
transform 1 0 55200 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1172
timestamp 1688980957
transform 1 0 6256 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1173
timestamp 1688980957
transform 1 0 11408 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1174
timestamp 1688980957
transform 1 0 16560 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1175
timestamp 1688980957
transform 1 0 21712 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1176
timestamp 1688980957
transform 1 0 26864 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1177
timestamp 1688980957
transform 1 0 32016 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1178
timestamp 1688980957
transform 1 0 37168 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1179
timestamp 1688980957
transform 1 0 42320 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1180
timestamp 1688980957
transform 1 0 47472 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1181
timestamp 1688980957
transform 1 0 52624 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1182
timestamp 1688980957
transform 1 0 57776 0 -1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1183
timestamp 1688980957
transform 1 0 3680 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1184
timestamp 1688980957
transform 1 0 8832 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1185
timestamp 1688980957
transform 1 0 13984 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1186
timestamp 1688980957
transform 1 0 19136 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1187
timestamp 1688980957
transform 1 0 24288 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1188
timestamp 1688980957
transform 1 0 29440 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1189
timestamp 1688980957
transform 1 0 34592 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1190
timestamp 1688980957
transform 1 0 39744 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1191
timestamp 1688980957
transform 1 0 44896 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1192
timestamp 1688980957
transform 1 0 50048 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1193
timestamp 1688980957
transform 1 0 55200 0 1 50048
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1194
timestamp 1688980957
transform 1 0 6256 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1195
timestamp 1688980957
transform 1 0 11408 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1196
timestamp 1688980957
transform 1 0 16560 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1197
timestamp 1688980957
transform 1 0 21712 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1198
timestamp 1688980957
transform 1 0 26864 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1199
timestamp 1688980957
transform 1 0 32016 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1200
timestamp 1688980957
transform 1 0 37168 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1201
timestamp 1688980957
transform 1 0 42320 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1202
timestamp 1688980957
transform 1 0 47472 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1203
timestamp 1688980957
transform 1 0 52624 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1204
timestamp 1688980957
transform 1 0 57776 0 -1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1205
timestamp 1688980957
transform 1 0 3680 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1206
timestamp 1688980957
transform 1 0 8832 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1207
timestamp 1688980957
transform 1 0 13984 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1208
timestamp 1688980957
transform 1 0 19136 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1209
timestamp 1688980957
transform 1 0 24288 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1210
timestamp 1688980957
transform 1 0 29440 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1211
timestamp 1688980957
transform 1 0 34592 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1212
timestamp 1688980957
transform 1 0 39744 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1213
timestamp 1688980957
transform 1 0 44896 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1214
timestamp 1688980957
transform 1 0 50048 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1215
timestamp 1688980957
transform 1 0 55200 0 1 51136
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1216
timestamp 1688980957
transform 1 0 6256 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1217
timestamp 1688980957
transform 1 0 11408 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1218
timestamp 1688980957
transform 1 0 16560 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1219
timestamp 1688980957
transform 1 0 21712 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1220
timestamp 1688980957
transform 1 0 26864 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1221
timestamp 1688980957
transform 1 0 32016 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1222
timestamp 1688980957
transform 1 0 37168 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1223
timestamp 1688980957
transform 1 0 42320 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1224
timestamp 1688980957
transform 1 0 47472 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1225
timestamp 1688980957
transform 1 0 52624 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1226
timestamp 1688980957
transform 1 0 57776 0 -1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1227
timestamp 1688980957
transform 1 0 3680 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1228
timestamp 1688980957
transform 1 0 8832 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1229
timestamp 1688980957
transform 1 0 13984 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1230
timestamp 1688980957
transform 1 0 19136 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1231
timestamp 1688980957
transform 1 0 24288 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1232
timestamp 1688980957
transform 1 0 29440 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1233
timestamp 1688980957
transform 1 0 34592 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1234
timestamp 1688980957
transform 1 0 39744 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1235
timestamp 1688980957
transform 1 0 44896 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1236
timestamp 1688980957
transform 1 0 50048 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1237
timestamp 1688980957
transform 1 0 55200 0 1 52224
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1238
timestamp 1688980957
transform 1 0 6256 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1239
timestamp 1688980957
transform 1 0 11408 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1240
timestamp 1688980957
transform 1 0 16560 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1241
timestamp 1688980957
transform 1 0 21712 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1242
timestamp 1688980957
transform 1 0 26864 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1243
timestamp 1688980957
transform 1 0 32016 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1244
timestamp 1688980957
transform 1 0 37168 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1245
timestamp 1688980957
transform 1 0 42320 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1246
timestamp 1688980957
transform 1 0 47472 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1247
timestamp 1688980957
transform 1 0 52624 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1248
timestamp 1688980957
transform 1 0 57776 0 -1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1249
timestamp 1688980957
transform 1 0 3680 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1250
timestamp 1688980957
transform 1 0 8832 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1251
timestamp 1688980957
transform 1 0 13984 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1252
timestamp 1688980957
transform 1 0 19136 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1253
timestamp 1688980957
transform 1 0 24288 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1254
timestamp 1688980957
transform 1 0 29440 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1255
timestamp 1688980957
transform 1 0 34592 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1256
timestamp 1688980957
transform 1 0 39744 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1257
timestamp 1688980957
transform 1 0 44896 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1258
timestamp 1688980957
transform 1 0 50048 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1259
timestamp 1688980957
transform 1 0 55200 0 1 53312
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1260
timestamp 1688980957
transform 1 0 6256 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1261
timestamp 1688980957
transform 1 0 11408 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1262
timestamp 1688980957
transform 1 0 16560 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1263
timestamp 1688980957
transform 1 0 21712 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1264
timestamp 1688980957
transform 1 0 26864 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1265
timestamp 1688980957
transform 1 0 32016 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1266
timestamp 1688980957
transform 1 0 37168 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1267
timestamp 1688980957
transform 1 0 42320 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1268
timestamp 1688980957
transform 1 0 47472 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1269
timestamp 1688980957
transform 1 0 52624 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1270
timestamp 1688980957
transform 1 0 57776 0 -1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1271
timestamp 1688980957
transform 1 0 3680 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1272
timestamp 1688980957
transform 1 0 8832 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1273
timestamp 1688980957
transform 1 0 13984 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1274
timestamp 1688980957
transform 1 0 19136 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1275
timestamp 1688980957
transform 1 0 24288 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1276
timestamp 1688980957
transform 1 0 29440 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1277
timestamp 1688980957
transform 1 0 34592 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1278
timestamp 1688980957
transform 1 0 39744 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1279
timestamp 1688980957
transform 1 0 44896 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1280
timestamp 1688980957
transform 1 0 50048 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1281
timestamp 1688980957
transform 1 0 55200 0 1 54400
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1282
timestamp 1688980957
transform 1 0 6256 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1283
timestamp 1688980957
transform 1 0 11408 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1284
timestamp 1688980957
transform 1 0 16560 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1285
timestamp 1688980957
transform 1 0 21712 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1286
timestamp 1688980957
transform 1 0 26864 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1287
timestamp 1688980957
transform 1 0 32016 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1288
timestamp 1688980957
transform 1 0 37168 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1289
timestamp 1688980957
transform 1 0 42320 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1290
timestamp 1688980957
transform 1 0 47472 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1291
timestamp 1688980957
transform 1 0 52624 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1292
timestamp 1688980957
transform 1 0 57776 0 -1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1293
timestamp 1688980957
transform 1 0 3680 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1294
timestamp 1688980957
transform 1 0 8832 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1295
timestamp 1688980957
transform 1 0 13984 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1296
timestamp 1688980957
transform 1 0 19136 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1297
timestamp 1688980957
transform 1 0 24288 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1298
timestamp 1688980957
transform 1 0 29440 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1299
timestamp 1688980957
transform 1 0 34592 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1300
timestamp 1688980957
transform 1 0 39744 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1301
timestamp 1688980957
transform 1 0 44896 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1302
timestamp 1688980957
transform 1 0 50048 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1303
timestamp 1688980957
transform 1 0 55200 0 1 55488
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1304
timestamp 1688980957
transform 1 0 6256 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1305
timestamp 1688980957
transform 1 0 11408 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1306
timestamp 1688980957
transform 1 0 16560 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1307
timestamp 1688980957
transform 1 0 21712 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1308
timestamp 1688980957
transform 1 0 26864 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1309
timestamp 1688980957
transform 1 0 32016 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1310
timestamp 1688980957
transform 1 0 37168 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1311
timestamp 1688980957
transform 1 0 42320 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1312
timestamp 1688980957
transform 1 0 47472 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1313
timestamp 1688980957
transform 1 0 52624 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1314
timestamp 1688980957
transform 1 0 57776 0 -1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1315
timestamp 1688980957
transform 1 0 3680 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1316
timestamp 1688980957
transform 1 0 8832 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1317
timestamp 1688980957
transform 1 0 13984 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1318
timestamp 1688980957
transform 1 0 19136 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1319
timestamp 1688980957
transform 1 0 24288 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1320
timestamp 1688980957
transform 1 0 29440 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1321
timestamp 1688980957
transform 1 0 34592 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1322
timestamp 1688980957
transform 1 0 39744 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1323
timestamp 1688980957
transform 1 0 44896 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1324
timestamp 1688980957
transform 1 0 50048 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1325
timestamp 1688980957
transform 1 0 55200 0 1 56576
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1326
timestamp 1688980957
transform 1 0 3680 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1327
timestamp 1688980957
transform 1 0 6256 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1328
timestamp 1688980957
transform 1 0 8832 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1329
timestamp 1688980957
transform 1 0 11408 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1330
timestamp 1688980957
transform 1 0 13984 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1331
timestamp 1688980957
transform 1 0 16560 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1332
timestamp 1688980957
transform 1 0 19136 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1333
timestamp 1688980957
transform 1 0 21712 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1334
timestamp 1688980957
transform 1 0 24288 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1335
timestamp 1688980957
transform 1 0 26864 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1336
timestamp 1688980957
transform 1 0 29440 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1337
timestamp 1688980957
transform 1 0 32016 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1338
timestamp 1688980957
transform 1 0 34592 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1339
timestamp 1688980957
transform 1 0 37168 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1340
timestamp 1688980957
transform 1 0 39744 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1341
timestamp 1688980957
transform 1 0 42320 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1342
timestamp 1688980957
transform 1 0 44896 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1343
timestamp 1688980957
transform 1 0 47472 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1344
timestamp 1688980957
transform 1 0 50048 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1345
timestamp 1688980957
transform 1 0 52624 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1346
timestamp 1688980957
transform 1 0 55200 0 -1 57664
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_1347
timestamp 1688980957
transform 1 0 57776 0 -1 57664
box -38 -48 130 592
<< labels >>
flabel metal2 s 14922 59200 14978 60000 0 FreeSans 224 90 0 0 clk_i
port 0 nsew signal input
flabel metal2 s 44914 59200 44970 60000 0 FreeSans 224 90 0 0 nrst_i
port 1 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 spi_clk_o
port 2 nsew signal tristate
flabel metal2 s 7562 0 7618 800 0 FreeSans 224 90 0 0 spi_cs_o
port 3 nsew signal tristate
flabel metal2 s 12530 0 12586 800 0 FreeSans 224 90 0 0 spi_dqsm_i
port 4 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 spi_dqsm_o
port 5 nsew signal tristate
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 spi_miso_i[0]
port 6 nsew signal input
flabel metal2 s 32402 0 32458 800 0 FreeSans 224 90 0 0 spi_miso_i[1]
port 7 nsew signal input
flabel metal2 s 42338 0 42394 800 0 FreeSans 224 90 0 0 spi_miso_i[2]
port 8 nsew signal input
flabel metal2 s 52274 0 52330 800 0 FreeSans 224 90 0 0 spi_miso_i[3]
port 9 nsew signal input
flabel metal2 s 27434 0 27490 800 0 FreeSans 224 90 0 0 spi_mosi_o[0]
port 10 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 spi_mosi_o[1]
port 11 nsew signal tristate
flabel metal2 s 47306 0 47362 800 0 FreeSans 224 90 0 0 spi_mosi_o[2]
port 12 nsew signal tristate
flabel metal2 s 57242 0 57298 800 0 FreeSans 224 90 0 0 spi_mosi_o[3]
port 13 nsew signal tristate
flabel metal3 s 59200 7080 60000 7200 0 FreeSans 480 0 0 0 sport_i[0]
port 14 nsew signal input
flabel metal3 s 59200 15240 60000 15360 0 FreeSans 480 0 0 0 sport_i[10]
port 15 nsew signal input
flabel metal3 s 59200 16056 60000 16176 0 FreeSans 480 0 0 0 sport_i[11]
port 16 nsew signal input
flabel metal3 s 59200 16872 60000 16992 0 FreeSans 480 0 0 0 sport_i[12]
port 17 nsew signal input
flabel metal3 s 59200 17688 60000 17808 0 FreeSans 480 0 0 0 sport_i[13]
port 18 nsew signal input
flabel metal3 s 59200 18504 60000 18624 0 FreeSans 480 0 0 0 sport_i[14]
port 19 nsew signal input
flabel metal3 s 59200 19320 60000 19440 0 FreeSans 480 0 0 0 sport_i[15]
port 20 nsew signal input
flabel metal3 s 59200 20136 60000 20256 0 FreeSans 480 0 0 0 sport_i[16]
port 21 nsew signal input
flabel metal3 s 59200 20952 60000 21072 0 FreeSans 480 0 0 0 sport_i[17]
port 22 nsew signal input
flabel metal3 s 59200 21768 60000 21888 0 FreeSans 480 0 0 0 sport_i[18]
port 23 nsew signal input
flabel metal3 s 59200 22584 60000 22704 0 FreeSans 480 0 0 0 sport_i[19]
port 24 nsew signal input
flabel metal3 s 59200 7896 60000 8016 0 FreeSans 480 0 0 0 sport_i[1]
port 25 nsew signal input
flabel metal3 s 59200 23400 60000 23520 0 FreeSans 480 0 0 0 sport_i[20]
port 26 nsew signal input
flabel metal3 s 59200 24216 60000 24336 0 FreeSans 480 0 0 0 sport_i[21]
port 27 nsew signal input
flabel metal3 s 59200 25032 60000 25152 0 FreeSans 480 0 0 0 sport_i[22]
port 28 nsew signal input
flabel metal3 s 59200 25848 60000 25968 0 FreeSans 480 0 0 0 sport_i[23]
port 29 nsew signal input
flabel metal3 s 59200 26664 60000 26784 0 FreeSans 480 0 0 0 sport_i[24]
port 30 nsew signal input
flabel metal3 s 59200 27480 60000 27600 0 FreeSans 480 0 0 0 sport_i[25]
port 31 nsew signal input
flabel metal3 s 59200 28296 60000 28416 0 FreeSans 480 0 0 0 sport_i[26]
port 32 nsew signal input
flabel metal3 s 59200 29112 60000 29232 0 FreeSans 480 0 0 0 sport_i[27]
port 33 nsew signal input
flabel metal3 s 59200 29928 60000 30048 0 FreeSans 480 0 0 0 sport_i[28]
port 34 nsew signal input
flabel metal3 s 59200 30744 60000 30864 0 FreeSans 480 0 0 0 sport_i[29]
port 35 nsew signal input
flabel metal3 s 59200 8712 60000 8832 0 FreeSans 480 0 0 0 sport_i[2]
port 36 nsew signal input
flabel metal3 s 59200 31560 60000 31680 0 FreeSans 480 0 0 0 sport_i[30]
port 37 nsew signal input
flabel metal3 s 59200 32376 60000 32496 0 FreeSans 480 0 0 0 sport_i[31]
port 38 nsew signal input
flabel metal3 s 59200 33192 60000 33312 0 FreeSans 480 0 0 0 sport_i[32]
port 39 nsew signal input
flabel metal3 s 59200 34008 60000 34128 0 FreeSans 480 0 0 0 sport_i[33]
port 40 nsew signal input
flabel metal3 s 59200 34824 60000 34944 0 FreeSans 480 0 0 0 sport_i[34]
port 41 nsew signal input
flabel metal3 s 59200 35640 60000 35760 0 FreeSans 480 0 0 0 sport_i[35]
port 42 nsew signal input
flabel metal3 s 59200 36456 60000 36576 0 FreeSans 480 0 0 0 sport_i[36]
port 43 nsew signal input
flabel metal3 s 59200 37272 60000 37392 0 FreeSans 480 0 0 0 sport_i[37]
port 44 nsew signal input
flabel metal3 s 59200 38088 60000 38208 0 FreeSans 480 0 0 0 sport_i[38]
port 45 nsew signal input
flabel metal3 s 59200 38904 60000 39024 0 FreeSans 480 0 0 0 sport_i[39]
port 46 nsew signal input
flabel metal3 s 59200 9528 60000 9648 0 FreeSans 480 0 0 0 sport_i[3]
port 47 nsew signal input
flabel metal3 s 59200 39720 60000 39840 0 FreeSans 480 0 0 0 sport_i[40]
port 48 nsew signal input
flabel metal3 s 59200 40536 60000 40656 0 FreeSans 480 0 0 0 sport_i[41]
port 49 nsew signal input
flabel metal3 s 59200 41352 60000 41472 0 FreeSans 480 0 0 0 sport_i[42]
port 50 nsew signal input
flabel metal3 s 59200 42168 60000 42288 0 FreeSans 480 0 0 0 sport_i[43]
port 51 nsew signal input
flabel metal3 s 59200 42984 60000 43104 0 FreeSans 480 0 0 0 sport_i[44]
port 52 nsew signal input
flabel metal3 s 59200 43800 60000 43920 0 FreeSans 480 0 0 0 sport_i[45]
port 53 nsew signal input
flabel metal3 s 59200 44616 60000 44736 0 FreeSans 480 0 0 0 sport_i[46]
port 54 nsew signal input
flabel metal3 s 59200 45432 60000 45552 0 FreeSans 480 0 0 0 sport_i[47]
port 55 nsew signal input
flabel metal3 s 59200 46248 60000 46368 0 FreeSans 480 0 0 0 sport_i[48]
port 56 nsew signal input
flabel metal3 s 59200 47064 60000 47184 0 FreeSans 480 0 0 0 sport_i[49]
port 57 nsew signal input
flabel metal3 s 59200 10344 60000 10464 0 FreeSans 480 0 0 0 sport_i[4]
port 58 nsew signal input
flabel metal3 s 59200 47880 60000 48000 0 FreeSans 480 0 0 0 sport_i[50]
port 59 nsew signal input
flabel metal3 s 59200 48696 60000 48816 0 FreeSans 480 0 0 0 sport_i[51]
port 60 nsew signal input
flabel metal3 s 59200 49512 60000 49632 0 FreeSans 480 0 0 0 sport_i[52]
port 61 nsew signal input
flabel metal3 s 59200 50328 60000 50448 0 FreeSans 480 0 0 0 sport_i[53]
port 62 nsew signal input
flabel metal3 s 59200 51144 60000 51264 0 FreeSans 480 0 0 0 sport_i[54]
port 63 nsew signal input
flabel metal3 s 59200 51960 60000 52080 0 FreeSans 480 0 0 0 sport_i[55]
port 64 nsew signal input
flabel metal3 s 59200 52776 60000 52896 0 FreeSans 480 0 0 0 sport_i[56]
port 65 nsew signal input
flabel metal3 s 59200 11160 60000 11280 0 FreeSans 480 0 0 0 sport_i[5]
port 66 nsew signal input
flabel metal3 s 59200 11976 60000 12096 0 FreeSans 480 0 0 0 sport_i[6]
port 67 nsew signal input
flabel metal3 s 59200 12792 60000 12912 0 FreeSans 480 0 0 0 sport_i[7]
port 68 nsew signal input
flabel metal3 s 59200 13608 60000 13728 0 FreeSans 480 0 0 0 sport_i[8]
port 69 nsew signal input
flabel metal3 s 59200 14424 60000 14544 0 FreeSans 480 0 0 0 sport_i[9]
port 70 nsew signal input
flabel metal3 s 0 3000 800 3120 0 FreeSans 480 0 0 0 sport_o[0]
port 71 nsew signal tristate
flabel metal3 s 0 19320 800 19440 0 FreeSans 480 0 0 0 sport_o[10]
port 72 nsew signal tristate
flabel metal3 s 0 20952 800 21072 0 FreeSans 480 0 0 0 sport_o[11]
port 73 nsew signal tristate
flabel metal3 s 0 22584 800 22704 0 FreeSans 480 0 0 0 sport_o[12]
port 74 nsew signal tristate
flabel metal3 s 0 24216 800 24336 0 FreeSans 480 0 0 0 sport_o[13]
port 75 nsew signal tristate
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 sport_o[14]
port 76 nsew signal tristate
flabel metal3 s 0 27480 800 27600 0 FreeSans 480 0 0 0 sport_o[15]
port 77 nsew signal tristate
flabel metal3 s 0 29112 800 29232 0 FreeSans 480 0 0 0 sport_o[16]
port 78 nsew signal tristate
flabel metal3 s 0 30744 800 30864 0 FreeSans 480 0 0 0 sport_o[17]
port 79 nsew signal tristate
flabel metal3 s 0 32376 800 32496 0 FreeSans 480 0 0 0 sport_o[18]
port 80 nsew signal tristate
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 sport_o[19]
port 81 nsew signal tristate
flabel metal3 s 0 4632 800 4752 0 FreeSans 480 0 0 0 sport_o[1]
port 82 nsew signal tristate
flabel metal3 s 0 35640 800 35760 0 FreeSans 480 0 0 0 sport_o[20]
port 83 nsew signal tristate
flabel metal3 s 0 37272 800 37392 0 FreeSans 480 0 0 0 sport_o[21]
port 84 nsew signal tristate
flabel metal3 s 0 38904 800 39024 0 FreeSans 480 0 0 0 sport_o[22]
port 85 nsew signal tristate
flabel metal3 s 0 40536 800 40656 0 FreeSans 480 0 0 0 sport_o[23]
port 86 nsew signal tristate
flabel metal3 s 0 42168 800 42288 0 FreeSans 480 0 0 0 sport_o[24]
port 87 nsew signal tristate
flabel metal3 s 0 43800 800 43920 0 FreeSans 480 0 0 0 sport_o[25]
port 88 nsew signal tristate
flabel metal3 s 0 45432 800 45552 0 FreeSans 480 0 0 0 sport_o[26]
port 89 nsew signal tristate
flabel metal3 s 0 47064 800 47184 0 FreeSans 480 0 0 0 sport_o[27]
port 90 nsew signal tristate
flabel metal3 s 0 48696 800 48816 0 FreeSans 480 0 0 0 sport_o[28]
port 91 nsew signal tristate
flabel metal3 s 0 50328 800 50448 0 FreeSans 480 0 0 0 sport_o[29]
port 92 nsew signal tristate
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 sport_o[2]
port 93 nsew signal tristate
flabel metal3 s 0 51960 800 52080 0 FreeSans 480 0 0 0 sport_o[30]
port 94 nsew signal tristate
flabel metal3 s 0 53592 800 53712 0 FreeSans 480 0 0 0 sport_o[31]
port 95 nsew signal tristate
flabel metal3 s 0 55224 800 55344 0 FreeSans 480 0 0 0 sport_o[32]
port 96 nsew signal tristate
flabel metal3 s 0 56856 800 56976 0 FreeSans 480 0 0 0 sport_o[33]
port 97 nsew signal tristate
flabel metal3 s 0 7896 800 8016 0 FreeSans 480 0 0 0 sport_o[3]
port 98 nsew signal tristate
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 sport_o[4]
port 99 nsew signal tristate
flabel metal3 s 0 11160 800 11280 0 FreeSans 480 0 0 0 sport_o[5]
port 100 nsew signal tristate
flabel metal3 s 0 12792 800 12912 0 FreeSans 480 0 0 0 sport_o[6]
port 101 nsew signal tristate
flabel metal3 s 0 14424 800 14544 0 FreeSans 480 0 0 0 sport_o[7]
port 102 nsew signal tristate
flabel metal3 s 0 16056 800 16176 0 FreeSans 480 0 0 0 sport_o[8]
port 103 nsew signal tristate
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 sport_o[9]
port 104 nsew signal tristate
flabel metal4 s 4208 2128 4528 57712 0 FreeSans 1920 90 0 0 vccd1
port 105 nsew power bidirectional
flabel metal4 s 34928 2128 35248 57712 0 FreeSans 1920 90 0 0 vccd1
port 105 nsew power bidirectional
flabel metal4 s 19568 2128 19888 57712 0 FreeSans 1920 90 0 0 vssd1
port 106 nsew ground bidirectional
flabel metal4 s 50288 2128 50608 57712 0 FreeSans 1920 90 0 0 vssd1
port 106 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 60000 60000
<< end >>
