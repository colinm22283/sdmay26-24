module word_stripe_cache_m #(
    parameter STRIPE_SIZE = 8
) (
    input wire clk_i,
    input wire nrst_i,

    input  wire [`BUS_MOPORT] cached_mport_i,
    output reg  [`BUS_MIPORT] cached_mport_o,

    input  wire [`BUS_MIPORT] mport_i,
    output reg  [`BUS_MOPORT] mport_o
);

    localparam STATE_READY       = 3'b000;
    localparam STATE_WRITE       = 3'b001;
    localparam STATE_WRITE_FLUSH = 3'b010;
    localparam STATE_READ        = 3'b011;
    localparam STATE_READ_FLUSH  = 3'b100;
    localparam STATE_DONE = 3'b011;

    localparam STATE_PASSTHROUGH = 3'b111;

    reg [2:0] state;

    reg [`BUS_ADDR_PORT] write_stripe_addr;
    reg [$clog2(STRIPE_SIZE + 1) - 1:0] write_stripe_size;
    reg [31:0] write_stripe [STRIPE_SIZE - 1:0];

    reg [$clog2(STRIPE_SIZE + 1) - 1:0] write_stripe_index;
    reg [1:0] write_stripe_state;

    reg [`BUS_ADDR_PORT] read_stripe_addr;
    reg [$clog2(STRIPE_SIZE + 1) - 1:0] read_stripe_size;
    reg [31:0] read_stripe [STRIPE_SIZE - 1:0];

    reg [$clog2(STRIPE_SIZE + 1) - 1:0] read_stripe_index;
    reg [1:0] read_stripe_state;

    always @(posedge clk_i, negedge nrst_i) begin
        if (!nrst_i) begin
            state <= STATE_READY;

            cached_mport_o <= 0;

            write_stripe_addr  <= 0;
            write_stripe_size  <= 0;

            write_stripe_index <= 0;
            write_stripe_state <= 0;
        end
        else if (clk_i) begin
            case (state)
                STATE_READY: begin
                    if (write_stripe_size == STRIPE_SIZE) begin
                        state <= STATE_WRITE_FLUSH;
                                    
                        write_stripe_index <= 0;
                    end
                    else begin
                        if (cached_mport_i[`BUS_MO_REQ]) begin
                            if (cached_mport_i[`BUS_MO_RW] == `BUS_READ) begin
                                if (cached_mport_i[`BUS_MO_SIZE] != `BUS_SIZE_WORD) begin
                                    state <= STATE_PASSTHROUGH;
                                end
                                else begin
                                    if (
                                        cached_mport_i[`BUS_MO_ADDR] != read_stripe_addr + (write_stripe_size * 4) &&
                                        write_stripe_size != 0
                                    ) begin
                                        state <= STATE_WRITE_FLUSH;
                                        
                                        write_stripe_index <= 0;
                                    end
                                    else begin
                                        state <= STATE_WRITE;

                                        if (write_stripe_size == 0) write_stripe_addr <= cached_mport_i[`BUS_MO_ADDR];

                                        cached_mport_o[`BUS_MI_ACK] <= 1;
                                    end
                                end
                            end
                            else begin
                                if (cached_mport_i[`BUS_MO_SIZE] != `BUS_SIZE_WORD) begin
                                    state <= STATE_PASSTHROUGH;
                                end
                                else begin
                                    if (
                                        cached_mport_i[`BUS_MO_ADDR] != write_stripe_addr + (write_stripe_size * 4) &&
                                        write_stripe_size != 0
                                    ) begin
                                        state <= STATE_WRITE_FLUSH;
                                        
                                        write_stripe_index <= 0;
                                    end
                                    else begin
                                        state <= STATE_WRITE;

                                        if (write_stripe_size == 0) write_stripe_addr <= cached_mport_i[`BUS_MO_ADDR];

                                        cached_mport_o[`BUS_MI_ACK] <= 1;
                                    end
                                end
                            end
                        end
                    end
                end

                STATE_WRITE: begin
                    state <= STATE_DONE;

                    write_stripe[write_stripe_size] <= cached_mport_i[`BUS_MO_DATA];

                    write_stripe_size <= write_stripe_size + 1;
                end

                STATE_WRITE_FLUSH: begin
                    case (write_stripe_state)
                        0: begin
                            if (mport_i[`BUS_MI_ACK]) begin
                                write_stripe_state <= 1;

                                write_stripe_index <= write_stripe_index + 1;
                            end

                            mport_o[`BUS_MO_ADDR] <= write_stripe_addr;
                            mport_o[`BUS_MO_DATA] <= write_stripe[write_stripe_index];
                            mport_o[`BUS_MO_RW]   <= `BUS_WRITE;
                            mport_o[`BUS_MO_SIZE] <= `BUS_SIZE_STREAM;

                            mport_o[`BUS_MO_REQ] <= 1;
                        end

                        1: begin
                            if (mport_i[`BUS_MI_SEQSLV]) begin
                                if (write_stripe_index == write_stripe_size) begin
                                    write_stripe_state <= 3;
                                end
                                else begin
                                    write_stripe_state <= 2;

                                    $display("Attempt write 0x%h", write_stripe[write_stripe_index]);
                                    mport_o[`BUS_MO_DATA] <= write_stripe[write_stripe_index];
                                end
                            end
                        end

                        2: begin
                            write_stripe_state <= 1;

                            write_stripe_index <= write_stripe_index + 1;
                        end

                        3: begin
                            if (!mport_i[`BUS_MI_ACK]) begin
                                state <= STATE_READY;
                                write_stripe_state <= 0;
                            end

                            mport_o[`BUS_MO_REQ] <= 0;

                            write_stripe_size <= 0;
                        end
                    endcase
                end

                STATE_DONE: begin
                    if (!cached_mport_i[`BUS_MO_REQ]) state <= STATE_READY;

                    cached_mport_o[`BUS_MI_ACK] <= 0;
                end

                STATE_PASSTHROUGH: begin
                    if (!cached_mport_i[`BUS_MO_REQ]) begin
                        state <= STATE_READY;
                    end

                    cached_mport_o <= mport_i;
                    mport_o <= cached_mport_i;
                end
            endcase
        end
    end

endmodule