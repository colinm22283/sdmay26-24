// This is the unpowered netlist.
module busarb_2_2 (clk_i,
    nrst_i,
    mports_i,
    mports_o,
    sports_i,
    sports_o);
 input clk_i;
 input nrst_i;
 input [227:0] mports_i;
 output [135:0] mports_o;
 input [135:0] sports_i;
 output [227:0] sports_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire _3757_;
 wire _3758_;
 wire _3759_;
 wire _3760_;
 wire _3761_;
 wire _3762_;
 wire _3763_;
 wire _3764_;
 wire _3765_;
 wire _3766_;
 wire _3767_;
 wire _3768_;
 wire _3769_;
 wire _3770_;
 wire _3771_;
 wire _3772_;
 wire _3773_;
 wire _3774_;
 wire _3775_;
 wire _3776_;
 wire _3777_;
 wire _3778_;
 wire _3779_;
 wire _3780_;
 wire _3781_;
 wire _3782_;
 wire _3783_;
 wire _3784_;
 wire _3785_;
 wire _3786_;
 wire _3787_;
 wire _3788_;
 wire _3789_;
 wire _3790_;
 wire _3791_;
 wire _3792_;
 wire _3793_;
 wire _3794_;
 wire _3795_;
 wire _3796_;
 wire _3797_;
 wire _3798_;
 wire _3799_;
 wire _3800_;
 wire _3801_;
 wire _3802_;
 wire _3803_;
 wire _3804_;
 wire _3805_;
 wire _3806_;
 wire _3807_;
 wire _3808_;
 wire _3809_;
 wire _3810_;
 wire _3811_;
 wire _3812_;
 wire _3813_;
 wire _3814_;
 wire _3815_;
 wire _3816_;
 wire _3817_;
 wire _3818_;
 wire _3819_;
 wire _3820_;
 wire _3821_;
 wire _3822_;
 wire _3823_;
 wire _3824_;
 wire _3825_;
 wire _3826_;
 wire _3827_;
 wire _3828_;
 wire _3829_;
 wire _3830_;
 wire _3831_;
 wire _3832_;
 wire _3833_;
 wire _3834_;
 wire _3835_;
 wire _3836_;
 wire _3837_;
 wire _3838_;
 wire _3839_;
 wire _3840_;
 wire _3841_;
 wire _3842_;
 wire _3843_;
 wire _3844_;
 wire _3845_;
 wire _3846_;
 wire _3847_;
 wire _3848_;
 wire _3849_;
 wire _3850_;
 wire _3851_;
 wire _3852_;
 wire _3853_;
 wire _3854_;
 wire _3855_;
 wire _3856_;
 wire _3857_;
 wire _3858_;
 wire _3859_;
 wire _3860_;
 wire _3861_;
 wire _3862_;
 wire _3863_;
 wire _3864_;
 wire _3865_;
 wire _3866_;
 wire _3867_;
 wire _3868_;
 wire _3869_;
 wire _3870_;
 wire _3871_;
 wire _3872_;
 wire _3873_;
 wire _3874_;
 wire _3875_;
 wire _3876_;
 wire _3877_;
 wire _3878_;
 wire _3879_;
 wire _3880_;
 wire _3881_;
 wire _3882_;
 wire _3883_;
 wire _3884_;
 wire _3885_;
 wire _3886_;
 wire _3887_;
 wire _3888_;
 wire _3889_;
 wire _3890_;
 wire _3891_;
 wire _3892_;
 wire _3893_;
 wire _3894_;
 wire _3895_;
 wire _3896_;
 wire _3897_;
 wire _3898_;
 wire _3899_;
 wire _3900_;
 wire _3901_;
 wire _3902_;
 wire _3903_;
 wire _3904_;
 wire _3905_;
 wire _3906_;
 wire _3907_;
 wire _3908_;
 wire _3909_;
 wire _3910_;
 wire _3911_;
 wire _3912_;
 wire _3913_;
 wire _3914_;
 wire _3915_;
 wire _3916_;
 wire _3917_;
 wire _3918_;
 wire _3919_;
 wire _3920_;
 wire _3921_;
 wire _3922_;
 wire _3923_;
 wire _3924_;
 wire _3925_;
 wire _3926_;
 wire _3927_;
 wire _3928_;
 wire _3929_;
 wire _3930_;
 wire _3931_;
 wire _3932_;
 wire _3933_;
 wire _3934_;
 wire _3935_;
 wire _3936_;
 wire _3937_;
 wire _3938_;
 wire _3939_;
 wire _3940_;
 wire _3941_;
 wire _3942_;
 wire _3943_;
 wire _3944_;
 wire _3945_;
 wire _3946_;
 wire _3947_;
 wire _3948_;
 wire _3949_;
 wire _3950_;
 wire _3951_;
 wire _3952_;
 wire _3953_;
 wire _3954_;
 wire _3955_;
 wire _3956_;
 wire _3957_;
 wire _3958_;
 wire _3959_;
 wire _3960_;
 wire _3961_;
 wire _3962_;
 wire _3963_;
 wire _3964_;
 wire _3965_;
 wire _3966_;
 wire _3967_;
 wire _3968_;
 wire _3969_;
 wire _3970_;
 wire _3971_;
 wire _3972_;
 wire _3973_;
 wire _3974_;
 wire _3975_;
 wire _3976_;
 wire _3977_;
 wire _3978_;
 wire _3979_;
 wire _3980_;
 wire _3981_;
 wire _3982_;
 wire _3983_;
 wire _3984_;
 wire _3985_;
 wire _3986_;
 wire _3987_;
 wire _3988_;
 wire _3989_;
 wire _3990_;
 wire _3991_;
 wire _3992_;
 wire _3993_;
 wire _3994_;
 wire _3995_;
 wire _3996_;
 wire _3997_;
 wire _3998_;
 wire _3999_;
 wire _4000_;
 wire _4001_;
 wire _4002_;
 wire _4003_;
 wire _4004_;
 wire _4005_;
 wire _4006_;
 wire _4007_;
 wire _4008_;
 wire _4009_;
 wire _4010_;
 wire _4011_;
 wire _4012_;
 wire _4013_;
 wire _4014_;
 wire _4015_;
 wire _4016_;
 wire _4017_;
 wire _4018_;
 wire _4019_;
 wire _4020_;
 wire _4021_;
 wire _4022_;
 wire _4023_;
 wire _4024_;
 wire _4025_;
 wire _4026_;
 wire _4027_;
 wire _4028_;
 wire _4029_;
 wire _4030_;
 wire _4031_;
 wire _4032_;
 wire _4033_;
 wire _4034_;
 wire _4035_;
 wire _4036_;
 wire _4037_;
 wire _4038_;
 wire _4039_;
 wire _4040_;
 wire _4041_;
 wire _4042_;
 wire _4043_;
 wire _4044_;
 wire _4045_;
 wire _4046_;
 wire _4047_;
 wire _4048_;
 wire _4049_;
 wire _4050_;
 wire _4051_;
 wire _4052_;
 wire _4053_;
 wire _4054_;
 wire _4055_;
 wire _4056_;
 wire _4057_;
 wire _4058_;
 wire _4059_;
 wire _4060_;
 wire _4061_;
 wire _4062_;
 wire _4063_;
 wire _4064_;
 wire _4065_;
 wire _4066_;
 wire _4067_;
 wire _4068_;
 wire _4069_;
 wire _4070_;
 wire _4071_;
 wire _4072_;
 wire _4073_;
 wire _4074_;
 wire _4075_;
 wire _4076_;
 wire _4077_;
 wire _4078_;
 wire _4079_;
 wire _4080_;
 wire _4081_;
 wire _4082_;
 wire _4083_;
 wire _4084_;
 wire _4085_;
 wire _4086_;
 wire _4087_;
 wire _4088_;
 wire _4089_;
 wire _4090_;
 wire _4091_;
 wire _4092_;
 wire _4093_;
 wire _4094_;
 wire _4095_;
 wire _4096_;
 wire _4097_;
 wire _4098_;
 wire _4099_;
 wire _4100_;
 wire _4101_;
 wire _4102_;
 wire _4103_;
 wire _4104_;
 wire _4105_;
 wire _4106_;
 wire _4107_;
 wire _4108_;
 wire _4109_;
 wire _4110_;
 wire _4111_;
 wire _4112_;
 wire _4113_;
 wire _4114_;
 wire _4115_;
 wire _4116_;
 wire _4117_;
 wire _4118_;
 wire _4119_;
 wire _4120_;
 wire _4121_;
 wire _4122_;
 wire _4123_;
 wire _4124_;
 wire _4125_;
 wire _4126_;
 wire _4127_;
 wire _4128_;
 wire _4129_;
 wire _4130_;
 wire _4131_;
 wire _4132_;
 wire _4133_;
 wire _4134_;
 wire _4135_;
 wire _4136_;
 wire _4137_;
 wire _4138_;
 wire _4139_;
 wire _4140_;
 wire _4141_;
 wire _4142_;
 wire _4143_;
 wire _4144_;
 wire _4145_;
 wire _4146_;
 wire _4147_;
 wire _4148_;
 wire _4149_;
 wire _4150_;
 wire _4151_;
 wire _4152_;
 wire _4153_;
 wire _4154_;
 wire _4155_;
 wire _4156_;
 wire _4157_;
 wire _4158_;
 wire _4159_;
 wire _4160_;
 wire _4161_;
 wire _4162_;
 wire _4163_;
 wire _4164_;
 wire _4165_;
 wire _4166_;
 wire _4167_;
 wire _4168_;
 wire _4169_;
 wire _4170_;
 wire _4171_;
 wire _4172_;
 wire _4173_;
 wire _4174_;
 wire _4175_;
 wire _4176_;
 wire _4177_;
 wire _4178_;
 wire _4179_;
 wire _4180_;
 wire _4181_;
 wire _4182_;
 wire _4183_;
 wire _4184_;
 wire _4185_;
 wire _4186_;
 wire _4187_;
 wire _4188_;
 wire _4189_;
 wire _4190_;
 wire _4191_;
 wire _4192_;
 wire _4193_;
 wire _4194_;
 wire _4195_;
 wire _4196_;
 wire _4197_;
 wire _4198_;
 wire _4199_;
 wire _4200_;
 wire _4201_;
 wire _4202_;
 wire _4203_;
 wire _4204_;
 wire _4205_;
 wire _4206_;
 wire _4207_;
 wire _4208_;
 wire _4209_;
 wire _4210_;
 wire _4211_;
 wire _4212_;
 wire _4213_;
 wire _4214_;
 wire _4215_;
 wire _4216_;
 wire _4217_;
 wire _4218_;
 wire _4219_;
 wire _4220_;
 wire _4221_;
 wire _4222_;
 wire _4223_;
 wire _4224_;
 wire _4225_;
 wire _4226_;
 wire _4227_;
 wire _4228_;
 wire _4229_;
 wire _4230_;
 wire _4231_;
 wire _4232_;
 wire _4233_;
 wire _4234_;
 wire _4235_;
 wire _4236_;
 wire _4237_;
 wire _4238_;
 wire _4239_;
 wire _4240_;
 wire _4241_;
 wire _4242_;
 wire _4243_;
 wire _4244_;
 wire _4245_;
 wire _4246_;
 wire _4247_;
 wire _4248_;
 wire _4249_;
 wire _4250_;
 wire _4251_;
 wire _4252_;
 wire _4253_;
 wire _4254_;
 wire _4255_;
 wire _4256_;
 wire _4257_;
 wire _4258_;
 wire _4259_;
 wire _4260_;
 wire _4261_;
 wire _4262_;
 wire _4263_;
 wire _4264_;
 wire _4265_;
 wire _4266_;
 wire _4267_;
 wire _4268_;
 wire _4269_;
 wire _4270_;
 wire _4271_;
 wire _4272_;
 wire _4273_;
 wire _4274_;
 wire _4275_;
 wire _4276_;
 wire _4277_;
 wire _4278_;
 wire _4279_;
 wire _4280_;
 wire _4281_;
 wire _4282_;
 wire _4283_;
 wire _4284_;
 wire _4285_;
 wire _4286_;
 wire _4287_;
 wire _4288_;
 wire _4289_;
 wire \arbiter.crossbar[0] ;
 wire \arbiter.crossbar[1] ;
 wire \arbiter.crossbar[2] ;
 wire \arbiter.crossbar[3] ;
 wire \arbiter.master_handled[0] ;
 wire \arbiter.master_handled[1] ;
 wire \arbiter.master_handled[2] ;
 wire \arbiter.master_handled[3] ;
 wire \arbiter.master_sel[0][0] ;
 wire \arbiter.master_sel[0][1] ;
 wire \arbiter.master_sel[1][0] ;
 wire \arbiter.master_sel[1][1] ;
 wire \arbiter.master_sel[2][0] ;
 wire \arbiter.master_sel[2][1] ;
 wire \arbiter.master_sel[3][0] ;
 wire \arbiter.master_sel[3][1] ;
 wire \arbiter.slave_handled[0] ;
 wire \arbiter.slave_handled[1] ;
 wire \arbiter.slave_handled[2] ;
 wire \arbiter.slave_handled[3] ;
 wire \arbiter.slave_sel[0][0] ;
 wire \arbiter.slave_sel[0][1] ;
 wire \arbiter.slave_sel[1][0] ;
 wire \arbiter.slave_sel[1][1] ;
 wire \arbiter.slave_sel[2][0] ;
 wire \arbiter.slave_sel[2][1] ;
 wire \arbiter.slave_sel[3][0] ;
 wire \arbiter.slave_sel[3][1] ;
 wire \arbiter.state[0][0] ;
 wire \arbiter.state[0][1] ;
 wire \arbiter.state[1][0] ;
 wire \arbiter.state[1][1] ;
 wire \arbiter.state[2][0] ;
 wire \arbiter.state[2][1] ;
 wire \arbiter.state[3][0] ;
 wire \arbiter.state[3][1] ;
 wire clknet_0_clk_i;
 wire clknet_2_0__leaf_clk_i;
 wire clknet_2_1__leaf_clk_i;
 wire clknet_2_2__leaf_clk_i;
 wire clknet_2_3__leaf_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(_2573_));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(_2573_));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(_2932_));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(_0737_));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(_2807_));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(_2196_));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(_2569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(_2569_));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(_2569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4291__A (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__A (.DIODE(_4095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__4294__A (.DIODE(\arbiter.slave_handled[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__A (.DIODE(_4098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__4297__A (.DIODE(_4100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4303__A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__A1 (.DIODE(_4106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__A2 (.DIODE(_4107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4306__A (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__B (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4312__B (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__A (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__B (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__A (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4317__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__B (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__B (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__B (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A1 (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A2 (.DIODE(_4107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__B1 (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__B (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4327__B (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4329__B (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__4331__B (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4333__B (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4335__B (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__A (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4337__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4339__B1 (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4342__A (.DIODE(\arbiter.master_sel[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A (.DIODE(\arbiter.master_sel[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__A (.DIODE(_4147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4344__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__A (.DIODE(\arbiter.master_sel[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__B (.DIODE(\arbiter.master_sel[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__B (.DIODE(_4150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__A (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__B (.DIODE(\arbiter.master_sel[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4352__A (.DIODE(\arbiter.master_sel[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__B1 (.DIODE(_4156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__B (.DIODE(_4150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4366__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__B1 (.DIODE(_4145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A (.DIODE(_4106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__B (.DIODE(_4107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__B (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__4383__B (.DIODE(_4184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__A (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__B (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__A (.DIODE(_4145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__B (.DIODE(_4186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__B (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__C (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4392__B (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__B (.DIODE(_4095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__A (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__B (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__A (.DIODE(_4145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__B (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__B (.DIODE(\arbiter.slave_handled[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__B (.DIODE(_4098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__B (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__A (.DIODE(_4145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__B (.DIODE(_4213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__B (.DIODE(_4100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__A (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__B (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__A (.DIODE(_4223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A (.DIODE(_4145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__B (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__B (.DIODE(_4106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__C (.DIODE(_4107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__B (.DIODE(_4184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A (.DIODE(_4235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__B (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A (.DIODE(_4238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__A (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__B (.DIODE(_4245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A (.DIODE(_4243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__B (.DIODE(_4253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A0 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__B (.DIODE(\arbiter.slave_sel[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A (.DIODE(_4263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__B (.DIODE(_4245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__B1 (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__B2 (.DIODE(_4265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A1 (.DIODE(_4245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__B (.DIODE(_4107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__B1 (.DIODE(\arbiter.slave_sel[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__A (.DIODE(_4245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A (.DIODE(_4253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__B (.DIODE(_4245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A1 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__A2 (.DIODE(_4271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__B1 (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__4472__B2 (.DIODE(_4272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4473__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__A2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__B1 (.DIODE(_4245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4476__B (.DIODE(_4253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__A (.DIODE(_4272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__A (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4478__B (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__A (.DIODE(_4271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__A (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A (.DIODE(_4265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__B (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__B (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__B1 (.DIODE(_4253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__C (.DIODE(_4245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A (.DIODE(_4265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__A2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__B1 (.DIODE(_4150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4493__B2 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__B2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A (.DIODE(_4287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__B (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__A1 (.DIODE(_4286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A (.DIODE(_4235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__4502__B (.DIODE(\arbiter.crossbar[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__A (.DIODE(_4272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__B (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__A1 (.DIODE(_4286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__B (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__A (.DIODE(_4271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__B (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A1 (.DIODE(_4286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__B (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A (.DIODE(_0068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__A (.DIODE(_4263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__B (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__A1 (.DIODE(_4286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__B (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__A1 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__A2 (.DIODE(_4107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__B1 (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__A (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__B (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__A (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__B (.DIODE(_4107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__B (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__C (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4557__B (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__B (.DIODE(\arbiter.slave_sel[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A (.DIODE(_4107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__A (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4561__B (.DIODE(\arbiter.slave_sel[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4562__A (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__A (.DIODE(\arbiter.slave_sel[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__B (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4567__B (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__B2 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A2 (.DIODE(_0111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__B (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__C (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A1 (.DIODE(_0110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__B2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__A (.DIODE(_4150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__B (.DIODE(_0128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__A2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__B1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__B2 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__B (.DIODE(_0131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__B1 (.DIODE(_0079_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__B (.DIODE(_0134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4591__B (.DIODE(_4107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__B (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B (.DIODE(_0068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A2 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__B1 (.DIODE(_0068_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__B (.DIODE(_0134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__A (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__B (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A (.DIODE(_0111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__B (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__B (.DIODE(_0166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__A (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__B (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A (.DIODE(_4243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__A1_N (.DIODE(\arbiter.crossbar[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__B (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__B (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__A (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__B1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__B2 (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__A1 (.DIODE(_4150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__A2 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__B1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4646__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__A (.DIODE(\arbiter.slave_sel[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__B (.DIODE(\arbiter.slave_sel[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A (.DIODE(\arbiter.slave_sel[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__B (.DIODE(\arbiter.slave_sel[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__A (.DIODE(\arbiter.slave_sel[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A (.DIODE(\arbiter.slave_sel[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__A (.DIODE(\arbiter.slave_sel[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4654__A (.DIODE(\arbiter.slave_sel[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__A (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__B (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__A1 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__A2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__B2 (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__A1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__B2 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__B (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4658__C (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__A1 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A2 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__B2 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__B (.DIODE(_0191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__C (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__B (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4671__B (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4674__C (.DIODE(_4156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4685__B (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A (.DIODE(_4145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__B (.DIODE(_4150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__B (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4698__A (.DIODE(_4147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__B (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4700__A (.DIODE(_4145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4702__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__B (.DIODE(\arbiter.master_sel[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__B (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4709__C (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4710__B (.DIODE(_4145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4712__C (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__A (.DIODE(\arbiter.master_sel[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4717__B (.DIODE(\arbiter.master_sel[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4719__A (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4720__B (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__A (.DIODE(_4145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__B1 (.DIODE(_4243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4739__A (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4740__B (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4741__A1 (.DIODE(_4286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4742__B (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__B (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4746__B (.DIODE(_4150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4747__B (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4753__A (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4754__B (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__A1 (.DIODE(_4286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4756__B (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4760__A (.DIODE(_4243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4765__B (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__A1 (.DIODE(_4286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4767__B (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__A1 (.DIODE(_4286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4776__B (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4778__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A (.DIODE(_0131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__B (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__B (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__B (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A2 (.DIODE(_4150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__B1 (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4810__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4818__B (.DIODE(_4150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4821__B (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4822__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__B (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__B (.DIODE(_0166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__B (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__B1 (.DIODE(_4243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A2 (.DIODE(_4286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__B2 (.DIODE(_4235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__A1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__A2 (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__B1 (.DIODE(_0134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A1_N (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__4843__A2_N (.DIODE(_0026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A (.DIODE(_0020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4846__B1 (.DIODE(net737));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__A (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__B (.DIODE(_0020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__B (.DIODE(_0026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__A (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__A (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__A (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__A (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__A (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__B (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__A (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__A (.DIODE(_4184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__B (.DIODE(_4263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__B (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__A (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__A (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A (.DIODE(_4147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__A (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__A (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4896__A (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A1 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B2 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4898__B2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__A (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4901__A (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4903__B (.DIODE(_4223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A2 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__B2 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A (.DIODE(_0128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__A (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__A (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__A (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__A (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__A (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__A2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__B2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__A (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__B (.DIODE(_0134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A (.DIODE(_0460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__A (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__B (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__A (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__A (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__B (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4926__S (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4927__A (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4930__A (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__A (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__A (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4935__A (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__A (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__A (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__A (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__B1 (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__B2 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__B2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__A (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4944__B (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__A (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4947__B (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4948__A (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__A (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A1 (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__B2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4956__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__A1 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__A2 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__B1 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4958__B2 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__B2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__A1 (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__A2 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4961__B2 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__B2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__A1 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__S (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__B1 (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__4965__B2 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A1 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__B2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__A1 (.DIODE(_0505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__B2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4971__B (.DIODE(_4272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__B (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4975__A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__B (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A (.DIODE(\arbiter.master_sel[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4979__B1 (.DIODE(_4156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__B2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4980__C1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__B (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__A (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__B (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__A (.DIODE(_4235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4987__B (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__A2 (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4988__B1 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4989__A2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A1 (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__A2 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4991__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__A2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4992__B2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__S (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__B1 (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__B2 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A1 (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__B1 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__B2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A0 (.DIODE(_0531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4996__A1 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__4999__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__B2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5002__A (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A1 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__A2 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__B1 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5005__B2 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__A2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5006__B2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5007__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__B (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__A1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5010__B (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A (.DIODE(_4235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__B (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__B1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__A2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5016__B2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A (.DIODE(_4253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5019__B (.DIODE(_4272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5020__A (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5021__A (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5022__A (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5023__A1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5026__A1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__B1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__B2 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__B1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__B2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A1 (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__B2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5036__A (.DIODE(_0111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5038__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5041__A (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A (.DIODE(_0110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__B1 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__B2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__B1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5044__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A1 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5045__B2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A1 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__A2 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__B1 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5048__B2 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5049__B2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__S (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__A (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5054__A (.DIODE(_4223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__A1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5057__B1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5058__A3 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5061__A1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__A (.DIODE(_4184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__B (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__C (.DIODE(_4245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5062__D (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__A1 (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5063__C1 (.DIODE(_0598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__A (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5064__B (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__B (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__A1 (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5067__B1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A2 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A1 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A2 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__B1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__B2 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5073__B2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__A (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__A (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5075__B (.DIODE(_0608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A3 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5077__A (.DIODE(_4265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5079__A (.DIODE(_4287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5081__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A2 (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__5085__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__A (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5087__B (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A1 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__A2 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__B1 (.DIODE(_4271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5088__B2 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5089__A (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5091__A (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5093__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__B (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5095__A1 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5098__A (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A1 (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__A2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5099__B1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__A1 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__B2 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5101__A (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5104__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5105__A (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5106__A (.DIODE(_0110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A1 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__B1 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__B2 (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5108__A (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__B (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5111__A (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__B1 (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__5112__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A1 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A2 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__B1 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5114__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A2 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5117__A (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5120__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A (.DIODE(_0656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A1 (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A2 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__B1 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__B2 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__A (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A2 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__B2 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5127__A2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A (.DIODE(_4147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A2 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__A2 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__B1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__B2 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5133__A (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A1 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A2 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__B2 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__C1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__A2 (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A2 (.DIODE(_0656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A1 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A2 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__B1 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__B2 (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__B2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5143__A (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5145__A (.DIODE(_4223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__B (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A2 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__B2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__B (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5149__A (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__B (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A2 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__B1 (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A2 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__A2 (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5154__B1_N (.DIODE(_0686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__A2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5156__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__A (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__B (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A2 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__B1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__B2 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A (.DIODE(_4186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__A1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__B1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5163__B2 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A2 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A2 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__B2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__A2 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__B1 (.DIODE(_4147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__B2 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__B1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__B2 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A1 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__A2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5170__B1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__A (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5171__B (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__S (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__A2 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5175__B2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__B (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__B2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A1 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__B1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__B2 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5182__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__B2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__B1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__B2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__B (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__B (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__A (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5190__B (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5193__A (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__B1 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A1 (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A (.DIODE(_0111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__A (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A1 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__B1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__B2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A1 (.DIODE(_0460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__B2 (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__C1 (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A2 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5204__B2 (.DIODE(_0189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A2 (.DIODE(_0182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A1 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A2 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__B1 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__B2 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__B1 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A1 (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A1 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__S (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5211__A (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__B (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5213__C (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__A2 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__B2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5214__C1 (.DIODE(_0744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__B2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A2 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__B1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__B1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__B1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__B2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__B1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__B2 (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A1 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__B1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__B2 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__A (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5230__B (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5232__S (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A2 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__B1 (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__C1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A2 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__B2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5238__A (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__A (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__A (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A2 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__B2 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A1 (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__B1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__B2 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__B1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5246__B2 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__S (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__A (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__B (.DIODE(_0460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__B1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__5250__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__B1 (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__B2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A1 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__B1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__B2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A (.DIODE(_4272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__5258__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__A (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5260__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__S (.DIODE(_4253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__B (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5263__A1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__A1 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__B1 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5267__B2 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__A2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5268__B2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__A2 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5270__A (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5271__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__A (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__B2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A2 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__B1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__B2 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__B (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5282__B (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5283__A2 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__S (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__B2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A1 (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5287__B1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__B (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A1 (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__B1 (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__A2 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__B1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__A (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__B (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A2 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__B1 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5296__B2 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__B (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5300__A2 (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__A2 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5304__B2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5305__A (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__A2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__B1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5306__B2 (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A1 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__B1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__B2 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5308__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__A1 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__A2 (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__B2 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__A2 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5312__B1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5315__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__A (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5317__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__S (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__B (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A1 (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__B (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5323__A (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__B (.DIODE(_0460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__B1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__A2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5326__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__B (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__A1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A2 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__B2 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__A (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5333__B (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__B1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A1 (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__A2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__B1 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5339__B2 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5340__B2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__A (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5341__B (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__A2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__B2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5343__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5346__B (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A1_N (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5347__A2_N (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5348__B (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__5349__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5350__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__A2 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__B1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5351__B2 (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__B (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A1 (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__B (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__B (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A1 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__B (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5360__A (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5363__A (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__B1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A1 (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__A (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5370__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5371__S (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5372__B (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5373__A1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__B2 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__A2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__B2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__B1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5378__B2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__B1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A1 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5380__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A1 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__B1 (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__B2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__C1 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5382__A1 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5385__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5386__A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__B (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__B1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5393__A1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__B2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__C1 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A1 (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A2 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__B1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5397__B (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A2 (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5399__A2 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__A (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__B2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__B (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__S (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__A1 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5407__S (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__B (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__B (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5410__B1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A1 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A (.DIODE(_0936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__B (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A2 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A2 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__A2 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__B1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5416__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__A2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__B2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5418__B2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__A2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5419__B2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__B2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__A2 (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__B1 (.DIODE(_4265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5421__B2 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__A (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__B (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5422__C (.DIODE(\arbiter.slave_sel[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5423__A2 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__A (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__A (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__B (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5425__C (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__A2 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5427__B2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A1 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__A2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5428__B1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__A1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5429__B2 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5430__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A2 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__A2 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__B1 (.DIODE(_0953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A1 (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A2 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__A2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__B2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__B (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5443__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__B (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__S (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A0 (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__S (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A1 (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A2 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A1 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__A2 (.DIODE(_4265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__B1 (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__B2 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__B2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__A2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__B2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__A2 (.DIODE(_4265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__B1 (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5451__B2 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A1 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__A2 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5455__B2 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__A2 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5456__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__B2 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A1 (.DIODE(_0980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__S (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A0 (.DIODE(_0981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5463__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A2 (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__B2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A1 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__A2 (.DIODE(_4265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__B1 (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__B2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5474__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A1 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__B1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5476__B2 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__A2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5477__B2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__A2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5478__B2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__A2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5480__B2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__A2 (.DIODE(_4265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B1 (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5481__B2 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5482__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5483__A1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5484__S (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5486__S (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5487__B (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__A2 (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__B1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5488__C1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5489__B2 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__A (.DIODE(_1011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5490__B (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A1 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__A2 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5491__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__B1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__B2 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A2 (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A2 (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__A2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5496__B2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A2 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A2 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__B1 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__B2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__B2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__A1 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__B1 (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__B2 (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__S (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A2 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__B2 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__C1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A1 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__B1 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__B2 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__B (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A2 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__B1 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__A (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__B (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__S (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__A (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5517__A1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5518__A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5519__A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A1 (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__A2 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__B1 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5520__B2 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5521__B2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5522__A (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5525__B2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5526__B (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A2 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__C1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A2 (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__B1 (.DIODE(_1048_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__B2 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5530__B2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5531__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5532__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A1 (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__B1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5533__B2 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A1_N (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A2_N (.DIODE(_1055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__B1 (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__B2 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__A2 (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__B1 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A1 (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__A3 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5542__B1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__A2 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5543__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A1 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__A2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__B1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5544__B2 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__A2 (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__A2 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__5547__B2 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5548__B2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5549__A (.DIODE(_1029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__A3 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5550__B1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A1 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__B1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__B2 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__S (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A2 (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__B2 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__A2 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5556__B1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__A2 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__B1 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__5557__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A1 (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__B1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__B2 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__A2 (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__B1 (.DIODE(_0111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5559__B2 (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__B2 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__A2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A1 (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A2 (.DIODE(_0111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__B1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__B2 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__A2 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__B1 (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__C1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A2 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__B1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__B2 (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__S (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5575__A (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A2 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__B (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__S (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__A (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A2 (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__A3 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5582__B1 (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5583__A (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5584__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__A1 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5585__B2 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A0 (.DIODE(_1103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__A1 (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5586__S (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5587__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A1 (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__A2 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5588__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A1 (.DIODE(_1106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A1 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__A2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__B1 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5593__B2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A (.DIODE(_1111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A1 (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A2 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__B1 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__B2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5601__A (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A1 (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__A2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5604__B2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__A (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5605__B (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5606__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__A3 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__A (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5609__B (.DIODE(_1111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5610__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5612__A1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5613__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5614__A1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5615__A (.DIODE(_4186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__B (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__B2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A1 (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__B1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5619__B2 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__S (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A2 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__B2 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__A2 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__B1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A2 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__B2 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__A (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__B (.DIODE(_0111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A1 (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__B (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A1 (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__B (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__B (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A1 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__B1 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5636__A1 (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A1 (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A1 (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A1 (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__A (.DIODE(_1158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__S (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__A (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__A (.DIODE(_1106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5645__B (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5646__A1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A2 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A2 (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__B2 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A1 (.DIODE(_1139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5650__A2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A1 (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__A2 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__B1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__B2 (.DIODE(_1158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5653__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5654__A (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5655__B (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__S (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__A (.DIODE(_1121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__B (.DIODE(_4106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5660__B (.DIODE(_4235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A2 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__B2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5665__B (.DIODE(_1180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__B (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__C (.DIODE(_1116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5668__A1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5669__S (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5670__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5671__A1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5673__B1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5674__A (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5675__A1 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__A1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__B1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__A2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__B1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__B1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__B2 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A (.DIODE(_1158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__B1 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__B2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__B (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__S (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5685__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__A1 (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__A2 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__B1 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__B2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__B (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__A1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__S (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__B2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__C1 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A1 (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A2 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__B1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A1 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5697__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A1 (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5699__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__B2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A1 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__B1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5701__B2 (.DIODE(_1215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__B (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5703__A1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__A2 (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__B1 (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5705__C1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A1 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A2 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__B2 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__C1 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5709__A (.DIODE(_1180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5710__S (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__A (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5712__A1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5714__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__B (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__A2 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__B2 (.DIODE(_1229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5716__C1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A2 (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__B1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A1 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5718__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A1 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__B1 (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__B2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A1 (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__A2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__B1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5720__B2 (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A2 (.DIODE(_4106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__B1 (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5722__A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A1 (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__A2 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5724__B1 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__B2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__A (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5726__B (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5728__A1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__S (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__A (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5730__B (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5731__B2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__B2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5733__B2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A1 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__B1 (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__B2 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5735__A (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5737__B (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__B (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__C (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5739__B1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A2 (.DIODE(_1215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__B1 (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5741__A (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__B1 (.DIODE(_1252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__5743__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__B1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A2 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__B1 (.DIODE(_4147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__A2 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__B1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5747__B2 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5749__B (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A1 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A2 (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5751__A3 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5753__A1 (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A1 (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__B1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__B2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A1 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A2 (.DIODE(_4265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__B1 (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__B2 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5760__B (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A1 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__A2 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__B2 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A1 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A2 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__B1 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A1 (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__B1 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__B2 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__A1 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__S (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5767__A (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__A2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__B1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5772__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A1 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__A2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__B1 (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__B2 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A1 (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__B1 (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__B2 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__B (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5777__A1 (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__B (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A2 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__B1 (.DIODE(_1278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__B2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A (.DIODE(_4263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__B (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5783__A (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__A1 (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__B2 (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A1 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__B2 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A1 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__B1 (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__B2 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A1 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__B1 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__5788__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__B1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__B2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A1 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A1 (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__A2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__B1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__5793__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A1 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__A2 (.DIODE(_0111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__B1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__B2 (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__B (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5798__B (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__A (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__B (.DIODE(_0460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A2 (.DIODE(_1297_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A2 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__B1 (.DIODE(_1312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5803__A (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5804__A (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__A2 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__A2 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5811__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__B (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__S (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5815__S (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__B (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__B (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__B1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5819__A1 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A (.DIODE(_1329_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__B (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A2 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__A2 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5823__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__B2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A2 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__B1 (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__B2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__B (.DIODE(_4106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5828__B (.DIODE(_4235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__B (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__C (.DIODE(_1259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__A1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5832__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__B (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A1 (.DIODE(_0548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__B2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__A2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__B2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A2 (.DIODE(_0039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__B2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__B2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5838__B2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A1 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__B1 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__B2 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A2 (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__B1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__B2 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__B (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__B (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__B (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__B1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A2 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__B1 (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A1 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__B1 (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__B2 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A2 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__B1 (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A2 (.DIODE(_4265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__B1 (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__B2 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5856__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__B2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__B (.DIODE(_4272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A1 (.DIODE(_4287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__B1 (.DIODE(_4253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__B (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A2 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A2 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5875__B (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__S (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__S (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A1 (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__A (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__B (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__B2 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__A1 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__B1 (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__A0 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__A1 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__S (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__B1 (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__B2 (.DIODE(_1395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__B1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__B2 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5891__B (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A1 (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5893__B (.DIODE(_0487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A2 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__B2 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A1 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__A2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__B1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__B2 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A (.DIODE(_1395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__B (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__A1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__S (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A1 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__B1 (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__B (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__B (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__A (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__B (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__B2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5913__S (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__B (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A1 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A1 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__B2 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A (.DIODE(_1424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__B (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A2 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__B1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__A (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__S (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A1 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__B1 (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5931__A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A1 (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A2 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__B1 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__B2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__B (.DIODE(_1440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A1 (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A2 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__B1 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__B2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__A (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__B (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__C (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__S (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A2 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__B2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A (.DIODE(_1452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__B (.DIODE(_4272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__A1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__B (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A1 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A1 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__A2 (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__B2 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A2 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__B1 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__A2 (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__B1 (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__C1 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A2 (.DIODE(_1395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__B1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__A (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__S (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A2 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A1 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A1 (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__B1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__B2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__A (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__A (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A1 (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A2 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__B1 (.DIODE(_0434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__B2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__B (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A2 (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A3 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A1 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A2 (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__B1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__A1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A1 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__S (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__A (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__B (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A1 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__A1 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__A2 (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__B2 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__A2 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__B1 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A2 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__B1 (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__C1 (.DIODE(_1490_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A2 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__B1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5988__A (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A2 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__A (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__B (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__C (.DIODE(_1473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__S (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__B (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5998__A (.DIODE(_1440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__B (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6000__B1 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__B (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__A (.DIODE(_1452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__A2 (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__B1_N (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6004__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__A2 (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__A (.DIODE(_1509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6006__B (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A1 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__A1 (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__B1 (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__A2 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__A1 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__A2 (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__B2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__B (.DIODE(_4272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__A1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__S (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A1 (.DIODE(_0263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A2 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__A2 (.DIODE(_0424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__B2 (.DIODE(_0429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__A (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__B (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__S (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__S (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__A1 (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__A1 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__B2 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A1 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A1 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A0 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__A1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__S (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__A1 (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__A2 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__S (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__A (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__B (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__A2 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A2 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A3 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__S (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A1 (.DIODE(_0677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__B2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__A1 (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__A2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__B1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__B2 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__A (.DIODE(_1539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__A (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__B (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__A1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A1 (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__A1 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__B1 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__A (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6063__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__B (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__A1 (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__A2 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__A2 (.DIODE(_1539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__B1 (.DIODE(_1559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__B2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__B (.DIODE(_4272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__S (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__A (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A2 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__B1 (.DIODE(_0804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__B2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__A2 (.DIODE(_0425_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__B2 (.DIODE(_0430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__B (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6081__S (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__S (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A1 (.DIODE(_0441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__B2 (.DIODE(_0443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__B (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__A1 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__B2 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A2 (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__B2 (.DIODE(_0725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A2 (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A1 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__S (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A1 (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__A0 (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__A1 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__A2 (.DIODE(_0186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__B2 (.DIODE(_0477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A2 (.DIODE(_0467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__B2 (.DIODE(_0185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__A (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__B (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A1 (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A2 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__A2 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__B2 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__A2 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__A2 (.DIODE(_0128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__B2 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__A (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__B (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6103__S (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A1 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A1 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__A (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__A (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6107__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__A (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__A1 (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__B (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__A1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__B (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__A (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__A1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__B (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A1 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__A2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A2 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__B1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__B2 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__B (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A2 (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__S (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__A (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__B (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__A2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6126__B1 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A1 (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A2 (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__B1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__B (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A1 (.DIODE(_0463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__B1 (.DIODE(_0601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A2 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__B1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6131__A1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__A1 (.DIODE(_0550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__B2 (.DIODE(_0706_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__B (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__A1 (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__B1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__B1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__B2 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A1 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__B1 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A1 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__B1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6139__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A1 (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__B1 (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__6140__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6141__A1 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__A1 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__A2 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__B1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__B2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A2 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__B1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__B2 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__S (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A1 (.DIODE(_0645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__A2 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6145__B2 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__A1 (.DIODE(_1634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__A2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__6147__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__A2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6148__B2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__A (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6149__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A2 (.DIODE(_0411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__B1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__B2 (.DIODE(_0413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A2 (.DIODE(_0409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__B2 (.DIODE(_0492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6152__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__S (.DIODE(_4253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__B (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A1 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__A2 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__B1 (.DIODE(_0435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6159__B2 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__A2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__B2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6161__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__A2 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6162__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A2 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__B1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__B2 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__A1 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6164__B1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__A1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__B (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A1 (.DIODE(_0703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__A2 (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6168__C1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__A1 (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__A2 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6169__B1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6170__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__A2 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__6171__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__A2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__B2 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6173__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A1 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A2 (.DIODE(_0123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__B1 (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__B2 (.DIODE(_0122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__A2 (.DIODE(_0365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__B1 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__6175__B2 (.DIODE(_0449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__S (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__S (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__B (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6180__A (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6181__B (.DIODE(_0460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__A1 (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__A2 (.DIODE(_0474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__B1 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__6182__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__A1 (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__A (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6185__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__S (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__A2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__B1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6187__B2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6188__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6189__A1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__B2 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__A2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__S (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A2 (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6195__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__A (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6196__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__S (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__S (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__B (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__C (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__A1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6200__B1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6201__B1 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6202__B (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__A (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__B (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6206__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__A (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__S (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6209__B (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6210__A1 (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6211__B (.DIODE(_0462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__A (.DIODE(_0461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6212__B (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A1 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__B1 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6213__B2 (.DIODE(_0478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__A2 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6214__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__S (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6218__A1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A2 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__B2 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__A2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__A1 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__A2 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__B1 (.DIODE(_1717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6222__B2 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__A1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6223__S (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A0 (.DIODE(_1719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6224__A1 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6226__A (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A1 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A2 (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__B1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__B2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__B2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__A (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__B (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__C (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__D (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A1 (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A2 (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6233__B (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__A (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6234__B (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__A2 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6235__B1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6236__A2 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6237__A1 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__A2 (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6238__B2 (.DIODE(_0456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__A2 (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__B2 (.DIODE(_0452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A2 (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6242__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A2 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__B1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__B2 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A1 (.DIODE(_1735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A2 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__B1 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__B2 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__C1 (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A1 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A2 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__A1 (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__B1 (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__B2 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__B1 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__B2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__A1 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6249__S (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__6251__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__A2 (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6254__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A1 (.DIODE(_0432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A2 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__B1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__B2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__B2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6258__A2 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6258__B2 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6258__C1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__A2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6260__B2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__A (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6261__B (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__A1 (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__B1 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__6262__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A2 (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__B1 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__A (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__A1 (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__A2 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6265__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6266__B (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__B (.DIODE(_1759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__B2 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__B2 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__A2 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__B1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6272__B2 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__6273__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6274__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A2 (.DIODE(_0036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__B2 (.DIODE(_4289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A2 (.DIODE(_0407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__B2 (.DIODE(_0038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A (.DIODE(_1768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__A (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__B2 (.DIODE(_0626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6280__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6280__A2 (.DIODE(_0408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6280__B2 (.DIODE(_0624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6281__A1 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6281__S (.DIODE(_0557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__A1 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__A2 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6282__B2 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6283__A (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__A1 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__B2 (.DIODE(_0631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__A1 (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__B1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__A2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__B1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__B2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__S (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__A1 (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__A2 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__B (.DIODE(_1759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6291__A2 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A2 (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6294__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__A2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__B2 (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__6296__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A2 (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__A1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__A2 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__B2 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__C1 (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A1 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A2 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__B1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__B2 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__A2 (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6302__B2 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__A (.DIODE(_0591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__B (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6305__A3 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__A2 (.DIODE(_1768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__B2 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__A2 (.DIODE(_0604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__B1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__A1 (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__A2 (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6308__B1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__B1 (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A1 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__B2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__A1_N (.DIODE(_1759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__B1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6311__B2 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6312__A (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__A1 (.DIODE(_0660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__A (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__A (.DIODE(\arbiter.master_sel[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__B (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__B1 (.DIODE(_4156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__A2 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__B2 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6318__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__A2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__B2 (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__B (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6322__A (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A1 (.DIODE(_4271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A2 (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__C1 (.DIODE(_0419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__A1 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__A2 (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__B1 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__B2 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__A1 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__B1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__6325__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A1 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__B2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A1 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__S (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A1 (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__A2 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6328__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__B (.DIODE(_1759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__A2 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6331__B2 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__A2 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__B1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__6332__B2 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__A2 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__B1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__A2 (.DIODE(_0417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__B1 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A1 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__A2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__B2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__S (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__A1 (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6339__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__B (.DIODE(_1759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__A (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__B (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__C (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__D (.DIODE(\arbiter.slave_sel[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A1 (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A2 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__B1 (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__B2 (.DIODE(_0632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__C1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A1 (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__A2 (.DIODE(_0191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__B (.DIODE(_1759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A1 (.DIODE(_0131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A2 (.DIODE(_0682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__B1 (.DIODE(_1830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A1 (.DIODE(_0191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A2 (.DIODE(_0567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__A2 (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__B2 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__A2 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__B1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__B2 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__A1 (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__A2 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6353__B2 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__A2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__B2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__S (.DIODE(_0465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A1 (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__B1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__B2 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__B1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__B2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__A1 (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__S (.DIODE(_0489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__A2 (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__B2 (.DIODE(_0479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A2 (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__B2 (.DIODE(_0472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6363__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__B2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__B2 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A2 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__B1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__B2 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A1 (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__B1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6368__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A2 (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__B1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A1 (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__A2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6370__B1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A1 (.DIODE(_0418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__B1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A1 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__B1 (.DIODE(_0420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__A1 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A1 (.DIODE(_4105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__B (.DIODE(_1759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6377__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6378__A2 (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6378__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__6378__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A1 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A2 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__B1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__B2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A2 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__B2 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__A1 (.DIODE(_0592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__A2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__6384__B2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__S (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A1 (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__B1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__B2 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__B1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__B2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__A (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__A2 (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6391__B2 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A2 (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__B2 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A2 (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__B2 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__A2 (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__B2 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__B (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__B2 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A2 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__B1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__B2 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__A2 (.DIODE(_0422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__B2 (.DIODE(_0447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6398__C1 (.DIODE(_0633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__A1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A1 (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__B1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__B2 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__B1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__B2 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__A (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__B (.DIODE(_1885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__A2 (.DIODE(_0636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__A (.DIODE(_4100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6404__B (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__A (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__A (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__B (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__B (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__A (.DIODE(_4100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__A (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6411__A (.DIODE(_4213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__A (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__B (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__B (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__A2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__B2 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__A (.DIODE(_4100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__B (.DIODE(_0134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6418__A (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__A (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__B (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__B (.DIODE(_1902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__S (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__A (.DIODE(_4100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__B (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6424__A (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__A (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__B (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__B (.DIODE(_1908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__A1 (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__S (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__A (.DIODE(_1912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__B (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__B1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A (.DIODE(_4235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__B (.DIODE(_4100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6436__A (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__A1 (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__A2 (.DIODE(_0498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__B (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__A (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__B (.DIODE(_4272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__A (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6443__B (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__B1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6449__A (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__A1 (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__A2 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__B1 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__A1 (.DIODE(_0505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6452__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__A1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A3 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__B1 (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__A2 (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__B (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__B (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__A (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__B2 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__A (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A2 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__B2 (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6464__S (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A1 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__S (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__A (.DIODE(_1946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__A2 (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__B2 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__C1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__A (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__B (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A1 (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A2 (.DIODE(_0438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__B1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__B1 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A3 (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__B2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6477__B (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__C1 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A1 (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A2 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__B2 (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6481__B (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__A1 (.DIODE(_0718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__A2 (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__A1_N (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6483__B2 (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A1 (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6485__S (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__A1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__S (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A (.DIODE(_1965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6489__A (.DIODE(_0621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6490__S (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6491__B (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A1 (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A2 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__B1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6494__A (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__A (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6495__C (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__B (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6498__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__A (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__A1 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__A2 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__B1 (.DIODE(_0597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__B2 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__C1 (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__A1 (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6502__A2 (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__A (.DIODE(_1902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6505__A (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__A (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__B (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A1 (.DIODE(_1980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__B1 (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__A (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__A (.DIODE(_1908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__B (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__A2 (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__A3 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__B (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__A1_N (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__B2 (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__A2 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__B1 (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A2 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__A1 (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__C1 (.DIODE(_1996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__A (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__A1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__B2 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6525__B (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__A (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A1_N (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__B2 (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__A (.DIODE(_1902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__A2 (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__B2 (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__C1 (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__A2 (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A1 (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A2 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__B1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__B2 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__A1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__A (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__A1 (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__A1 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__A2 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__B1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__B2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__S (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__A1 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__B2 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__B (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__A (.DIODE(_1976_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__B (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__S (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A1 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A2 (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__B1 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__B2 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__A (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__B1 (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__A (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__A (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__B (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__A (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__A1 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__A2 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__B1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__B2 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A2 (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__C1 (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__B2 (.DIODE(_1908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__B (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__B (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__A (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__B (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__B (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__A1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__A (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__B (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__A (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__S (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__A (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__A2 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A2 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__A (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__A (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__B (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__C (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__B (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__A (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6578__B (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A2 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A (.DIODE(_2051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__B (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6581__B (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__A1 (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6584__B (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__B (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__A1 (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A2 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6589__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__A3 (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__B1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6592__B2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A (.DIODE(_0781_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6594__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__A1_N (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__B1 (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__B2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__A2 (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__B1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__A (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__B (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A1 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A2 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__B2 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__A1 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__B2 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A2 (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__B1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A2 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__B1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__B2 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__B2 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A2 (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__B1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__A2 (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__B1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__B (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A1 (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__B (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__B (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A (.DIODE(_2087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__B (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__B (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__A1 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__A2 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__B (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__S (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__B (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__B (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A1 (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__B2 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__B (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6633__B (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__A (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6634__B (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__A (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__B1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__B2 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A2 (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__C1 (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__A2 (.DIODE(_1908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6640__C1 (.DIODE(_2106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A1 (.DIODE(_0980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A2 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__B1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__B2 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__S (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__B (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6646__B (.DIODE(_0929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__A (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__B (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6649__A2 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__A2 (.DIODE(_0980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__B1 (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__A2 (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__B2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__A (.DIODE(_0966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6654__A2 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__B2 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__B2 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A2 (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__B1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A (.DIODE(_0980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6660__S (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6661__S (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6662__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A1 (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A2 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__B1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A1 (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__B1 (.DIODE(_2122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A1 (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A2 (.DIODE(_0111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__B1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__B2 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6667__S (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__B (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__B (.DIODE(_0961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__A (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6671__B (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6672__A2 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__A2 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6673__B1 (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__A2 (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__B1 (.DIODE(_2136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6674__B2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A1 (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__A (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__B (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__C (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__D_N (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__B (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__A (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6679__B (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A2 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__B (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__B1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__B2 (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6683__A (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__A2 (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6684__B1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__B1 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6685__B2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__A1_N (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6686__B2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A1 (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6687__B2 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__A2 (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6688__B1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__S (.DIODE(_0761_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A2 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__B1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A0 (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__S (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__B (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__B (.DIODE(_1096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__A (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6697__B (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A1 (.DIODE(_1055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A2 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__B (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__A2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__B1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6700__B2 (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__A2 (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6702__B1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__B1 (.DIODE(_1106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__B2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__A2 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__B1 (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6705__S (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__A2 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__B2 (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A2 (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__B2 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__A2 (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6708__B1 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A2 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__C1 (.DIODE(_2168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A1 (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6711__S (.DIODE(_0813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A2 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__B2 (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__B (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A1 (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__A2 (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__B2 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6714__C1 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A1 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A1 (.DIODE(_1158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__C1 (.DIODE(_2174_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__A1_N (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6717__B2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A1 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A2 (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__B2 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A2 (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__B1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6720__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__B (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A1 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A2 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A1 (.DIODE(_2177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__A (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__B (.DIODE(_1180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__A (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__B (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__A2 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__A (.DIODE(_2185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__B (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A1 (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__A2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__B1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__B2 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__A (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__A (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__B (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A1 (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__A2 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__A2 (.DIODE(_1215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__B1 (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__A (.DIODE(_1203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__A2 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__B2 (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__A2 (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__B2 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__A2 (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__B1 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__A2 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A1 (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__A (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__B (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__A1 (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__A1 (.DIODE(_1215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__A2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__B1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__B2 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__A2 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__B1 (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__A (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__B (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__A2 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__B2 (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__B (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__A2 (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6752__B1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__A2 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__C1 (.DIODE(_2207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A1 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__B (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__B (.DIODE(_1238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__A (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__B (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__A2 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__A (.DIODE(_2213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__B (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__B (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A1 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__A2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__B1 (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__B2 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__B (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__A1 (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A1 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__A2 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6769__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__A (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__B (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__A1 (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__A2 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__B1 (.DIODE(_1930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A1 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__A2 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__B2 (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__A1_N (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__B1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__B2 (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__A2 (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6776__B1 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__A2 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__A1 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__A1 (.DIODE(_0719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__A (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__A2 (.DIODE(_0704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__C1 (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__B (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__A2 (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__B1 (.DIODE(_2231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__B2 (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__A (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__B (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__S (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__A1_N (.DIODE(_1908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__B1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__B2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__A1 (.DIODE(_2238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__B2 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__A1_N (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__B1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__B2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__A2 (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__B1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A1 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__B1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__B2 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__B (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__A1 (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__A (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__B (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__B (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__A1 (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__A1 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__A2 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A1 (.DIODE(_2246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__A (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__B1 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__B (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__A (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__A2 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__A (.DIODE(_2262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__B (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A1 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__A2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__B1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__B2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__A (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__A (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__B (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__B (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__A1 (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__A2 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__A1 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__B1 (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A1 (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__B2 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__A1 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__A2 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__B2 (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__A2 (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__B1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__A (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__A (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__S (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__S (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__A1 (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__A2 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__B1 (.DIODE(_2273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__A1 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__B1 (.DIODE(_2281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__A1 (.DIODE(_4100_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__A2 (.DIODE(_0166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__B1 (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__B (.DIODE(_2283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__A1 (.DIODE(_1395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__A (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__B (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__A2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__B1 (.DIODE(_1895_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__B (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__A (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__B (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6842__A2 (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__A (.DIODE(_2290_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__B (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__A1 (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__B1 (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__B2 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6846__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__A (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__B (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__A1 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__A2 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__B (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__A (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__B (.DIODE(_1440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6854__A (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__A (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__B (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__A2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__B1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__B2 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__A (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__B (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__A1 (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__A2 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__B2 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__A1 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__A2 (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__B2 (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__A2 (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__B1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__A (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__A (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__B (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__S (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__S (.DIODE(_0841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__B (.DIODE(_2004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__A1 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__A2 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__B1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__A1 (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__B2 (.DIODE(_1988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__A1 (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__B (.DIODE(_0833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__C (.DIODE(_1923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__A2 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__A1 (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__A2 (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__A1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__B1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__B2 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__A1 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__B1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__B2 (.DIODE(_2324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__A1 (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__A2 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__A1 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__B1 (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__B (.DIODE(_2283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__A1 (.DIODE(_1539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__B2 (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__B (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__B (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__A (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__B (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__A (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__A1 (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__A1 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__A2 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__B1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__A1 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__B1_N (.DIODE(_2339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__A (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__B2 (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__B (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__B (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__A (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__B (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__A2 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__B1 (.DIODE(_1902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__B1_N (.DIODE(_2346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__A1 (.DIODE(_1539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__A2 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__B1 (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__B2 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__A (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__A1 (.DIODE(_0887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__A (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__B (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__B2 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__B (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__B (.DIODE(_1924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__B (.DIODE(_2023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__A (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__A1 (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__A1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__A2 (.DIODE(_1983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__B1 (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__C1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__A2 (.DIODE(_1908_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__C1 (.DIODE(_2359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__B (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__A1 (.DIODE(_1914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__B1 (.DIODE(_1917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__A2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__A3 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__A1 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__A2 (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__B2 (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__A (.DIODE(_1981_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__B (.DIODE(_1900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6926__A (.DIODE(_0886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__A1 (.DIODE(_1280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__A1 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__A2 (.DIODE(_1906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__A1 (.DIODE(_2364_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__A2 (.DIODE(_1932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__A2 (.DIODE(_1955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__B2 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__A (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__A2 (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__B1 (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__A1 (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__A2 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__B1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__A1 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__A (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__B (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__A1 (.DIODE(_1717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__A2 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__B2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__A1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__A (.DIODE(_2283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__A (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__B (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__A1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__B1 (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__A1 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__A (.DIODE(_1725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__A1 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__A2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__B2 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__A1 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__A (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__B (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__A1 (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__A2 (.DIODE(_1986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__A1 (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__A1 (.DIODE(_1735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__A2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__B1 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__B2 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__A1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__S (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__A1 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__S (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__A1 (.DIODE(_1973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__B1 (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__A1 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__A3 (.DIODE(_1997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__A2 (.DIODE(_1999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6958__B (.DIODE(_1929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__A1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__A2 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__B1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__A1 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__A1 (.DIODE(_1766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__A2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__B2 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__S (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__A1 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__S (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__A (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__B (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__A2 (.DIODE(_1892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__B2 (.DIODE(_1953_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__C1 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__A1 (.DIODE(_1768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__A2 (.DIODE(_1920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__B2 (.DIODE(_1889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__A (.DIODE(_1926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__A1 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__A2 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__B1 (.DIODE(_1931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__A1 (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__A2 (.DIODE(_1911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__A (.DIODE(_1772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__B (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__A1 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__A2 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__B2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__C1 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__A1 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__A1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__S (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__A2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__B2 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__S (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6978__S (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__A (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__A1 (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__A2 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__B1 (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__B2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__C1 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6982__A1 (.DIODE(_0131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6982__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__A0 (.DIODE(_2413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__A1 (.DIODE(_0191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__S (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__A1 (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__A2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__B2 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__C1 (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__A2 (.DIODE(_1947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__A1 (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__S (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__B (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6990__A2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__S (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__S (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__B (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__A2 (.DIODE(_1941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__S (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6997__S (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__A2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__B2 (.DIODE(_1898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__S (.DIODE(_1904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__A1 (.DIODE(_1885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__S (.DIODE(_1910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__A1 (.DIODE(_4235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__A2 (.DIODE(_4098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__B1 (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__B2 (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__A (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__A (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__A1 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__A2 (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__B2 (.DIODE(_4098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__B (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__A1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__B2 (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__A1 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__A2 (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__B2 (.DIODE(_4098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__A (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7012__S (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__A (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__A2 (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__B1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__B2 (.DIODE(_4098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7016__A (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__A1 (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7018__A (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7019__A (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7020__A (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__A1 (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__B2 (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__C1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7022__A (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__A1 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__A2 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__B1_N (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__A1 (.DIODE(_0505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__A1 (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__A (.DIODE(_2454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__A1 (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__A (.DIODE(_2458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__A (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__A2 (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__B2 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__C1 (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__A2 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7041__A1 (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7041__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__A (.DIODE(_2463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__A (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__A2 (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__B2 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__C1 (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__A1 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__A2 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__A1 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__A2 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__B1 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__A_N (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__A1 (.DIODE(_0576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__A0 (.DIODE(_2471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__A1 (.DIODE(_0656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7054__A2 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7054__B1 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__A1 (.DIODE(_0639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__A0 (.DIODE(_2475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__A1 (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__A (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__A (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7061__A (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__A1 (.DIODE(_0715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__B1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__B2 (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__C1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__A1 (.DIODE(_0727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__A0 (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__A1 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__A1 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__B1 (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__B2 (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__C1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__A1 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__A1 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__A1 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__A1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__A0 (.DIODE(_2488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__A1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__A1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__B2 (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__C1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__A1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__A1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__A1 (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__B1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__B2 (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__C1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__A1 (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__A1 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__A1 (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7084__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7085__A1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7085__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__A0 (.DIODE(_2498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__A1 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__A (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__A (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__A1 (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7090__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__A1 (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__A1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7094__A (.DIODE(_0867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__A1 (.DIODE(_0906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__A1 (.DIODE(_0877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7096__B1 (.DIODE(_2506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__A1 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__S (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__A (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__A1 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__A1 (.DIODE(_0955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7102__A (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__A0 (.DIODE(_2511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__A1 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__A (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__A1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__A1 (.DIODE(_0980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__A0 (.DIODE(_2516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__A1 (.DIODE(_0942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__A1 (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__A0 (.DIODE(_2520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__A1 (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__B (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__A1 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7118__A1 (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7118__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__A (.DIODE(_2525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7120__A (.DIODE(_1034_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7121__B (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__A1 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__A1 (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__A1 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__A (.DIODE(_2530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__A1 (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__B1 (.DIODE(_2531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7128__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7128__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__A (.DIODE(_2533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__A1 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__A1 (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__B1 (.DIODE(_2534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__A1 (.DIODE(_1106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7132__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__A1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__A1 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__B1 (.DIODE(_2537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7136__A1 (.DIODE(_1153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7136__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7137__A (.DIODE(_2539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7138__A (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7139__B (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__A1 (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7140__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__A1 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__A0 (.DIODE(_2543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__A1 (.DIODE(_1158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__A1 (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__A1 (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7146__A0 (.DIODE(_2546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7146__A1 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7146__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7148__B (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7149__A1 (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7149__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7149__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__A1 (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__A0 (.DIODE(_2550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__A1 (.DIODE(_1169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7153__B (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__A1 (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7155__A1 (.DIODE(_1215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7155__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__A0 (.DIODE(_2554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__A1 (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__A1 (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__A1 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__B1 (.DIODE(_2556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__A1 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__A1 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__A1 (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__B1 (.DIODE(_2559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__A1 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__A (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7166__A1 (.DIODE(_1269_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7166__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7166__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__A (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7168__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7168__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__A0 (.DIODE(_2564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__A1 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7170__A (.DIODE(_2565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7171__A (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__B (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7173__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7173__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7173__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7174__A1 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7174__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__A0 (.DIODE(_2569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__A1 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__S (.DIODE(_2512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__B (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__A1 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7179__A1 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7179__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__A (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__A0 (.DIODE(_2573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__A1 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__A (.DIODE(_2575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7183__B (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__A1 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__B1 (.DIODE(_2437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7185__A1 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7185__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7186__A0 (.DIODE(_2578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7186__A1 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7186__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7187__A (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7188__A1 (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7188__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7188__B1 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7188__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7188__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7189__A1 (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7189__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7190__A0 (.DIODE(_2581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7190__A1 (.DIODE(_1395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7190__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7191__A (.DIODE(_2582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7192__B (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__A1 (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__A2 (.DIODE(_2444_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7194__A1 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7194__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__A0 (.DIODE(_2585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__A1 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7196__A (.DIODE(_2586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__A1 (.DIODE(_1452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7198__A1 (.DIODE(_1512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7198__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7198__B1 (.DIODE(_2587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7199__A1 (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7199__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7200__A (.DIODE(_2589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7201__A1 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7201__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7201__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7201__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7202__A1 (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7202__A2 (.DIODE(_2448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7202__B1 (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7203__A1 (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7203__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7204__A (.DIODE(_2592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__A1 (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7205__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__A1 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__A0 (.DIODE(_2594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__A1 (.DIODE(_1539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7208__A (.DIODE(_2595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7209__B (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__A1 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7211__A1 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7211__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7212__A0 (.DIODE(_2598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7212__A1 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7212__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7213__A (.DIODE(_2599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__A1 (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7215__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7215__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__A0 (.DIODE(_2601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__A1 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7217__A (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7218__B (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__A1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__A0 (.DIODE(_2605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__A1 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__A (.DIODE(_2606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__A1 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__A_N (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7224__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__A1 (.DIODE(_1598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__A0 (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__A1 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7227__A (.DIODE(_2610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7228__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7229__A1 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7229__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7230__A0 (.DIODE(_2612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7230__A1 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7230__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7231__A (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7232__A1 (.DIODE(_1717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7232__A2 (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7232__B2 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7232__C1 (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7233__A1 (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7233__A2 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7235__A1 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7235__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7236__A (.DIODE(_2617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__A1 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__A1 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7239__A1 (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7239__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7240__A (.DIODE(_2620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7241__A1 (.DIODE(_1735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7241__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7241__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7242__A (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7242__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7243__A1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7243__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7244__A1 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7244__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7245__A (.DIODE(_2624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7246__B (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7247__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7247__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7248__A1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7248__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7249__A1 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7249__S (.DIODE(_2574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7250__A (.DIODE(_2628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7251__A (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__A2 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__B2 (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7252__C1 (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7253__A2 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__A1 (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7255__S (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7256__A (.DIODE(_2633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__A1 (.DIODE(_1768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__B2 (.DIODE(_2500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7257__C1 (.DIODE(_2501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7258__A1 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7258__A2 (.DIODE(_2450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7259__A1 (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7259__S (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7260__A (.DIODE(_2636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7261__A1 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7261__A2 (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7261__B2 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7261__C1 (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7262__A1 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7262__A2 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7264__A1 (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7264__S (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7265__A (.DIODE(_2640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7266__B (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__A2 (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__B2 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7267__C1 (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7268__A2 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7270__S (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7271__A (.DIODE(_2645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__B (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7272__C (.DIODE(_2432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7273__A1 (.DIODE(_0041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7273__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7273__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7274__A1 (.DIODE(_0131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7274__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7275__A0 (.DIODE(_2648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7275__A1 (.DIODE(_0191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7275__S (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__A1 (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7277__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7278__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7279__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__A1 (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7280__S (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7281__A (.DIODE(_2653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7282__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7282__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7283__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7284__A2 (.DIODE(_2540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7285__S (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7286__A (.DIODE(_2657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7287__A2 (.DIODE(_2477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7287__B1 (.DIODE(_2479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7288__B (.DIODE(_2445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7289__A2 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7290__S (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7291__A (.DIODE(_2661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7292__A2 (.DIODE(_2429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7292__B2 (.DIODE(_2434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7292__C1 (.DIODE(_2436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7293__A2 (.DIODE(_2447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7295__A1 (.DIODE(_1885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7295__S (.DIODE(_2441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7296__A (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7297__A (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7297__B (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7298__A (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7299__A (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7299__B (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7300__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7300__B (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7301__A (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7302__A (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7303__A (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7304__A (.DIODE(_4186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7304__B (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7305__A (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7305__B (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7306__A (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7307__A (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7308__A1 (.DIODE(_0416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7308__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7308__B2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7309__A (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7309__B (.DIODE(_0134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7310__A (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7311__A (.DIODE(_0111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7311__B (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7312__A (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7312__B (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7314__S (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7315__A (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7315__B (.DIODE(_4095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7316__A (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7317__B (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7318__A1 (.DIODE(_0482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7318__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7320__A1 (.DIODE(_0494_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7320__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7320__B2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7321__A1 (.DIODE(_0502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7321__S (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7322__A1 (.DIODE(_0505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7322__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7325__A (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7326__A (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7327__A2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7327__B2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7327__C1 (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7328__A2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7329__A (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7331__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7332__A (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7332__B (.DIODE(_0533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7333__A1 (.DIODE(_2695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7333__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7334__A (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7335__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7335__B2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7336__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7337__A1 (.DIODE(_0565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7337__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7339__A2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7339__B2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7339__C1 (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7340__A1 (.DIODE(_0571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7340__A2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7341__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7341__B (.DIODE(_0569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7342__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7343__A2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7343__B2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7343__C1 (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7344__A1 (.DIODE(_0574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7344__A2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7345__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7345__B (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7346__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7347__A (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7348__A (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7349__A (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7350__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7350__A2 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7350__B1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7350__B2 (.DIODE(net730));
 sky130_fd_sc_hd__diode_2 ANTENNA__7351__S (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7352__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7352__B (.DIODE(_0656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7353__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7354__A1 (.DIODE(_0619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7354__A2 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7354__B1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7354__B2 (.DIODE(_0675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7355__S (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7356__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7356__B (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7357__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7358__A (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7359__A (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7360__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7362__A (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7364__A (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7365__A1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7365__A2 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7365__B2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7366__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7367__A2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7367__B2 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7368__A (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7369__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7369__B2 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7370__A (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7371__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7371__A2 (.DIODE(_0688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7371__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7372__A (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7372__B (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7373__A (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7374__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7375__A (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7376__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7377__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7378__A (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7379__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7379__A2 (.DIODE(_0736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7379__B1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7380__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7381__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7382__A (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7383__A (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7383__B (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7384__A (.DIODE(_4235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7384__B (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7386__A2 (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7386__A3 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7386__B1 (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7387__A2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7388__A1 (.DIODE(_0710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7388__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7388__B2 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7389__A (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7390__A2 (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7390__B2 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7391__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7391__B2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7392__A1 (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7393__A1_N (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7393__B2 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7394__A (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7395__A1 (.DIODE(_0712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7395__A2 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7395__B2 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7396__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7397__A1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7397__A2 (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7397__B2 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7398__A (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7399__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7399__A2 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7399__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7400__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7401__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7402__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7403__A1 (.DIODE(_0797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7403__A2 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7403__B1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7403__C1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7404__A1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7404__A2 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7404__B1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7405__A2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7406__A1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7406__A2 (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7406__B2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7407__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7407__A2 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7407__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7408__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7409__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7410__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7411__A (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7412__A1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7412__A2 (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7412__B2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7413__A (.DIODE(_0788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7413__B (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7414__A2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7414__B2 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7415__A (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7416__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7416__B2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7417__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7417__A2 (.DIODE(_0854_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7417__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7418__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7419__A1_N (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7419__B1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7421__A2 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7421__B2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7422__A (.DIODE(_0784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7422__B (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7423__A2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7423__B2 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7425__A1 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7425__A2 (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7425__B2 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7426__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7426__A2 (.DIODE(_0885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7426__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7427__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7428__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7429__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7430__A1 (.DIODE(_0843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7430__A2 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7430__B1 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7430__C1 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7431__A (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7431__B (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7431__C (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7432__A (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7432__B (.DIODE(_0825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7433__A2 (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7433__B1 (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7435__A1_N (.DIODE(_0628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7435__A2_N (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7436__B (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7437__A1 (.DIODE(_0896_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7437__A2 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7438__A2 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7438__B2 (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7439__A (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7440__A2 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7440__B2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7441__A (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7442__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7442__B1 (.DIODE(_2794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7442__B2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7443__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7443__A2 (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7443__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7444__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7445__A1 (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7445__B1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7447__A (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7448__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7448__A2 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7448__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7450__A (.DIODE(_0931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7450__B (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7451__A (.DIODE(_0948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7451__B (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7452__A1 (.DIODE(_0904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7452__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7452__B1 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7452__C1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7453__A1 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7454__A2 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7454__B2 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7455__B1 (.DIODE(_0940_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7455__B2 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7456__A1 (.DIODE(_0957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7456__A2 (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7456__B2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7457__A1 (.DIODE(_0944_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7457__A2 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7457__B2 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7458__A2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7459__A (.DIODE(_0980_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7459__B (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7460__A1 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7461__A1 (.DIODE(_2810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7461__A2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7462__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7462__A2 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7462__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7463__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7464__A1 (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7464__A2 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7465__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7465__A2 (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7465__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7466__B (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7467__A2 (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7467__B2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7468__B (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7469__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7469__B1 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7470__A (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7470__B (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7471__A2 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7471__B1 (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7471__B2 (.DIODE(_2820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7472__B1 (.DIODE(_0986_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7472__B2 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7473__A2 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7473__B2 (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7474__A (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7475__A1 (.DIODE(_0973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7475__A2 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7475__B2 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7477__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7477__A2 (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7477__B2 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7478__A1 (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7478__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7480__A2 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7480__B2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7481__A1 (.DIODE(_0990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7481__A2 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7482__A1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7483__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7484__A1 (.DIODE(_1064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7484__A2 (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7484__B2 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7485__A1 (.DIODE(_1050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7485__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7487__A2 (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7487__B2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7487__C1 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7488__B (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7489__A1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7489__A2 (.DIODE(_1021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7489__B1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7490__A1 (.DIODE(_1077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7490__A2 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7492__A1 (.DIODE(_1067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7492__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7494__A1 (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7494__A2 (.DIODE(_1106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7494__B1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7495__A1 (.DIODE(_1052_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7495__A2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7495__B1 (.DIODE(_4184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7496__A2 (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7496__B2 (.DIODE(_0288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7498__B (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7499__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7500__A1_N (.DIODE(_1081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7500__A2_N (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7500__B1 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7501__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7501__B1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7501__B2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7502__A1 (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7502__B1 (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7503__A2 (.DIODE(_1111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7503__B1 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7504__A1 (.DIODE(_1071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7504__A2 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7504__B1 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7505__A (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7505__B (.DIODE(_2850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7506__A1 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7506__A2 (.DIODE(_1083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7508__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7509__B (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7510__B (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7512__A (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7513__A1 (.DIODE(_1090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7513__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7513__B1 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7514__B (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7515__A2 (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7515__A3 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7515__B1 (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7516__A1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7518__A1 (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7518__A2 (.DIODE(_1158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7518__B1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7519__A1_N (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7519__B1 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7519__B2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7520__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7521__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7522__A1 (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7522__A2 (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7522__B1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7523__A2 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7523__B2 (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7524__A (.DIODE(_0995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7524__B (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7525__A2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7525__B2 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7526__A (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7527__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7527__B1 (.DIODE(_2869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7527__B2 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7529__A (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7530__A1 (.DIODE(_4095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7531__B (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7532__A (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7532__B (.DIODE(_1180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7533__A2 (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7533__B1 (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7535__A1_N (.DIODE(_0997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7535__A2_N (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7536__B (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7537__A1 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7537__B1 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7538__A1 (.DIODE(_2878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7538__A2 (.DIODE(_2856_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7538__B1 (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7539__A2 (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7539__C1 (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7540__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7541__A2 (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7541__B2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7542__A (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7543__A2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7543__B2 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7544__A (.DIODE(_1215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7544__B (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7545__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7545__B1 (.DIODE(_2885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7545__B2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7546__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7546__A2 (.DIODE(_1232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7546__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7547__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7548__A1_N (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7548__B1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7550__A2 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7550__B2 (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7551__A (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7551__B (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7552__A2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7552__B2 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7553__A0 (.DIODE(_2893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7553__A1 (.DIODE(_1277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7553__S (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7554__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7554__A2 (.DIODE(_1256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7554__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7555__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7556__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7557__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7558__B (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7559__A1 (.DIODE(_1246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7559__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7559__B1 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7560__B (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7561__A2 (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7561__A3 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7561__B1 (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7562__A1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7563__B1 (.DIODE(_2899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7563__B2 (.DIODE(_2902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7564__A1 (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7564__A2 (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7564__B1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7565__A1_N (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7565__B1 (.DIODE(_1304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7565__B2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7566__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7567__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7568__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7569__A1 (.DIODE(_1260_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7569__A2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7569__B1 (.DIODE(_2231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7569__B2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7570__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7571__A1 (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7571__A2 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7571__B2 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7572__A1 (.DIODE(_1284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7572__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7574__A2 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7574__B2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7575__A (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7576__A1 (.DIODE(_1335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7576__A2 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7576__B2 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7577__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7578__A1 (.DIODE(_1301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7578__A2 (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7578__B1 (.DIODE(_2914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7578__B2 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7579__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7579__A2 (.DIODE(_1333_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7579__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7580__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7581__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7582__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7583__A2 (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7583__B2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7583__C1 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7584__B (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7585__A1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7585__A2 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7585__B1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7586__A1 (.DIODE(_1390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7586__A2 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7586__B2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7588__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7588__A2 (.DIODE(_1361_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7588__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7589__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7590__A (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7591__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7591__B1 (.DIODE(_2924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7592__B (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7593__A1 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7593__A2 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7593__B1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7594__A1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7594__A2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7594__B1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7595__B2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7596__A2 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7596__B2 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7596__C1 (.DIODE(_2931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7597__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7597__A2 (.DIODE(_1393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7597__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7598__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7599__A (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7600__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7601__A1 (.DIODE(_4094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7601__A2 (.DIODE(_1395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7601__B1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7602__A1 (.DIODE(_1436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7602__A2 (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7602__B1 (.DIODE(_1479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7602__B2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7602__C1 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7603__A1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7603__A2 (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7603__B1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7604__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7605__A1 (.DIODE(_1435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7605__A2 (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7607__A (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7608__A1 (.DIODE(_4095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7609__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7609__A2 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7609__B1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7610__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7611__B (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7612__A2 (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7612__A3 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7612__B1 (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7613__A1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7614__A1 (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7614__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7614__B1 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7615__A2 (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7615__B2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7616__A1 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7616__B1 (.DIODE(_2948_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7616__B2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7617__A1 (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7618__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7618__A2 (.DIODE(_1428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7618__B1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7619__B (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7620__B (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7621__A2 (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7621__A3 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7621__B1 (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7622__B (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7623__A (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7624__A2 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7625__A2 (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7625__B2 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7626__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7626__B1 (.DIODE(_2957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7626__B2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7627__A1 (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7628__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7628__A2 (.DIODE(_1462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7628__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7629__B (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7630__B (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7631__A2 (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7631__A3 (.DIODE(_2668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7631__B1 (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7632__A (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7633__A2 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7634__A1_N (.DIODE(_1535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7634__A2_N (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7634__B1 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7635__A1 (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7635__B1 (.DIODE(_2965_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7635__B2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7636__A1 (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7636__B1 (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7637__A (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7638__B (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7639__B (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7640__B (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7641__A1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7641__A2 (.DIODE(_1518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7641__B1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7642__A1 (.DIODE(_1564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7642__A2 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7642__B2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7644__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7644__A2 (.DIODE(_1539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7644__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7645__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7646__A (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7647__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7647__B1 (.DIODE(_2974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7648__A (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7649__A1 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7649__A2 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7649__B1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7650__A (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7652__A1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7652__A2 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7652__B1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7653__A1 (.DIODE(_1588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7653__A2 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7653__B2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7655__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7655__A2 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7655__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7656__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7657__A (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7658__A1 (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7658__B1 (.DIODE(_2984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7659__A2 (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7659__B2 (.DIODE(_2725_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7660__A (.DIODE(_1541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7660__B (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7661__A2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7661__B2 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7662__A1 (.DIODE(_1605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7662__A2 (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7662__B2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7663__A2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7664__A1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7664__A2 (.DIODE(_1594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7664__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7665__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7666__A1 (.DIODE(_2736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7666__B1 (.DIODE(_2685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7667__A1 (.DIODE(_2992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7668__B (.DIODE(_2768_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7669__A2 (.DIODE(_0056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7669__A3 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7669__B1 (.DIODE(_2745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7670__A1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7671__A2 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7671__B1 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7672__A (.DIODE(_2999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7672__B (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7673__A (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7674__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7674__A2 (.DIODE(_1636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7674__B1 (.DIODE(_0168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7675__A1 (.DIODE(_1601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7675__A2 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7676__A1 (.DIODE(_4095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7676__B2 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7678__B (.DIODE(_1621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7679__A1 (.DIODE(_1614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7679__A2 (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7679__B1 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7679__C1 (.DIODE(_2691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7680__B (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7681__A (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7682__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7683__A (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7683__B (.DIODE(_4095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7683__C (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7684__A2 (.DIODE(_2720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7684__B2 (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7685__A1_N (.DIODE(_2673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7685__B2 (.DIODE(_2671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7686__A (.DIODE(_2667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7687__A2 (.DIODE(_2724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7687__B2 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7688__A1_N (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7688__B1 (.DIODE(_1673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7688__B2 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7689__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7690__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7690__A2 (.DIODE(_1638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7690__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7691__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7692__A (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7693__A2 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7694__A (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7695__A1 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7695__A2 (.DIODE(_2666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7695__B1 (.DIODE(_1717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7695__B2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7696__A (.DIODE(_1670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7696__B (.DIODE(_2749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7697__A1 (.DIODE(_2680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7698__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7699__A1 (.DIODE(_2738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7699__A2 (.DIODE(_1681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7699__B1 (.DIODE(_2757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7700__B (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7701__A (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7702__A2 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7703__A1 (.DIODE(_1692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7703__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7703__B2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7703__C1 (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7704__A1 (.DIODE(_1703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7704__A2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7705__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7705__B (.DIODE(_1711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7706__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7707__A (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7707__B (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7707__C (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7707__D (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7708__A1 (.DIODE(_1735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7708__A2 (.DIODE(_2669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7708__B1 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7708__B2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7709__A1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7709__A2 (.DIODE(_2679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7710__A1 (.DIODE(_1742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7710__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7712__A1 (.DIODE(_2672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7712__B1 (.DIODE(_2710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7713__A1 (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7713__A2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7714__A2 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7715__A1 (.DIODE(_1753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7716__A1 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7716__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7718__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7718__B2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7718__C1 (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7719__A2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7720__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7720__B (.DIODE(_1762_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7721__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7722__A1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7722__A2 (.DIODE(_1793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7722__B1 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7723__B (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7724__A1 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7724__A2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7725__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7725__B (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7726__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7727__A1 (.DIODE(_1807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7727__A2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7727__B2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7727__C1 (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7728__A1 (.DIODE(_1816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7728__A2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7729__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7729__B (.DIODE(_1784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7730__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7731__A2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7731__B2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7731__C1 (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7732__A2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7733__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7734__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7735__A1 (.DIODE(_0229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7735__A2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7735__B1 (.DIODE(_2411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7735__B2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7735__C1 (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7736__A1 (.DIODE(_0131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7736__A2 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7737__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7737__B (.DIODE(_0191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7738__A1 (.DIODE(_3053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7738__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7739__A1 (.DIODE(_1836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7739__A2 (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7739__B2 (.DIODE(_2676_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7740__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7741__A1 (.DIODE(_1845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7741__S (.DIODE(_2686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7743__B (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7744__A1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7744__B1 (.DIODE(_2692_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7745__A2_N (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7746__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7747__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7748__A1 (.DIODE(_2711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7748__B1 (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7749__S (.DIODE(_2682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7750__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7751__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7752__A1 (.DIODE(_2742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7752__B1 (.DIODE(_2741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7752__C1 (.DIODE(_2674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7753__B (.DIODE(_2670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7754__A (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7755__A2 (.DIODE(_2700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7756__A (.DIODE(_2697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7756__B (.DIODE(_1885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7757__A2 (.DIODE(_2698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7758__A (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7758__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7760__A (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7761__A (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7762__A2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7762__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__7762__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7762__B2 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7763__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__7763__A2 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7763__B1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__7763__B2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7764__A1 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7764__A2 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7764__B1 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7764__B2 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__7765__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__7765__A2 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7765__B1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__7765__B2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7766__A (.DIODE(_4184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7766__B (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7767__A (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7767__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7769__A (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7770__A1 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7770__A2 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__7770__B1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__7770__B2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7771__A1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7771__A2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7771__B2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7773__A (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7773__B (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7774__A (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7775__A1 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7775__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7775__B1 (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7775__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7775__C1 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7776__A (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7778__A (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7779__A2 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7779__A3 (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA__7779__B1 (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA__7779__B2 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7780__A1 (.DIODE(net233));
 sky130_fd_sc_hd__diode_2 ANTENNA__7780__A2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7780__B1 (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA__7780__B2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7781__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7781__A2 (.DIODE(_3092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7781__B1_N (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7782__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7782__A2 (.DIODE(_3075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7783__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7783__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7783__B1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7783__B2 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__7784__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__7784__A2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7784__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__7784__B2 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7785__A1 (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7785__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7785__B1 (.DIODE(_4186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7785__B2 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__7786__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__7786__A2 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7786__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__7786__B2 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7787__A1 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7787__A2 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__7787__B1 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7787__B2 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__7788__A1 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__7788__A2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7788__B1 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7788__B2 (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7789__A1 (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7789__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7789__B1 (.DIODE(_3099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7789__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7789__C1 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7790__A1 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7790__A2 (.DIODE(net277));
 sky130_fd_sc_hd__diode_2 ANTENNA__7790__B1 (.DIODE(_0111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7790__B2 (.DIODE(net331));
 sky130_fd_sc_hd__diode_2 ANTENNA__7791__A1 (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA__7791__A2 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7791__B1 (.DIODE(net234));
 sky130_fd_sc_hd__diode_2 ANTENNA__7791__B2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7793__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7793__A2 (.DIODE(_3102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7793__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7794__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7794__A2 (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7795__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7795__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__7795__B1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7795__B2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__7796__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__7796__A2 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7796__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__7796__B2 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7797__A1 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7797__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__7797__B1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7797__B2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__7798__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__7798__A2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7798__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__7798__B2 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7799__A1 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7799__A2 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__7799__B1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__7799__B2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7800__A1 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__7800__A2 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7800__B1 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__7800__B2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7801__A1 (.DIODE(_3108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7801__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7801__B1 (.DIODE(_3110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7801__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7801__C1 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7802__A1 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7802__A2 (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA__7802__B1 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7802__B2 (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA__7803__A1 (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA__7803__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7803__B1 (.DIODE(net235));
 sky130_fd_sc_hd__diode_2 ANTENNA__7803__B2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7804__A1 (.DIODE(_3113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7804__A2 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7804__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7805__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7805__A2 (.DIODE(_3106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7806__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7806__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__7806__B1 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7807__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__7807__A2 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7807__B1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__7807__B2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7808__A1 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7808__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__7808__B1 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7809__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__7809__A2 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7809__B1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__7809__B2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7810__A1 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7810__B1 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__7810__B2 (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7811__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__7811__A2 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7811__B1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__7811__B2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7812__A1 (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7812__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7812__B1 (.DIODE(_3120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7812__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7812__C1 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7813__A1 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7813__A2 (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA__7813__B1 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7814__A1 (.DIODE(net236));
 sky130_fd_sc_hd__diode_2 ANTENNA__7814__A2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7814__B1 (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA__7814__B2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7815__A1 (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7815__A2 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7815__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7816__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7816__A2 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7817__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7817__B (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7818__A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA__7818__B (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7819__B1 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7820__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__7820__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7820__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7821__A (.DIODE(_3128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7822__A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7823__B (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7824__B1 (.DIODE(\arbiter.slave_sel[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7825__A1 (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__7825__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7825__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7827__A (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 ANTENNA__7829__A (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7829__B (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA__7830__B1 (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7831__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7831__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7833__A1 (.DIODE(_3133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7833__A2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7833__B1 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7833__B2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7833__C1 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7834__S (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7835__A (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7836__B (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7837__A2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7837__B2 (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7838__A1 (.DIODE(_3145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7838__A2 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7838__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7839__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7839__A2 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7842__A (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7842__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__7843__A (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7843__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__7844__B1 (.DIODE(\arbiter.slave_sel[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7845__A1 (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7845__A2 (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7845__B2 (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7846__A1 (.DIODE(_3152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7846__A2 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7846__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7847__A (.DIODE(_4114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7847__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__7848__A (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7848__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__7849__B1 (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7850__A1 (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7850__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7850__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7851__A (.DIODE(_3157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7852__A (.DIODE(_4253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7852__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__7853__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__7854__B1 (.DIODE(\arbiter.slave_sel[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7855__A1 (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7855__A2 (.DIODE(_4263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7855__B2 (.DIODE(_4287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7856__A (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7857__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7857__B1 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7857__C1 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7858__B (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA__7859__A (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7859__B (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA__7860__B1 (.DIODE(\arbiter.slave_sel[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__7861__A1 (.DIODE(_3147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7861__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7861__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7862__A (.DIODE(_3168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7863__B1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7866__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7866__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7866__B1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__7866__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7867__A2 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7867__B2 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7868__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7868__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7868__B1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__7868__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7869__A2 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7869__B2 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7870__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7870__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7870__B1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__7870__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7871__A2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7871__B2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7872__A (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7873__A1 (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7873__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7873__B1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7873__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7873__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7874__A (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7875__A (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7876__A (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7877__A1 (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 ANTENNA__7877__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7877__B1 (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA__7877__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7878__A2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7878__B2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7879__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7879__A2 (.DIODE(_3184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7879__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7880__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7880__A2 (.DIODE(_3173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7882__A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA__7883__A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA__7885__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7885__B1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7886__A1 (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7886__A2 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7886__B2 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7887__A1 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7887__B1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7888__A1 (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7888__A2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7888__B2 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7889__A1 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7889__B1 (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7889__B2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7890__A2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7890__B2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7891__A1 (.DIODE(_3193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7891__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7891__B1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7891__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7891__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7892__A1 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7893__A1 (.DIODE(_3186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7893__A2 (.DIODE(_0111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7893__B2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7894__A1 (.DIODE(_3198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7894__A2 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7894__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7895__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7895__A2 (.DIODE(_3191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7898__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7898__B1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__7899__A2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7899__B2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7900__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7900__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7900__B1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__7900__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7901__A2 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7901__B2 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7902__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7902__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7902__B1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__7902__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7903__A2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7903__B2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7904__A1 (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7904__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7904__B1 (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7904__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7904__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7905__A1 (.DIODE(net242));
 sky130_fd_sc_hd__diode_2 ANTENNA__7905__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7905__B1 (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA__7905__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7906__A2 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7906__B2 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7907__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7907__A2 (.DIODE(_3210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7907__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7908__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7908__A2 (.DIODE(_3203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7911__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7911__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7911__B1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__7911__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7912__A2 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7912__B2 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7913__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7913__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7913__B1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__7913__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7914__A2 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7914__B2 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7915__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7915__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7915__B1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__7915__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7916__A2 (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7916__B2 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7917__A1 (.DIODE(_3217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7917__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7917__B1 (.DIODE(_3219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7917__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7917__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7918__A1 (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA__7918__A2 (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7918__B1 (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA__7918__B2 (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7919__A2 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7919__B2 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7920__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7920__A2 (.DIODE(_3222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7920__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7921__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7921__A2 (.DIODE(_3215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7922__A (.DIODE(net241));
 sky130_fd_sc_hd__diode_2 ANTENNA__7924__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7924__B1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__7925__A2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7926__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7926__A2 (.DIODE(_4223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7926__B1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__7927__A2 (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7927__B2 (.DIODE(_4213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7928__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7928__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7928__B1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__7928__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7929__A2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7929__B2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7930__A1 (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7930__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7930__B1 (.DIODE(_3231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7930__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7930__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7931__A1 (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 ANTENNA__7931__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7931__B1 (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA__7931__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7932__A2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7932__B2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7933__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7933__A2 (.DIODE(_3234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7933__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7934__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7934__A2 (.DIODE(_3227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7937__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7937__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7937__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__7937__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7938__A2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7938__B2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7939__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7939__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7939__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__7939__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7940__A2 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7940__B2 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7941__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7941__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7941__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__7941__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7942__A2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7942__B2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7943__A1 (.DIODE(_3241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7943__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7943__B1 (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7943__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7943__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7944__A1 (.DIODE(net245));
 sky130_fd_sc_hd__diode_2 ANTENNA__7944__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7944__B1 (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA__7944__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7945__A2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7945__B2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7946__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7946__A2 (.DIODE(_3246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7946__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7947__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7947__A2 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7948__A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA__7950__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7950__B1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__7951__A2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7951__B2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7952__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7952__A2 (.DIODE(_4223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7952__B1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__7953__A2 (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7953__B2 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7955__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7955__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7955__B1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__7955__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7956__A2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7956__B2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7957__A1 (.DIODE(_3253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7957__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7957__B1 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7957__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7957__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7958__A1 (.DIODE(net246));
 sky130_fd_sc_hd__diode_2 ANTENNA__7958__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7958__B1 (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA__7958__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7959__A2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7959__B2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7960__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7960__A2 (.DIODE(_3259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7960__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7961__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7961__A2 (.DIODE(_3251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7964__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7964__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7964__B1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__7964__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7965__A2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7965__B2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7966__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7966__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7966__B1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__7966__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7967__A2 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7967__B2 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7968__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7968__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7968__B1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__7968__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7969__A2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7969__B2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7970__A1 (.DIODE(_3266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7970__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7970__B1 (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7970__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7970__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7971__A1 (.DIODE(net247));
 sky130_fd_sc_hd__diode_2 ANTENNA__7971__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7971__B1 (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA__7971__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7972__A2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7972__B2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7973__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7973__A2 (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7973__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7974__A1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7974__A2 (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7975__A (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7978__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7978__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7978__B1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__7978__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7979__A2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7979__B2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7980__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7980__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7980__B1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__7980__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7981__A2 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7981__B2 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7982__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7982__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7982__B1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__7982__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7983__A2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7983__B2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7984__A1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7984__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7984__B1 (.DIODE(_3281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7984__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7984__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7985__A1 (.DIODE(net248));
 sky130_fd_sc_hd__diode_2 ANTENNA__7985__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7985__B1 (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA__7985__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7986__A2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7986__B2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7987__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7987__A2 (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7987__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7988__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7988__A2 (.DIODE(_3277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7991__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__7991__B1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__7992__A2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7992__B2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7993__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__7993__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7993__B1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__7993__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7994__A2 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7994__B2 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7995__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__7995__A2 (.DIODE(_4263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7995__B1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__7995__B2 (.DIODE(_4287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7996__A2 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7996__B2 (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7997__A1 (.DIODE(_3291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7997__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7997__B1 (.DIODE(_3293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7997__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7997__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7998__A1 (.DIODE(net249));
 sky130_fd_sc_hd__diode_2 ANTENNA__7998__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7998__B1 (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA__7998__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7999__A2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__7999__B2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8000__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8000__A2 (.DIODE(_3296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8000__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8001__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8001__A2 (.DIODE(_3289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8004__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__8004__B1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__8005__A2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8006__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__8006__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8006__B1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__8006__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8007__A2 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8007__B2 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8008__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__8008__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8008__B1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__8008__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8009__A2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8009__B2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8010__A1 (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8010__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8010__B1 (.DIODE(_3305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8010__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8010__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8011__A1 (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA__8011__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8011__B1 (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA__8011__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8012__A2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8012__B2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8013__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8013__A2 (.DIODE(_3308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8013__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8014__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8014__A2 (.DIODE(_3301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8017__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__8017__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8017__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8018__A2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8018__B2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8019__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__8019__A2 (.DIODE(_4223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8020__A2 (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8020__B2 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8021__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__8021__A2 (.DIODE(_4263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8021__B2 (.DIODE(_4287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8022__A2 (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8022__B2 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8023__A1 (.DIODE(_3315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8023__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8023__B1 (.DIODE(_3317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8023__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8023__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8024__A1 (.DIODE(net251));
 sky130_fd_sc_hd__diode_2 ANTENNA__8024__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8024__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8025__A2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8025__B2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8026__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8026__A2 (.DIODE(_3320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8026__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8027__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8027__A2 (.DIODE(_3313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8028__A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA__8029__A (.DIODE(net350));
 sky130_fd_sc_hd__diode_2 ANTENNA__8032__A1 (.DIODE(_0192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8033__A2 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8034__A1 (.DIODE(_4204_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8034__B1 (.DIODE(_4213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8035__A2 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8035__B2 (.DIODE(_4186_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8037__A1 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8037__B2 (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8038__A2 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8038__B2 (.DIODE(_4265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8040__A1 (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8040__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8040__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8040__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8041__A1 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8041__B1 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8042__A2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8042__B2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8043__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8043__A2 (.DIODE(_3336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8043__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8044__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8044__A2 (.DIODE(_3327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8047__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__8047__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8047__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8048__A2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8048__B2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8049__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__8049__A2 (.DIODE(_4223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8050__A2 (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8050__B2 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8051__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__8051__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8051__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8052__A2 (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8052__B2 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8053__A1 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8053__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8053__B1 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8053__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8053__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8054__A1 (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA__8054__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8054__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8055__A2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8055__B2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8056__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8056__A2 (.DIODE(_3348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8056__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8057__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8057__A2 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8060__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__8060__B1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__8061__A2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8062__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__8062__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8062__B1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__8062__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8063__A2 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8063__B2 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8064__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__8064__A2 (.DIODE(_4263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8064__B1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__8064__B2 (.DIODE(_4287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8065__A2 (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8065__B2 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8066__A1 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8066__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8066__B1 (.DIODE(_3357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8066__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8066__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8067__A1 (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA__8067__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8067__B1 (.DIODE(net352));
 sky130_fd_sc_hd__diode_2 ANTENNA__8067__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8068__A2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8068__B2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8069__A1 (.DIODE(_3089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8069__A2 (.DIODE(_3360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8069__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8070__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8070__A2 (.DIODE(_3353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8073__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__8073__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8073__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8074__A2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8074__B2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8075__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__8075__A2 (.DIODE(_4223_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8076__A2 (.DIODE(_0910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8076__B2 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8077__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__8077__A2 (.DIODE(_4263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8077__B2 (.DIODE(_4287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8078__A2 (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8078__B2 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8079__A1 (.DIODE(_3367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8079__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8079__B1 (.DIODE(_3369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8079__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8079__C1 (.DIODE(_3178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8080__A1 (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA__8080__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8080__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8081__A2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8081__B2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8082__A2 (.DIODE(_3372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8082__B1_N (.DIODE(_3103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8083__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8083__A2 (.DIODE(_3365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8086__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__8086__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__8087__B2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8088__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__8088__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8088__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__8088__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8089__A2 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8089__B2 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8090__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__8090__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8090__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__8090__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8091__A2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8091__B2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8092__A1 (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8092__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8092__B1 (.DIODE(_3381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8092__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8092__C1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8093__A1 (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA__8093__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8093__B1 (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA__8093__B2 (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8094__A2 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8094__B2 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8095__A2 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__8096__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8096__A2 (.DIODE(_3377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8099__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__8099__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8099__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8100__A2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8100__B2 (.DIODE(_0741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8101__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__8101__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8102__A2 (.DIODE(_1894_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8102__B2 (.DIODE(_0538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8103__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__8103__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8103__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8104__A2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8104__B2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8105__A1 (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8105__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8105__B1 (.DIODE(_3393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8105__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8105__C1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8106__A1 (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA__8106__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8106__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8107__A2 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8107__B2 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8108__A2 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8109__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8109__A2 (.DIODE(_3389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8112__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__8112__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8112__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__8112__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8113__A2 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8113__B1 (.DIODE(_3399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8113__B2 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8114__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__8114__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8114__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__8114__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8115__A2 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8115__B1 (.DIODE(_3399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8115__B2 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8116__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__8116__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8116__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__8116__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8117__A2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8117__B1 (.DIODE(_3399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8117__B2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8118__A1 (.DIODE(_3403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8118__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8118__B1 (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8118__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8118__C1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8119__A1 (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA__8119__A2 (.DIODE(_3182_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8119__B1 (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 ANTENNA__8119__B2 (.DIODE(_3143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8120__A2 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8120__B1 (.DIODE(_3399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8120__B2 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8121__A2 (.DIODE(_3408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8122__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8122__A2 (.DIODE(_3401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8125__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__8125__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8125__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__8125__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8126__A2 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8126__B2 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8127__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__8127__A2 (.DIODE(_0678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8127__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__8127__B2 (.DIODE(_1133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8128__A2 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8128__B2 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8129__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__8129__A2 (.DIODE(_1291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8129__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__8129__B2 (.DIODE(_0614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8130__A2 (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8130__B2 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8131__A1 (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8131__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8131__B1 (.DIODE(_3417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8131__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8131__C1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8132__A1 (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA__8132__A2 (.DIODE(_0107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8132__B1 (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA__8132__B2 (.DIODE(_0160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8133__A2 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8133__B2 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8134__A2 (.DIODE(_3420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8135__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8135__A2 (.DIODE(_3413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8136__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__8136__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8136__B1 (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__8136__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8137__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__8137__A2 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8137__B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__8137__B2 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8138__A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__8139__A (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8140__A (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8140__B (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__8141__B (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8142__A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__8143__A (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8144__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__8144__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8146__A (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8147__A1 (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__8147__A2 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8147__B1 (.DIODE(_4245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8148__A1 (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__8148__A2 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8148__B1 (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA__8148__B2 (.DIODE(_4271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8149__A1 (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8149__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8149__B1 (.DIODE(_3434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8149__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8149__C1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8150__A (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8150__B (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA__8151__A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA__8151__B (.DIODE(_0730_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8152__A1_N (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA__8152__A2_N (.DIODE(_0844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8152__B2 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8153__A1 (.DIODE(\arbiter.slave_sel[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8154__A1 (.DIODE(_3439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8154__A2 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8154__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8155__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8155__A2 (.DIODE(_3423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8156__A1 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__8156__A2 (.DIODE(_0486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8156__B1 (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__8156__B2 (.DIODE(_0654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8157__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__8157__A2 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8157__B1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__8157__B2 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8158__A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA__8159__A (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8160__A (.DIODE(_4127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8160__B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__8161__B (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8162__A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__8163__A (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8164__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__8164__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8167__A1 (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8167__A2 (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__8167__B1 (.DIODE(_4245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8168__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__8168__A2 (.DIODE(_4272_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8168__B1 (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA__8168__B2 (.DIODE(_4271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8170__A1 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8170__A2 (.DIODE(_3450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8170__B1 (.DIODE(_3454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8170__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8170__C1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8171__A (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8172__A (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8172__B (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA__8173__B (.DIODE(\arbiter.slave_sel[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8174__A (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8175__A1 (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA__8175__A2 (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8176__A1 (.DIODE(_3460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8176__A2 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8176__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8177__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8177__A2 (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8178__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__8178__B (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8180__A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__8181__A (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8182__B1 (.DIODE(\arbiter.slave_sel[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8183__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__8183__A2 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8183__B2 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8184__A1 (.DIODE(_3467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8184__A2 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8184__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8185__B (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8186__A1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8186__A2 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__8187__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__8187__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8188__A0 (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA__8188__A1 (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__8188__S (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8189__A (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8189__B (.DIODE(_4245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8189__C (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__8190__A2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8190__B2 (.DIODE(\arbiter.slave_sel[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8191__A1 (.DIODE(_3471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8191__A2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8191__B1 (.DIODE(_3474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8191__B2 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8191__C1 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8192__A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA__8192__B (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8194__A (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8195__B1 (.DIODE(\arbiter.slave_sel[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8196__A1 (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA__8196__A2 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8196__B2 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8197__B1 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8197__B2 (.DIODE(_3480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8198__B (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__8199__A1 (.DIODE(_0198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8199__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__8199__B1 (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8200__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__8200__A2 (.DIODE(_0888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8200__B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__8200__B2 (.DIODE(_0197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8201__A1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8201__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__8201__B1 (.DIODE(_4119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8202__A1 (.DIODE(_0522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8202__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__8203__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__8203__A2 (.DIODE(_0520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8203__B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__8204__A1 (.DIODE(_4253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8204__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__8204__B1 (.DIODE(_4245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8205__A1 (.DIODE(_0510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8205__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__8206__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__8206__A2 (.DIODE(_0785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8206__B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__8206__B2 (.DIODE(_4271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8207__A1 (.DIODE(_3486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8207__A2 (.DIODE(_3254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8207__B1 (.DIODE(_3489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8207__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8207__C1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8208__A1 (.DIODE(_0090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8208__A2 (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA__8208__B1 (.DIODE(_0096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8209__A1 (.DIODE(_0088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8209__A2 (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA__8210__A1 (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA__8210__A2 (.DIODE(_0152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8210__B1 (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA__8210__B2 (.DIODE(_0110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8211__A (.DIODE(_3493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8212__A2 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8212__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8213__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8213__A2 (.DIODE(_3483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8214__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8214__B1 (.DIODE(_0651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8214__B2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__8215__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__8215__A2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8215__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__8215__B2 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8216__A1 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8216__B1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8216__B2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__8217__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__8217__A2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8217__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__8217__B2 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8218__A1 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8218__A2 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__8218__B1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__8218__B2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8219__A1 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__8219__A2 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8219__B2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8220__A1 (.DIODE(_3499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8220__B1 (.DIODE(_3501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8220__B2 (.DIODE(_3134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8220__C1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8221__A1 (.DIODE(_0759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8221__B1 (.DIODE(_0143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8221__B2 (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA__8222__A1 (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA__8222__A2 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8222__B1 (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA__8222__B2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8223__A2 (.DIODE(_3504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8224__A1 (.DIODE(_3273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8224__A2 (.DIODE(_3497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8225__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8225__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__8225__B1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8225__B2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__8226__A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__8226__A2 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8226__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__8226__B2 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8227__A1 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8227__A2 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__8227__B1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__8227__B2 (.DIODE(_0612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8228__A1 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8228__A2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__8228__B1 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__8228__B2 (.DIODE(_4278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8231__A1 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8231__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__8231__B1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8231__B2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__8232__A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__8232__A2 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8232__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__8232__B2 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8233__A1 (.DIODE(_3084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8233__A2 (.DIODE(_3511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8233__B1 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8233__B2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8233__C1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8234__A1 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8234__A2 (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA__8234__B1 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8234__B2 (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA__8235__A1 (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA__8235__A2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8235__B1 (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA__8235__B2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8236__A1 (.DIODE(_3516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8236__A2 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8236__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8237__A1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8237__A2 (.DIODE(_3507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8238__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8238__A2 (.DIODE(_3086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8238__B1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8239__A (.DIODE(_4145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8240__A (.DIODE(_4286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8241__A1 (.DIODE(_3519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8241__B1 (.DIODE(_3520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8241__C1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8242__B1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8242__B2 (.DIODE(_3072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8243__A1 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8243__B1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8243__B2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__8244__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__8244__A2 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8244__B1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__8244__B2 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8245__A1 (.DIODE(_4268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8245__A2 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__8245__B1 (.DIODE(_4280_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8245__B2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__8246__A2 (.DIODE(_3081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8246__B1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__8246__B2 (.DIODE(_0613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8248__A1 (.DIODE(_0539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8248__B1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8248__B2 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__8249__A1 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__8249__A2 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8249__B1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__8249__B2 (.DIODE(_0590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8250__A1 (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8250__B1 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8250__B2 (.DIODE(_3080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8250__C1 (.DIODE(_3085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8251__A1 (.DIODE(_3180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8251__B1 (.DIODE(_3181_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8251__B2 (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA__8252__A1 (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 ANTENNA__8252__A2 (.DIODE(_0572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8252__B1 (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA__8252__B2 (.DIODE(_0108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8253__A2 (.DIODE(_3531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8254__A1 (.DIODE(_3071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8254__A2 (.DIODE(_3523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8255__A2 (.DIODE(_3504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8255__B1 (.DIODE(_3092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8256__B (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8257__B (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8257__C (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8258__A (.DIODE(_3535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8260__A1 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8260__A2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8260__B1 (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8260__B2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8261__B (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8262__S (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8263__A2 (.DIODE(_3497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8263__B1 (.DIODE(_3075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8263__B2 (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8264__A (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8264__B (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8265__A (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8266__S (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8268__A (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8270__A (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8271__A (.DIODE(_0637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8271__B (.DIODE(_0454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8272__A (.DIODE(_3102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8273__A1 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8273__A2 (.DIODE(_3516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8273__B1 (.DIODE(_3548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8274__A2 (.DIODE(_3511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8274__B1 (.DIODE(_3099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8275__A1 (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8275__A2 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8275__B1 (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8275__B2 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8276__A1 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8276__B2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8276__C1 (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8277__A1 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8278__A1 (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8278__S (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8280__A1 (.DIODE(_3108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8280__A2 (.DIODE(_3535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8280__B1 (.DIODE(_3110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8280__B2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8281__A1 (.DIODE(_3113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8281__A2 (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8282__A1 (.DIODE(_3106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8282__S (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8284__B (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8285__A1 (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8285__A2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8285__B1 (.DIODE(_3120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8285__B2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8285__C1 (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8286__A1 (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8287__A1 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8287__S (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8288__A (.DIODE(_3562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8289__A (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8290__A (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8290__B (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8291__A (.DIODE(_3564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8292__A1 (.DIODE(_3075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8292__B1 (.DIODE(_3565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8293__A1 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8293__A2 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8293__B1 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8293__B2 (.DIODE(_3106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8294__A (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8295__A (.DIODE(_3092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8296__A2 (.DIODE(_3113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8296__B1 (.DIODE(_3145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8297__A2 (.DIODE(_3548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8298__A1 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8298__A2 (.DIODE(_3571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8298__B1 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8299__A (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8300__A (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8302__A1 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8302__A2 (.DIODE(\arbiter.master_sel[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8303__A1 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8303__A2 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8303__B1 (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8303__B2 (.DIODE(_3108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8304__A (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8305__A1 (.DIODE(_3133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8305__A2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8305__B1 (.DIODE(_3577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8305__B2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8306__B (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8307__A1 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8308__A1 (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8308__A2 (.DIODE(\arbiter.master_sel[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8309__A1 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8309__B1 (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8309__B2 (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8310__A (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8310__B (.DIODE(_0412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8311__A (.DIODE(_3583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8312__A1 (.DIODE(_3099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8313__A1 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8313__B1 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8313__B2 (.DIODE(_3120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8314__A1 (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8314__A2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8314__B1 (.DIODE(_3586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8314__B2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8315__A (.DIODE(_3152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8316__B (.DIODE(_3548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8317__A1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8318__A1 (.DIODE(_3590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8318__S (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8319__A1 (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8319__B1 (.DIODE(_3565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8320__A1 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8320__B1 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8320__B2 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8321__A1 (.DIODE(_3593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8321__S (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8323__A (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8324__A1 (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8324__A2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8324__B1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8324__B2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8324__C1 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8325__A1 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8325__A2 (.DIODE(_3184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8325__B1 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8326__A1 (.DIODE(_3173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8326__A2 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8327__A1 (.DIODE(_3193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8327__A2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8327__B1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8327__B2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8327__C1 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8328__A1 (.DIODE(_3198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8328__A2 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8328__B1 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8329__A1 (.DIODE(_3191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8329__A2 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8330__A1 (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8330__A2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8330__B1 (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8330__B2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8330__C1 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8331__A1 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8331__A2 (.DIODE(_3210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8331__B1 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8332__A1 (.DIODE(_3203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8332__A2 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8333__A (.DIODE(_3198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8334__A (.DIODE(_3602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8334__B (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8335__A (.DIODE(_3222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8335__B (.DIODE(_0450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8338__A1 (.DIODE(_3217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8338__A2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8338__B1 (.DIODE(_3219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8338__B2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8339__A1 (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8340__A1 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8340__A2 (.DIODE(_3191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8340__B1 (.DIODE(_3215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8341__S (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8343__A1 (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8343__A2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8343__B1 (.DIODE(_3231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8343__B2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8343__C1 (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8344__A1 (.DIODE(_3234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8344__A2 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8345__A (.DIODE(_3227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8345__B (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8346__A (.DIODE(_3203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8346__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8347__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8349__A (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8350__A2 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8351__A (.DIODE(_3241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8351__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8352__A (.DIODE(_3217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8352__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8353__S (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8355__A1 (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8355__A2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8355__B2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8355__C1 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8356__A1 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8356__A2 (.DIODE(_3246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8356__B1 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8357__A1 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8357__A2 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8358__A (.DIODE(_3253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8358__B (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8359__A (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8359__B (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8360__S (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8362__A1 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8362__A2 (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8363__A1 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8363__A2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8363__B1 (.DIODE(_3628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8363__B2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8364__A (.DIODE(_3548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8365__A1 (.DIODE(_3210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8366__A1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8366__A2 (.DIODE(_3259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8366__B1 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8366__B2 (.DIODE(_3234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8367__A1 (.DIODE(_3632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8367__S (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8368__A (.DIODE(_0475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8369__A (.DIODE(_3251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8369__B (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8370__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8372__A2 (.DIODE(_3203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8372__B2 (.DIODE(_3565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8373__A1 (.DIODE(_3638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8373__S (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8375__A (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8375__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8376__A (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8376__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8377__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8379__A2 (.DIODE(_3215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8379__B2 (.DIODE(_3565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8380__A1 (.DIODE(_0453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8380__A2 (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8380__B1 (.DIODE(_0457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8380__B2 (.DIODE(_3246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8382__A1 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8382__A2 (.DIODE(_3646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8382__B1 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8383__A1 (.DIODE(_3219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8384__A1 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8384__A2 (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8384__B1 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8384__B2 (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8385__A2 (.DIODE(_3217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8385__B1 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8386__A1 (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8386__A2 (.DIODE(_3241_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8386__B1 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8386__B2 (.DIODE(_3266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8387__A1 (.DIODE(_3649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8387__A2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8387__B1 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8387__B2 (.DIODE(_3651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8388__B (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8389__A1 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8389__A2 (.DIODE(_3644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8390__A (.DIODE(_3277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8390__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8391__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8393__S (.DIODE(_3564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8394__A (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8394__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8395__S (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8396__B1 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8396__B2 (.DIODE(_3229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8397__A1 (.DIODE(_3281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8397__A2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8397__B2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8397__C1 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8398__A1 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8398__A2 (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8398__B1 (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8399__A1 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8400__A (.DIODE(_3289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8400__B (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8401__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8402__A1_N (.DIODE(_3564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8402__B2 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8403__A (.DIODE(_3291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8403__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8404__A (.DIODE(_3266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8404__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8405__S (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8409__A1 (.DIODE(_3293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8409__A2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8409__B2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8409__C1 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8410__A1 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8410__A2 (.DIODE(_3296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8410__B1 (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8411__A1 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8412__A (.DIODE(_3301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8412__B (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8413__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8415__A1 (.DIODE(_3564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8416__A (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8416__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8417__S (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8420__A1 (.DIODE(_3305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8420__A2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8420__B2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8420__C1 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8421__A1 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8421__A2 (.DIODE(_3308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8421__B1 (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8422__A1 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8423__A (.DIODE(_3317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8423__B (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8424__A (.DIODE(_3293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8424__B (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8427__A (.DIODE(_3315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8427__B (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8428__S (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8429__A (.DIODE(_3535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8431__A2 (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8432__A1 (.DIODE(_3320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8432__S (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8433__A (.DIODE(_3313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8433__B (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8434__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8436__A1 (.DIODE(_3564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8437__S (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8438__A (.DIODE(_3698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8439__A (.DIODE(_3327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8439__B (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8440__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8442__A1 (.DIODE(_3564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8443__A1 (.DIODE(_3336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8443__A2 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8443__B1 (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8444__A (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8445__A (.DIODE(_3704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8446__S (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8449__A (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8450__A1 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8451__A (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8451__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8452__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8453__B (.DIODE(_3565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8454__B (.DIODE(_3564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8455__A (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8455__B (.DIODE(_0426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8456__S (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8458__A (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8458__B (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8461__A2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8461__B2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8461__C1 (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8462__A1 (.DIODE(_3348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8462__A2 (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8462__B1 (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8463__A1 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8464__A (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8464__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8465__S (.DIODE(\arbiter.master_sel[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8467__B1 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8468__B (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8469__A (.DIODE(_3357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8469__B (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8472__A2 (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8472__B1 (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8473__A1 (.DIODE(_3360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8473__A2 (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8474__A1 (.DIODE(_3353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8474__S (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8475__A (.DIODE(_3732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8476__A (.DIODE(_3365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8476__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8477__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8478__S (.DIODE(_3564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8480__A (.DIODE(_3369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8480__B (.DIODE(_0615_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8483__A (.DIODE(_3367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8483__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8484__S (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8487__A1 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8487__B2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8487__C1 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8488__A1 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8488__A2 (.DIODE(_3372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8488__B1 (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8489__A1 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8490__A (.DIODE(_3377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8490__B (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8491__A (.DIODE(_3353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8491__B (.DIODE(_0646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8492__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8493__S (.DIODE(_3565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8495__A1 (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8495__A2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8495__B1 (.DIODE(_3381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8495__B2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8496__A1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__8496__S (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8497__S (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8498__A (.DIODE(_3753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8499__A (.DIODE(_3389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8499__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8500__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8501__S (.DIODE(_3564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8503__A (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8503__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8504__S (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8507__A1 (.DIODE(_3393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8507__A2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8507__B2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8507__C1 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8508__A1 (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8508__A2 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8508__B1 (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8509__A1 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8510__A (.DIODE(_3403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8510__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8511__A (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8511__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8512__S (.DIODE(_4153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8514__A1 (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8514__A2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8514__B2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8514__C1 (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8515__A (.DIODE(_3408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8515__B (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8516__A (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__8516__B (.DIODE(_0451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8518__B (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8519__A (.DIODE(_3401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8519__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8520__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8521__A2 (.DIODE(_3565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8521__B1 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8522__A2 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8523__A (.DIODE(_3413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8523__B (.DIODE(_0469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8524__S (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8525__A (.DIODE(_3777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8526__A1 (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8526__A2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8526__B1 (.DIODE(_3417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8526__B2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8526__C1 (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8527__A1 (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8527__A2 (.DIODE(_3420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8527__B1 (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8528__A1 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8529__A1 (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8529__A2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8529__B1 (.DIODE(_3434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8529__B2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8529__C1 (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8530__A1 (.DIODE(_3439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8530__A2 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8530__B1 (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8531__A1 (.DIODE(_3423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8531__A2 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8532__A1 (.DIODE(_3450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8532__A2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8532__B1 (.DIODE(_3454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8532__B2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8532__C1 (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8533__A1 (.DIODE(_3460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8533__A2 (.DIODE(_3547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8533__B1 (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8534__A1 (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8534__A2 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8535__B (.DIODE(_3564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8536__A1 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8536__A2 (.DIODE(_3480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8536__B1 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8536__B2 (.DIODE(_3423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8537__A2 (.DIODE(_3467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8537__B1 (.DIODE(_3439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8538__A2 (.DIODE(_3548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8539__A1 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8539__B1 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8541__A1 (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8541__A2 (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8541__B1 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8541__B2 (.DIODE(_3471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8542__A1 (.DIODE(_3474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8542__A2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8542__B2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8543__B (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8544__A1 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8545__A1 (.DIODE(_3420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8546__A2 (.DIODE(_3460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8548__A1 (.DIODE(_3417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8549__A1 (.DIODE(_0414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8549__A2 (.DIODE(_3454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8549__B1 (.DIODE(_0410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8549__B2 (.DIODE(_3489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8550__A (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8550__B (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8552__A1 (.DIODE(_0253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8552__A2 (.DIODE(_3450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8552__B1 (.DIODE(_0431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8552__B2 (.DIODE(_3486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8553__A2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8553__B2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8554__A1 (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8555__A (.DIODE(_3777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8555__B (.DIODE(_3564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8556__A1 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8556__A2 (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8556__B1 (.DIODE(_0473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8556__B2 (.DIODE(_3483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8557__S (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8559__A1 (.DIODE(_3499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8559__A2 (.DIODE(_3578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8559__B1 (.DIODE(_3501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8559__B2 (.DIODE(_3573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8559__C1 (.DIODE(_3546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8560__A1 (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8560__A2 (.DIODE(_3504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8560__B1 (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8561__A1 (.DIODE(_3497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8561__A2 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8562__A1 (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8562__A2 (.DIODE(_3516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8562__B1 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8563__A1 (.DIODE(_3511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8563__A2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8563__B1 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8563__B2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8564__B (.DIODE(_3568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8565__A1 (.DIODE(_3507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8565__A2 (.DIODE(_3563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8566__A1 (.DIODE(_3519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8566__A2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8566__B1 (.DIODE(_3520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8566__B2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8567__B (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8568__A1 (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8568__A2 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8568__B1 (.DIODE(_3542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8569__A1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8569__A2 (.DIODE(_3595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8570__A1 (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8570__A2 (.DIODE(_3537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8570__B1 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8570__B2 (.DIODE(_3536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8571__A1 (.DIODE(_3531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8571__A2 (.DIODE(_3539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8572__A1 (.DIODE(_3523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8572__S (.DIODE(_3543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8574__B (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8575__A (.DIODE(_3818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8577__A (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8578__B (.DIODE(_4233_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8579__B (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8579__C (.DIODE(_0436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8581__A (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8583__A (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8584__B (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8587__A (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8588__A1 (.DIODE(_3077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8588__A2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8588__B1 (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8588__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8590__A (.DIODE(_3818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8591__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8591__A2 (.DIODE(_3092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8591__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8592__A1 (.DIODE(_3075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8592__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8593__A1 (.DIODE(_3097_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8593__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8593__B1 (.DIODE(_3099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8593__B2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8594__A1 (.DIODE(_3102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8594__S (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8595__A1 (.DIODE(_3095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8595__S (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8597__A1 (.DIODE(_3110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8597__A2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8597__B1 (.DIODE(_3577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8597__B2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8598__A1 (.DIODE(_3571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8598__B1 (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8599__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8600__A1 (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8600__A2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8600__B1 (.DIODE(_3586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8600__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8601__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8601__A2 (.DIODE(_3590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8601__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8602__A1 (.DIODE(_3593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8602__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8603__A1 (.DIODE(_3133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8603__A2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8603__B1 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8603__B2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8604__A1 (.DIODE(_3145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8604__B1 (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8605__A1 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8605__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8606__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8606__B2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8608__S (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8610__A1 (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8610__A2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8610__B1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8610__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8611__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8611__A2 (.DIODE(_3184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8611__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8612__A1 (.DIODE(_3173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8612__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8613__A1 (.DIODE(_3193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8613__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8613__B1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8613__B2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8614__A1 (.DIODE(_3602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8614__S (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8615__A1 (.DIODE(_3191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8615__S (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8617__A1 (.DIODE(_3205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8617__A2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8617__B1 (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8617__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8618__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8618__A2 (.DIODE(_3210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8618__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8619__A1 (.DIODE(_3203_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8619__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8620__A1 (.DIODE(_3217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8620__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8620__B1 (.DIODE(_3219_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8620__B2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8621__A1 (.DIODE(_3222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8621__S (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8622__A1 (.DIODE(_3215_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8622__S (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8624__A1 (.DIODE(_3231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8624__A2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8624__B1 (.DIODE(_3628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8624__B2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8625__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8625__A2 (.DIODE(_3632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8625__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8626__A1 (.DIODE(_3638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8626__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8627__A1 (.DIODE(_3649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8627__A2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8627__B1 (.DIODE(_3651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8627__B2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8628__A1 (.DIODE(_3646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8628__B1 (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8629__A1 (.DIODE(_3644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8629__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8630__A1 (.DIODE(_3253_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8630__A2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8630__B1 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8630__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8631__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8631__A2 (.DIODE(_3259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8631__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8632__A1 (.DIODE(_3251_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8632__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8633__A1 (.DIODE(_3266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8633__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8633__B1 (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8633__B2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8634__A1 (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8635__A1 (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8637__A1 (.DIODE(_3279_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8637__A2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8637__B1 (.DIODE(_3281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8637__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8637__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8638__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8638__A2 (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8638__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8639__A1 (.DIODE(_3277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8639__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8640__A1 (.DIODE(_3291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8640__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8640__B2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8641__A1 (.DIODE(_3296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8642__A1 (.DIODE(_3289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8644__A1 (.DIODE(_3303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8644__A2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8644__B1 (.DIODE(_3305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8644__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8644__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8645__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8645__A2 (.DIODE(_3308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8645__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8646__A1 (.DIODE(_3301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8646__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8647__B1 (.DIODE(_3315_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8647__B2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8648__A1 (.DIODE(_3320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8649__A1 (.DIODE(_3313_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8651__A1 (.DIODE(_3330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8651__A2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8651__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8651__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8652__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8652__A2 (.DIODE(_3336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8652__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8653__A1 (.DIODE(_3327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8653__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8654__B1 (.DIODE(_3343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8654__B2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8655__A1 (.DIODE(_3348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8656__A1 (.DIODE(_3341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8658__A1 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8658__A2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8658__B1 (.DIODE(_3357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8658__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8658__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8659__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8659__A2 (.DIODE(_3360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8659__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8660__A1 (.DIODE(_3353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8660__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8661__A1 (.DIODE(_3367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8661__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8661__B1 (.DIODE(_3369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8661__B2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8662__A1 (.DIODE(_3372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8663__A1 (.DIODE(_3365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8665__A1 (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8665__A2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8665__B1 (.DIODE(_3381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8665__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8665__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8666__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8666__A2 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__8666__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8667__A1 (.DIODE(_3377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8667__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8668__A1 (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8668__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8668__B1 (.DIODE(_3393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8668__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8668__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8669__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8669__A2 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8669__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8670__A1 (.DIODE(_3389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8670__A2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8671__A1 (.DIODE(_3403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8671__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8671__B1 (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8671__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8671__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8672__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8672__A2 (.DIODE(_3408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8672__B1 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8673__A1 (.DIODE(_3401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8673__A2 (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8674__A1 (.DIODE(_3415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8674__B1 (.DIODE(_3417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8674__B2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8675__A1 (.DIODE(_3420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8676__A1 (.DIODE(_3413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8678__A1 (.DIODE(_3434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8678__A2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8678__B2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8678__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8679__B1 (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8680__A2 (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8681__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8681__B2 (.DIODE(_3827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8681__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8682__B1 (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8683__A2 (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8684__A1 (.DIODE(_3471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8684__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8684__B1 (.DIODE(_3474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8684__B2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8684__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8685__A (.DIODE(_3467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8686__A (.DIODE(_3480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8686__B (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8687__A2 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8688__A1 (.DIODE(_3486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8688__B1 (.DIODE(_3489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8688__B2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8689__A1 (.DIODE(_3493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8690__A1 (.DIODE(_3483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8692__A1 (.DIODE(_3499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8692__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8692__B1 (.DIODE(_3501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8692__B2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8693__A2 (.DIODE(_4239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8693__B1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8694__A1 (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8694__B2 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8695__A1 (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8695__B1 (.DIODE(_3818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8697__A2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8697__A3 (.DIODE(\arbiter.master_sel[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__8698__B (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8699__B1 (.DIODE(_3507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8699__B2 (.DIODE(_3834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8700__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8700__B1 (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8701__A1 (.DIODE(_3519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8701__A2 (.DIODE(_3824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8701__B1 (.DIODE(_3520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8701__B2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8701__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8702__B1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8702__B2 (.DIODE(_3821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8703__A1 (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8703__A2 (.DIODE(_3826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8703__B1 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8703__B2 (.DIODE(_3825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8703__C1 (.DIODE(_3830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8704__A1 (.DIODE(_3833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8704__A2 (.DIODE(_3531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8704__B1 (.DIODE(_3818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8705__A1 (.DIODE(_3523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8705__A2 (.DIODE(_3820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8706__A (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8706__B (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8708__A (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8709__A (.DIODE(_4184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8709__B (.DIODE(_0625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8713__B (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8713__C (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8716__A (.DIODE(_0083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8716__B (.DIODE(_0455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8717__A (.DIODE(_3926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8718__A1 (.DIODE(_3083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8718__A2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8718__B1 (.DIODE(_3577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8718__B2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8718__C1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8719__A1 (.DIODE(_3571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8719__A2 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8719__B1 (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8720__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8721__A1 (.DIODE(_3582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8721__A2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8721__B1 (.DIODE(_3586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8721__B2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8721__C1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8722__A (.DIODE(_3926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8726__A2 (.DIODE(_3590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8727__A1 (.DIODE(_3593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8727__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8728__A1 (.DIODE(_3108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8728__A2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8728__B1 (.DIODE(_3110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8728__B2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8728__C1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8729__A1 (.DIODE(_3113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8729__A2 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8729__B1 (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8730__A1 (.DIODE(_3106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8730__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8731__A2 (.DIODE(_3123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8732__A1 (.DIODE(_3118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8732__B1 (.DIODE(_3120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8734__A1 (.DIODE(_3116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8735__A1 (.DIODE(_3133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8735__A2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8735__B1 (.DIODE(_3140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8735__B2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8735__C1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8736__A1 (.DIODE(_3145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8736__A2 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8736__B1 (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8737__A1 (.DIODE(_3129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8737__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8739__A2 (.DIODE(_3162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8739__B1 (.DIODE(_3157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8740__A1 (.DIODE(_3152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8740__A2 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8740__B1 (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8741__A1 (.DIODE(_3168_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8742__A1 (.DIODE(_3175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8742__A2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8742__B1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8742__B2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8742__C1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8743__A2 (.DIODE(_3184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8744__A1 (.DIODE(_3173_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8744__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8745__A1 (.DIODE(_3193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8745__B1 (.DIODE(_3195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8745__C1 (.DIODE(_3926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8746__A1 (.DIODE(_3602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8747__A1 (.DIODE(_3191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8747__S (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8749__A1 (.DIODE(_3207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8749__A2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8749__B1 (.DIODE(_3628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8749__B2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8749__C1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8750__A2 (.DIODE(_3632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8751__A1 (.DIODE(_3638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8751__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8752__A1 (.DIODE(_3649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8752__A2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8752__B1 (.DIODE(_3651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8752__B2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8752__C1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8753__A1 (.DIODE(_3646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8753__A2 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8753__B1 (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8754__A1 (.DIODE(_3644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8754__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8755__C (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8756__A1 (.DIODE(_3231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8756__C1 (.DIODE(_3926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8757__A1 (.DIODE(_3234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8758__A1 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8758__A2 (.DIODE(_3227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8758__A3 (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8759__A (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8759__B (.DIODE(_3565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8760__A1 (.DIODE(_3243_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8761__A (.DIODE(_3926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8762__A1 (.DIODE(_3246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8762__S (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8764__A1 (.DIODE(_3256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8764__C1 (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8765__B (.DIODE(_3259_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8767__A1 (.DIODE(_3266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8767__A2 (.DIODE(_0427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8767__B1 (.DIODE(_3268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8768__A1 (.DIODE(_3271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8768__S (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8771__A1 (.DIODE(_3281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8771__B1 (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8772__B (.DIODE(_3284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8774__A1 (.DIODE(_3293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8774__A2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8774__B2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8774__C1 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8775__A2 (.DIODE(_3296_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8776__A1 (.DIODE(_3289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8776__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8777__A1 (.DIODE(_3305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8777__B1 (.DIODE(_3926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8778__A2 (.DIODE(_0589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8778__A3 (.DIODE(_0433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8779__A2 (.DIODE(_3308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8780__A1 (.DIODE(_3301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8780__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8781__A1 (.DIODE(_3317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8781__C1 (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8782__B (.DIODE(_3320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8784__A1 (.DIODE(_3704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8785__A1 (.DIODE(_3336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8785__S (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8787__A1 (.DIODE(_3345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8788__A1 (.DIODE(_3348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8788__S (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8790__A1 (.DIODE(_3355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8790__A2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8790__B1 (.DIODE(_3357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8790__B2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8790__C1 (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8791__A2 (.DIODE(_3360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8792__A1 (.DIODE(_3353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8792__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8793__A1 (.DIODE(_3367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8793__B1 (.DIODE(_3369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8794__A1 (.DIODE(_3372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8794__S (.DIODE(_3926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8795__A1 (.DIODE(_3365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8795__S (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8797__A1 (.DIODE(_3379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8797__A2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8797__B1 (.DIODE(_3381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8797__B2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8797__C1 (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8798__A2 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__8799__A1 (.DIODE(_3377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8799__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8800__A1 (.DIODE(_3391_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8800__A2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8800__B1 (.DIODE(_3393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8800__B2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8800__C1 (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8801__A2 (.DIODE(_3396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8802__A1 (.DIODE(_3389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8802__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8803__B (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8804__A1 (.DIODE(_3405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8804__A2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8804__B1 (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8805__A2 (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8806__B (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8807__A1 (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8809__S (.DIODE(_3926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8810__S (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8811__A (.DIODE(_3995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8812__A1 (.DIODE(_3431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8812__A2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8812__B1 (.DIODE(_3434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8812__B2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8812__C1 (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8813__A1 (.DIODE(_3439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8813__A2 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8813__B1 (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8814__A1 (.DIODE(_3423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8814__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8815__A2 (.DIODE(_3460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8816__A1 (.DIODE(_3450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8816__B1 (.DIODE(_3454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8818__A1 (.DIODE(_3442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8819__A1 (.DIODE(_3471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8819__A2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8819__B1 (.DIODE(_3474_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8819__B2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8819__C1 (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8820__A (.DIODE(_3467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8820__B (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8821__A (.DIODE(_3480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8821__B (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8823__A1 (.DIODE(_3486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8823__B1 (.DIODE(_3489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8824__A1 (.DIODE(_3493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8824__S (.DIODE(_3926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8825__A1 (.DIODE(_3483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8825__S (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8827__A1 (.DIODE(_3499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8827__B1 (.DIODE(_3501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8827__C1 (.DIODE(_3926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8828__A1 (.DIODE(_3504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8829__A1 (.DIODE(_3497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8829__S (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8831__A2 (.DIODE(_3516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8832__A1 (.DIODE(_3511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8832__B1 (.DIODE(_3513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8834__A1 (.DIODE(_3507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8835__A1 (.DIODE(_0118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8835__A2 (.DIODE(_3927_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8835__B1 (.DIODE(_3917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8836__A1 (.DIODE(_3519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8836__A2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8836__B1 (.DIODE(_3520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8836__B2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8836__C1 (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8837__B1 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8837__B2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8838__A1 (.DIODE(_3526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8838__A2 (.DIODE(_3921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8838__B1 (.DIODE(_3528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8838__B2 (.DIODE(_3925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8838__C1 (.DIODE(_3960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8839__A2 (.DIODE(_3531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8840__A1 (.DIODE(_3523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8840__A2 (.DIODE(_3918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8842__B (.DIODE(_0855_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8845__C (.DIODE(_0199_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8853__A2 (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8853__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8854__A1 (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8857__B (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8858__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8863__A2 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8863__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8864__A2 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8866__B1 (.DIODE(_0483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8867__A1 (.DIODE(_0194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8867__B1 (.DIODE(_1757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8875__B (.DIODE(_0183_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8878__A2 (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8882__A1 (.DIODE(_4150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8882__A2 (.DIODE(_0470_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8882__A3 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8882__B1 (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8883__A1 (.DIODE(_0166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8890__A1 (.DIODE(_0205_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8890__A3 (.DIODE(_0184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8890__B1 (.DIODE(_0138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8891__A1 (.DIODE(_0166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8896__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__8896__A2 (.DIODE(_0480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8896__A3 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8896__B1 (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8897__A1 (.DIODE(_0166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8901__A1 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__8901__A2 (.DIODE(_0476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8901__A3 (.DIODE(_0206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8901__B1 (.DIODE(_0209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8902__A1 (.DIODE(_0166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8911__A1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8915__A1 (.DIODE(_0523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8917__A1 (.DIODE(_4118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8919__A (.DIODE(_0287_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8919__B (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__8924__B (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8932__B1 (.DIODE(net743));
 sky130_fd_sc_hd__diode_2 ANTENNA__8940__A1 (.DIODE(_0771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8942__B (.DIODE(net745));
 sky130_fd_sc_hd__diode_2 ANTENNA__8944__CLK (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8944__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8945__CLK (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8945__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8946__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8946__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8947__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8947__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8948__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8948__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8949__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8949__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8950__CLK (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8950__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8951__CLK (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8951__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8952__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8952__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8953__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8953__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8954__CLK (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8954__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8955__CLK (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8955__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8956__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8957__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8958__CLK (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8958__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8959__CLK (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8959__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8960__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8960__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8961__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8961__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8962__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8962__SET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8963__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8963__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8964__CLK (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8964__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8965__CLK (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8965__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8966__CLK (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8966__D (.DIODE(_0020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8966__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8967__CLK (.DIODE(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8967__D (.DIODE(_0021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8967__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__8968__CLK (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8968__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__8969__CLK (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8969__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8970__CLK (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8970__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8971__CLK (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8971__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8972__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8973__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8974__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8975__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8976__D (.DIODE(_0026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__8976__RESET_B (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__8977__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8977__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA__8978__CLK (.DIODE(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8978__RESET_B (.DIODE(net732));
 sky130_fd_sc_hd__diode_2 ANTENNA__8979__CLK (.DIODE(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA__8979__RESET_B (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f_clk_i_A (.DIODE(clknet_0_clk_i));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout732_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout733_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold10_A (.DIODE(\arbiter.crossbar[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold12_A (.DIODE(\arbiter.slave_sel[2][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold23_A (.DIODE(\arbiter.slave_sel[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold26_A (.DIODE(\arbiter.master_sel[0][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold41_A (.DIODE(\arbiter.master_sel[0][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold44_A (.DIODE(\arbiter.slave_sel[3][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_output366_A (.DIODE(net366));
 sky130_fd_sc_hd__diode_2 ANTENNA_output377_A (.DIODE(net377));
 sky130_fd_sc_hd__diode_2 ANTENNA_output388_A (.DIODE(net388));
 sky130_fd_sc_hd__diode_2 ANTENNA_output395_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_output398_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_output399_A (.DIODE(net399));
 sky130_fd_sc_hd__diode_2 ANTENNA_output404_A (.DIODE(net404));
 sky130_fd_sc_hd__diode_2 ANTENNA_output406_A (.DIODE(net406));
 sky130_fd_sc_hd__diode_2 ANTENNA_output407_A (.DIODE(net407));
 sky130_fd_sc_hd__diode_2 ANTENNA_output408_A (.DIODE(net408));
 sky130_fd_sc_hd__diode_2 ANTENNA_output409_A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_output410_A (.DIODE(net410));
 sky130_fd_sc_hd__diode_2 ANTENNA_output411_A (.DIODE(net411));
 sky130_fd_sc_hd__diode_2 ANTENNA_output412_A (.DIODE(net412));
 sky130_fd_sc_hd__diode_2 ANTENNA_output413_A (.DIODE(net413));
 sky130_fd_sc_hd__diode_2 ANTENNA_output414_A (.DIODE(net414));
 sky130_fd_sc_hd__diode_2 ANTENNA_output415_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_output416_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_output417_A (.DIODE(net417));
 sky130_fd_sc_hd__diode_2 ANTENNA_output418_A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_output419_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_output420_A (.DIODE(net420));
 sky130_fd_sc_hd__diode_2 ANTENNA_output421_A (.DIODE(net421));
 sky130_fd_sc_hd__diode_2 ANTENNA_output422_A (.DIODE(net422));
 sky130_fd_sc_hd__diode_2 ANTENNA_output423_A (.DIODE(net423));
 sky130_fd_sc_hd__diode_2 ANTENNA_output424_A (.DIODE(net424));
 sky130_fd_sc_hd__diode_2 ANTENNA_output425_A (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_output426_A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_output427_A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_output428_A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_output435_A (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_output440_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_output441_A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_output444_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_output445_A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_output446_A (.DIODE(net446));
 sky130_fd_sc_hd__diode_2 ANTENNA_output447_A (.DIODE(net447));
 sky130_fd_sc_hd__diode_2 ANTENNA_output449_A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_output450_A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_output452_A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_output454_A (.DIODE(net454));
 sky130_fd_sc_hd__diode_2 ANTENNA_output455_A (.DIODE(net455));
 sky130_fd_sc_hd__diode_2 ANTENNA_output456_A (.DIODE(net456));
 sky130_fd_sc_hd__diode_2 ANTENNA_output457_A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_output459_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_output468_A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_output479_A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_output490_A (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_output499_A (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_output500_A (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 ANTENNA_output501_A (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 ANTENNA_output503_A (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 ANTENNA_output506_A (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_output507_A (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA_output508_A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_output509_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 ANTENNA_output510_A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_output511_A (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 ANTENNA_output514_A (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 ANTENNA_output515_A (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA_output516_A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_output517_A (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 ANTENNA_output518_A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_output520_A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA_output586_A (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_output587_A (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA_output589_A (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA_output592_A (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA_output593_A (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA_output594_A (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_output595_A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_output602_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_output604_A (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_output606_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_output608_A (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA_output611_A (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA_output613_A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_output628_A (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA_output629_A (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_output639_A (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA_output683_A (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_output686_A (.DIODE(net686));
 sky130_fd_sc_hd__diode_2 ANTENNA_output688_A (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_output704_A (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_output705_A (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA_output706_A (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_output711_A (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_output719_A (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA_output721_A (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA_output722_A (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_output723_A (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA_output728_A (.DIODE(net728));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_672 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_423 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_266 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_423 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_182 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_802 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_268 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_203 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_131_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_131_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_339 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_132_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_255 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_133_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_171 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_402 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_135_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_135_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_135_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_136_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_254 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_591 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_137_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_620 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_138_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_139_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_139_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_140_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_140_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_141_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_142_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_142_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_259 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_143_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_143_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_143_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_144_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_144_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_555 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_145_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_145_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_145_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_272 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_146_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_147_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_147_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_148_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_242 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_149_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_149_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_546 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_336 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_150_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_151_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_151_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_151_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_152_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_153_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_153_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_153_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_504 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_154_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_155_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_155_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_155_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_23 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_594 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_852 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_812 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_310 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_588 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_932 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_904 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_682 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_866 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_923 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_626 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_927 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_592 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_791 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_535 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_650 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_826 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_42 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_812 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_930 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_934 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_829 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_786 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_933 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_878 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_874 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_856 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_934 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_135 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_458 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_759 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_350 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_627 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_79 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_312 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_394 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_836 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_536 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_918 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_742 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_688 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_700 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_320 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_792 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_938 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_199 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_936 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_903 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_931 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_311 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_315 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_367 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_897 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_905 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_926 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_280 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_734 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_907 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_919 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_644 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_868 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_872 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_928 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_936 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_599 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_763 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_739 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_328 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_651 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_392 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_827 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_196 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_448 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_869 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_262 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_822 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_422 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_674 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_479 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_812 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_375 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_651 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_784 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_636 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_583 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_451 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_310 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_945 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_652 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_460 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_598 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_703 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__buf_12 _4290_ (.A(\arbiter.slave_handled[2] ),
    .X(_4094_));
 sky130_fd_sc_hd__clkinv_4 _4291_ (.A(_4094_),
    .Y(_4095_));
 sky130_fd_sc_hd__nand2_1 _4292_ (.A(_4095_),
    .B(net231),
    .Y(_4096_));
 sky130_fd_sc_hd__inv_2 _4293_ (.A(_4096_),
    .Y(_4097_));
 sky130_fd_sc_hd__clkinv_4 _4294_ (.A(\arbiter.slave_handled[0] ),
    .Y(_4098_));
 sky130_fd_sc_hd__nand2_1 _4295_ (.A(_4098_),
    .B(net291),
    .Y(_4099_));
 sky130_fd_sc_hd__clkbuf_16 _4296_ (.A(\arbiter.slave_handled[1] ),
    .X(_4100_));
 sky130_fd_sc_hd__inv_2 _4297_ (.A(_4100_),
    .Y(_4101_));
 sky130_fd_sc_hd__nand2_1 _4298_ (.A(_4101_),
    .B(net328),
    .Y(_4102_));
 sky130_fd_sc_hd__nand2_1 _4299_ (.A(_4099_),
    .B(_4102_),
    .Y(_4103_));
 sky130_fd_sc_hd__nor2_1 _4300_ (.A(_4097_),
    .B(_4103_),
    .Y(_4104_));
 sky130_fd_sc_hd__buf_12 _4301_ (.A(\arbiter.slave_handled[3] ),
    .X(_4105_));
 sky130_fd_sc_hd__inv_6 _4302_ (.A(_4105_),
    .Y(_4106_));
 sky130_fd_sc_hd__buf_4 _4303_ (.A(net268),
    .X(_4107_));
 sky130_fd_sc_hd__inv_2 _4304_ (.A(net778),
    .Y(_4108_));
 sky130_fd_sc_hd__a21oi_1 _4305_ (.A1(_4106_),
    .A2(_4107_),
    .B1(_4108_),
    .Y(_4109_));
 sky130_fd_sc_hd__inv_2 _4306_ (.A(net737),
    .Y(_4110_));
 sky130_fd_sc_hd__a21o_1 _4307_ (.A1(_4104_),
    .A2(_4109_),
    .B1(_4110_),
    .X(_4111_));
 sky130_fd_sc_hd__nor2_4 _4308_ (.A(net772),
    .B(_4108_),
    .Y(_4112_));
 sky130_fd_sc_hd__buf_6 _4309_ (.A(\arbiter.slave_sel[0][0] ),
    .X(_4113_));
 sky130_fd_sc_hd__inv_6 _4310_ (.A(_4113_),
    .Y(_4114_));
 sky130_fd_sc_hd__nand2_1 _4311_ (.A(_4114_),
    .B(net361),
    .Y(_4115_));
 sky130_fd_sc_hd__nand2_1 _4312_ (.A(_4113_),
    .B(net363),
    .Y(_4116_));
 sky130_fd_sc_hd__nand2_1 _4313_ (.A(_4115_),
    .B(_4116_),
    .Y(_4117_));
 sky130_fd_sc_hd__buf_8 _4314_ (.A(net770),
    .X(_4118_));
 sky130_fd_sc_hd__inv_6 _4315_ (.A(_4118_),
    .Y(_4119_));
 sky130_fd_sc_hd__nand2_1 _4316_ (.A(_4117_),
    .B(_4119_),
    .Y(_4120_));
 sky130_fd_sc_hd__nand2_1 _4317_ (.A(_4114_),
    .B(net231),
    .Y(_4121_));
 sky130_fd_sc_hd__nand2_1 _4318_ (.A(_4113_),
    .B(net233),
    .Y(_4122_));
 sky130_fd_sc_hd__nand2_1 _4319_ (.A(_4121_),
    .B(_4122_),
    .Y(_4123_));
 sky130_fd_sc_hd__nand2_1 _4320_ (.A(_4123_),
    .B(_4118_),
    .Y(_4124_));
 sky130_fd_sc_hd__nand2_1 _4321_ (.A(_4120_),
    .B(_4124_),
    .Y(_4125_));
 sky130_fd_sc_hd__nand2_1 _4322_ (.A(_4125_),
    .B(_4114_),
    .Y(_4126_));
 sky130_fd_sc_hd__buf_8 _4323_ (.A(_4113_),
    .X(_4127_));
 sky130_fd_sc_hd__a21oi_1 _4324_ (.A1(_4127_),
    .A2(_4107_),
    .B1(_4119_),
    .Y(_4128_));
 sky130_fd_sc_hd__nand2_1 _4325_ (.A(_4126_),
    .B(_4128_),
    .Y(_4129_));
 sky130_fd_sc_hd__nand2_1 _4326_ (.A(_4114_),
    .B(net295),
    .Y(_4130_));
 sky130_fd_sc_hd__nand2_1 _4327_ (.A(_4113_),
    .B(net297),
    .Y(_4131_));
 sky130_fd_sc_hd__nand2_1 _4328_ (.A(_4130_),
    .B(_4131_),
    .Y(_4132_));
 sky130_fd_sc_hd__nand2_1 _4329_ (.A(_4132_),
    .B(_4118_),
    .Y(_4133_));
 sky130_fd_sc_hd__nand2_1 _4330_ (.A(_4114_),
    .B(net291),
    .Y(_4134_));
 sky130_fd_sc_hd__nand2_1 _4331_ (.A(_4113_),
    .B(net293),
    .Y(_4135_));
 sky130_fd_sc_hd__nand2_1 _4332_ (.A(_4134_),
    .B(_4135_),
    .Y(_4136_));
 sky130_fd_sc_hd__nand2_1 _4333_ (.A(_4136_),
    .B(_4119_),
    .Y(_4137_));
 sky130_fd_sc_hd__nand2_1 _4334_ (.A(_4133_),
    .B(_4137_),
    .Y(_4138_));
 sky130_fd_sc_hd__nand2_1 _4335_ (.A(_4138_),
    .B(_4114_),
    .Y(_4139_));
 sky130_fd_sc_hd__nand2_1 _4336_ (.A(_4114_),
    .B(net326),
    .Y(_4140_));
 sky130_fd_sc_hd__nand2_1 _4337_ (.A(_4113_),
    .B(net328),
    .Y(_4141_));
 sky130_fd_sc_hd__nand2_1 _4338_ (.A(_4140_),
    .B(_4141_),
    .Y(_4142_));
 sky130_fd_sc_hd__a21oi_1 _4339_ (.A1(_4142_),
    .A2(_4113_),
    .B1(_4118_),
    .Y(_4143_));
 sky130_fd_sc_hd__nand2_1 _4340_ (.A(_4139_),
    .B(_4143_),
    .Y(_4144_));
 sky130_fd_sc_hd__nand2_4 _4341_ (.A(_4129_),
    .B(_4144_),
    .Y(_4145_));
 sky130_fd_sc_hd__inv_4 _4342_ (.A(\arbiter.master_sel[0][0] ),
    .Y(_4146_));
 sky130_fd_sc_hd__nor2_4 _4343_ (.A(\arbiter.master_sel[0][1] ),
    .B(_4146_),
    .Y(_4147_));
 sky130_fd_sc_hd__nand2_1 _4344_ (.A(_4147_),
    .B(net11),
    .Y(_4148_));
 sky130_fd_sc_hd__nor2_4 _4345_ (.A(\arbiter.master_sel[0][0] ),
    .B(\arbiter.master_sel[0][1] ),
    .Y(_4149_));
 sky130_fd_sc_hd__buf_6 _4346_ (.A(net176),
    .X(_4150_));
 sky130_fd_sc_hd__nand2_1 _4347_ (.A(_4149_),
    .B(_4150_),
    .Y(_4151_));
 sky130_fd_sc_hd__and2_1 _4348_ (.A(_4148_),
    .B(_4151_),
    .X(_4152_));
 sky130_fd_sc_hd__buf_8 _4349_ (.A(_4146_),
    .X(_4153_));
 sky130_fd_sc_hd__nand2_1 _4350_ (.A(_4153_),
    .B(net74),
    .Y(_4154_));
 sky130_fd_sc_hd__nand2_1 _4351_ (.A(net138),
    .B(\arbiter.master_sel[0][0] ),
    .Y(_4155_));
 sky130_fd_sc_hd__inv_2 _4352_ (.A(\arbiter.master_sel[0][1] ),
    .Y(_4156_));
 sky130_fd_sc_hd__a21o_1 _4353_ (.A1(_4154_),
    .A2(_4155_),
    .B1(_4156_),
    .X(_4157_));
 sky130_fd_sc_hd__inv_2 _4354_ (.A(\arbiter.state[0][1] ),
    .Y(_4158_));
 sky130_fd_sc_hd__nor2_1 _4355_ (.A(net778),
    .B(_4158_),
    .Y(_4159_));
 sky130_fd_sc_hd__nand3_2 _4356_ (.A(_4152_),
    .B(_4157_),
    .C(_4159_),
    .Y(_4160_));
 sky130_fd_sc_hd__inv_4 _4357_ (.A(_4160_),
    .Y(_4161_));
 sky130_fd_sc_hd__nor2_2 _4358_ (.A(net778),
    .B(net772),
    .Y(_4162_));
 sky130_fd_sc_hd__inv_2 _4359_ (.A(_4162_),
    .Y(_4163_));
 sky130_fd_sc_hd__nor2_1 _4360_ (.A(_4110_),
    .B(_4163_),
    .Y(_4164_));
 sky130_fd_sc_hd__inv_2 _4361_ (.A(_4164_),
    .Y(_4165_));
 sky130_fd_sc_hd__inv_2 _4362_ (.A(net766),
    .Y(_4166_));
 sky130_fd_sc_hd__nand2_2 _4363_ (.A(_4166_),
    .B(_4150_),
    .Y(_4167_));
 sky130_fd_sc_hd__nand2_1 _4364_ (.A(_4167_),
    .B(_4108_),
    .Y(_4168_));
 sky130_fd_sc_hd__inv_2 _4365_ (.A(\arbiter.master_handled[1] ),
    .Y(_4169_));
 sky130_fd_sc_hd__nand2_1 _4366_ (.A(_4169_),
    .B(net11),
    .Y(_4170_));
 sky130_fd_sc_hd__inv_2 _4367_ (.A(net768),
    .Y(_4171_));
 sky130_fd_sc_hd__nand2_1 _4368_ (.A(_4171_),
    .B(net74),
    .Y(_4172_));
 sky130_fd_sc_hd__inv_2 _4369_ (.A(net767),
    .Y(_4173_));
 sky130_fd_sc_hd__nand2_1 _4370_ (.A(_4173_),
    .B(net138),
    .Y(_4174_));
 sky130_fd_sc_hd__nand3_1 _4371_ (.A(_4170_),
    .B(_4172_),
    .C(_4174_),
    .Y(_4175_));
 sky130_fd_sc_hd__nor2_1 _4372_ (.A(_4168_),
    .B(_4175_),
    .Y(_4176_));
 sky130_fd_sc_hd__nor2_1 _4373_ (.A(_4165_),
    .B(_4176_),
    .Y(_4177_));
 sky130_fd_sc_hd__a221o_1 _4374_ (.A1(_4111_),
    .A2(_4112_),
    .B1(_4145_),
    .B2(_4161_),
    .C1(_4177_),
    .X(_4178_));
 sky130_fd_sc_hd__buf_2 _4375_ (.A(_4178_),
    .X(_0020_));
 sky130_fd_sc_hd__nand2_1 _4376_ (.A(_4106_),
    .B(_4107_),
    .Y(_4179_));
 sky130_fd_sc_hd__and2_1 _4377_ (.A(_4179_),
    .B(_4158_),
    .X(_4180_));
 sky130_fd_sc_hd__nand2_1 _4378_ (.A(net773),
    .B(net737),
    .Y(_4181_));
 sky130_fd_sc_hd__a21oi_1 _4379_ (.A1(_4104_),
    .A2(_4180_),
    .B1(_4181_),
    .Y(_4182_));
 sky130_fd_sc_hd__or2_1 _4380_ (.A(net779),
    .B(_4182_),
    .X(_4183_));
 sky130_fd_sc_hd__buf_2 _4381_ (.A(_4183_),
    .X(_0021_));
 sky130_fd_sc_hd__inv_4 _4382_ (.A(\arbiter.state[1][1] ),
    .Y(_4184_));
 sky130_fd_sc_hd__nor2_2 _4383_ (.A(net765),
    .B(_4184_),
    .Y(_4185_));
 sky130_fd_sc_hd__nor2_8 _4384_ (.A(_4127_),
    .B(_4119_),
    .Y(_4186_));
 sky130_fd_sc_hd__nand3_1 _4385_ (.A(_4145_),
    .B(_4186_),
    .C(_4161_),
    .Y(_4187_));
 sky130_fd_sc_hd__nand2_1 _4386_ (.A(_4187_),
    .B(_4094_),
    .Y(_4188_));
 sky130_fd_sc_hd__o21ai_2 _4387_ (.A1(_4109_),
    .A2(_4180_),
    .B1(_4104_),
    .Y(_4189_));
 sky130_fd_sc_hd__nand3_1 _4388_ (.A(_4179_),
    .B(_4096_),
    .C(_4119_),
    .Y(_4190_));
 sky130_fd_sc_hd__inv_2 _4389_ (.A(_4103_),
    .Y(_4191_));
 sky130_fd_sc_hd__nand2_1 _4390_ (.A(_4190_),
    .B(_4191_),
    .Y(_4192_));
 sky130_fd_sc_hd__nor2_1 _4391_ (.A(_4110_),
    .B(_4192_),
    .Y(_4193_));
 sky130_fd_sc_hd__nand2_1 _4392_ (.A(_4179_),
    .B(_4114_),
    .Y(_4194_));
 sky130_fd_sc_hd__nand2_1 _4393_ (.A(_4194_),
    .B(_4096_),
    .Y(_4195_));
 sky130_fd_sc_hd__nand2_1 _4394_ (.A(_4195_),
    .B(_4102_),
    .Y(_4196_));
 sky130_fd_sc_hd__nand2_1 _4395_ (.A(_4196_),
    .B(_4099_),
    .Y(_4197_));
 sky130_fd_sc_hd__nand3_1 _4396_ (.A(_4189_),
    .B(_4193_),
    .C(_4197_),
    .Y(_4198_));
 sky130_fd_sc_hd__nand2_1 _4397_ (.A(_4198_),
    .B(_4095_),
    .Y(_4199_));
 sky130_fd_sc_hd__nand2_1 _4398_ (.A(_4199_),
    .B(_4112_),
    .Y(_4200_));
 sky130_fd_sc_hd__nand3_1 _4399_ (.A(_4188_),
    .B(net231),
    .C(_4200_),
    .Y(_4201_));
 sky130_fd_sc_hd__inv_2 _4400_ (.A(_4201_),
    .Y(_4202_));
 sky130_fd_sc_hd__nor2_1 _4401_ (.A(_4127_),
    .B(_4118_),
    .Y(_4203_));
 sky130_fd_sc_hd__buf_12 _4402_ (.A(_4203_),
    .X(_4204_));
 sky130_fd_sc_hd__nand3_1 _4403_ (.A(_4145_),
    .B(_4204_),
    .C(_4161_),
    .Y(_4205_));
 sky130_fd_sc_hd__nand2_1 _4404_ (.A(_4205_),
    .B(\arbiter.slave_handled[0] ),
    .Y(_4206_));
 sky130_fd_sc_hd__inv_2 _4405_ (.A(_4192_),
    .Y(_4207_));
 sky130_fd_sc_hd__nor2_1 _4406_ (.A(_4110_),
    .B(_4207_),
    .Y(_4208_));
 sky130_fd_sc_hd__nand3_1 _4407_ (.A(_4208_),
    .B(_4189_),
    .C(_4197_),
    .Y(_4209_));
 sky130_fd_sc_hd__nand2_1 _4408_ (.A(_4209_),
    .B(_4098_),
    .Y(_4210_));
 sky130_fd_sc_hd__nand2_1 _4409_ (.A(_4210_),
    .B(_4112_),
    .Y(_4211_));
 sky130_fd_sc_hd__nand3_1 _4410_ (.A(_4206_),
    .B(net291),
    .C(_4211_),
    .Y(_4212_));
 sky130_fd_sc_hd__nor2_4 _4411_ (.A(_4118_),
    .B(_4114_),
    .Y(_4213_));
 sky130_fd_sc_hd__nand3_1 _4412_ (.A(_4145_),
    .B(_4213_),
    .C(_4161_),
    .Y(_4214_));
 sky130_fd_sc_hd__nand2_1 _4413_ (.A(_4214_),
    .B(_4100_),
    .Y(_4215_));
 sky130_fd_sc_hd__a21boi_2 _4414_ (.A1(_4195_),
    .A2(_4102_),
    .B1_N(_4099_),
    .Y(_4216_));
 sky130_fd_sc_hd__nand3_1 _4415_ (.A(_4208_),
    .B(_4189_),
    .C(_4216_),
    .Y(_4217_));
 sky130_fd_sc_hd__nand2_1 _4416_ (.A(_4217_),
    .B(_4101_),
    .Y(_4218_));
 sky130_fd_sc_hd__nand2_1 _4417_ (.A(_4218_),
    .B(_4112_),
    .Y(_4219_));
 sky130_fd_sc_hd__nand3_1 _4418_ (.A(_4215_),
    .B(net328),
    .C(_4219_),
    .Y(_4220_));
 sky130_fd_sc_hd__nand2_1 _4419_ (.A(_4212_),
    .B(_4220_),
    .Y(_4221_));
 sky130_fd_sc_hd__nor2_1 _4420_ (.A(_4202_),
    .B(_4221_),
    .Y(_4222_));
 sky130_fd_sc_hd__nand2_8 _4421_ (.A(_4127_),
    .B(_4118_),
    .Y(_4223_));
 sky130_fd_sc_hd__nor2_1 _4422_ (.A(_4223_),
    .B(_4160_),
    .Y(_4224_));
 sky130_fd_sc_hd__nand2_1 _4423_ (.A(_4145_),
    .B(_4224_),
    .Y(_4225_));
 sky130_fd_sc_hd__nand2_1 _4424_ (.A(_4225_),
    .B(_4105_),
    .Y(_4226_));
 sky130_fd_sc_hd__nand3_1 _4425_ (.A(_4216_),
    .B(_4189_),
    .C(_4193_),
    .Y(_4227_));
 sky130_fd_sc_hd__nand2_1 _4426_ (.A(_4227_),
    .B(_4106_),
    .Y(_4228_));
 sky130_fd_sc_hd__nand2_1 _4427_ (.A(_4228_),
    .B(_4112_),
    .Y(_4229_));
 sky130_fd_sc_hd__nand3_2 _4428_ (.A(_4226_),
    .B(_4229_),
    .C(_4107_),
    .Y(_4230_));
 sky130_fd_sc_hd__nand2_1 _4429_ (.A(_4230_),
    .B(_4184_),
    .Y(_4231_));
 sky130_fd_sc_hd__inv_2 _4430_ (.A(_4231_),
    .Y(_4232_));
 sky130_fd_sc_hd__buf_12 _4431_ (.A(\arbiter.state[1][1] ),
    .X(_4233_));
 sky130_fd_sc_hd__inv_2 _4432_ (.A(net765),
    .Y(_4234_));
 sky130_fd_sc_hd__nor2_8 _4433_ (.A(_4233_),
    .B(_4234_),
    .Y(_4235_));
 sky130_fd_sc_hd__nand2_1 _4434_ (.A(_4235_),
    .B(net743),
    .Y(_4236_));
 sky130_fd_sc_hd__a21oi_1 _4435_ (.A1(_4222_),
    .A2(_4232_),
    .B1(_4236_),
    .Y(_4237_));
 sky130_fd_sc_hd__or2_1 _4436_ (.A(_4185_),
    .B(_4237_),
    .X(_4238_));
 sky130_fd_sc_hd__buf_1 _4437_ (.A(_4238_),
    .X(_0027_));
 sky130_fd_sc_hd__clkbuf_16 _4438_ (.A(\arbiter.state[2][1] ),
    .X(_4239_));
 sky130_fd_sc_hd__inv_2 _4439_ (.A(net762),
    .Y(_4240_));
 sky130_fd_sc_hd__nor2_4 _4440_ (.A(_4239_),
    .B(_4240_),
    .Y(_4241_));
 sky130_fd_sc_hd__nand2_2 _4441_ (.A(_4241_),
    .B(net734),
    .Y(_4242_));
 sky130_fd_sc_hd__inv_2 _4442_ (.A(net743),
    .Y(_4243_));
 sky130_fd_sc_hd__inv_2 _4443_ (.A(_4221_),
    .Y(_4244_));
 sky130_fd_sc_hd__clkinv_8 _4444_ (.A(net756),
    .Y(_4245_));
 sky130_fd_sc_hd__nand3_1 _4445_ (.A(_4201_),
    .B(_4245_),
    .C(_4230_),
    .Y(_4246_));
 sky130_fd_sc_hd__nand2_1 _4446_ (.A(_4244_),
    .B(_4246_),
    .Y(_4247_));
 sky130_fd_sc_hd__nor2_1 _4447_ (.A(_4243_),
    .B(_4247_),
    .Y(_4248_));
 sky130_fd_sc_hd__nand2_1 _4448_ (.A(_4230_),
    .B(net765),
    .Y(_4249_));
 sky130_fd_sc_hd__inv_2 _4449_ (.A(_4249_),
    .Y(_4250_));
 sky130_fd_sc_hd__o21ai_2 _4450_ (.A1(_4232_),
    .A2(_4250_),
    .B1(_4222_),
    .Y(_4251_));
 sky130_fd_sc_hd__buf_8 _4451_ (.A(\arbiter.slave_sel[1][0] ),
    .X(_4252_));
 sky130_fd_sc_hd__inv_6 _4452_ (.A(_4252_),
    .Y(_4253_));
 sky130_fd_sc_hd__nand2_1 _4453_ (.A(_4230_),
    .B(_4253_),
    .Y(_4254_));
 sky130_fd_sc_hd__nand2_1 _4454_ (.A(_4254_),
    .B(_4201_),
    .Y(_4255_));
 sky130_fd_sc_hd__nand2_1 _4455_ (.A(_4255_),
    .B(_4220_),
    .Y(_4256_));
 sky130_fd_sc_hd__nand2_1 _4456_ (.A(_4256_),
    .B(_4212_),
    .Y(_4257_));
 sky130_fd_sc_hd__nand3_1 _4457_ (.A(_4248_),
    .B(_4251_),
    .C(_4257_),
    .Y(_4258_));
 sky130_fd_sc_hd__nand2_1 _4458_ (.A(_4188_),
    .B(_4200_),
    .Y(_4259_));
 sky130_fd_sc_hd__inv_2 _4459_ (.A(_4259_),
    .Y(_4260_));
 sky130_fd_sc_hd__nand2_1 _4460_ (.A(_4258_),
    .B(_4260_),
    .Y(_4261_));
 sky130_fd_sc_hd__mux2_1 _4461_ (.A0(net361),
    .A1(net363),
    .S(_4252_),
    .X(_4262_));
 sky130_fd_sc_hd__nand2_8 _4462_ (.A(_4252_),
    .B(\arbiter.slave_sel[1][1] ),
    .Y(_4263_));
 sky130_fd_sc_hd__inv_2 _4463_ (.A(_4263_),
    .Y(_4264_));
 sky130_fd_sc_hd__nor2_8 _4464_ (.A(_4252_),
    .B(_4245_),
    .Y(_4265_));
 sky130_fd_sc_hd__a22o_1 _4465_ (.A1(_4264_),
    .A2(net233),
    .B1(net231),
    .B2(_4265_),
    .X(_4266_));
 sky130_fd_sc_hd__a21oi_1 _4466_ (.A1(_4245_),
    .A2(_4262_),
    .B1(_4266_),
    .Y(_4267_));
 sky130_fd_sc_hd__buf_8 _4467_ (.A(_4264_),
    .X(_4268_));
 sky130_fd_sc_hd__nand2_1 _4468_ (.A(_4268_),
    .B(_4107_),
    .Y(_4269_));
 sky130_fd_sc_hd__o211ai_2 _4469_ (.A1(_4252_),
    .A2(_4267_),
    .B1(\arbiter.slave_sel[1][1] ),
    .C1(_4269_),
    .Y(_4270_));
 sky130_fd_sc_hd__nand2_8 _4470_ (.A(_4245_),
    .B(_4252_),
    .Y(_4271_));
 sky130_fd_sc_hd__nand2_8 _4471_ (.A(_4253_),
    .B(_4245_),
    .Y(_4272_));
 sky130_fd_sc_hd__o22a_1 _4472_ (.A1(net293),
    .A2(_4271_),
    .B1(net291),
    .B2(_4272_),
    .X(_4273_));
 sky130_fd_sc_hd__inv_2 _4473_ (.A(net297),
    .Y(_4274_));
 sky130_fd_sc_hd__nand2_1 _4474_ (.A(_4274_),
    .B(_4252_),
    .Y(_4275_));
 sky130_fd_sc_hd__a21o_1 _4475_ (.A1(_4275_),
    .A2(net295),
    .B1(_4245_),
    .X(_4276_));
 sky130_fd_sc_hd__and3_1 _4476_ (.A(_4273_),
    .B(_4253_),
    .C(_4276_),
    .X(_4277_));
 sky130_fd_sc_hd__clkinv_16 _4477_ (.A(_4272_),
    .Y(_4278_));
 sky130_fd_sc_hd__nand2_1 _4478_ (.A(_4278_),
    .B(net326),
    .Y(_4279_));
 sky130_fd_sc_hd__inv_12 _4479_ (.A(_4271_),
    .Y(_4280_));
 sky130_fd_sc_hd__nand2_1 _4480_ (.A(_4280_),
    .B(net328),
    .Y(_4281_));
 sky130_fd_sc_hd__nand2_1 _4481_ (.A(_4265_),
    .B(net330),
    .Y(_4282_));
 sky130_fd_sc_hd__nand2_1 _4482_ (.A(_4264_),
    .B(net333),
    .Y(_4283_));
 sky130_fd_sc_hd__a41o_1 _4483_ (.A1(_4279_),
    .A2(_4281_),
    .A3(_4282_),
    .A4(_4283_),
    .B1(_4253_),
    .X(_4284_));
 sky130_fd_sc_hd__nand3b_1 _4484_ (.A_N(_4277_),
    .B(_4284_),
    .C(_4245_),
    .Y(_4285_));
 sky130_fd_sc_hd__nand2_4 _4485_ (.A(_4270_),
    .B(_4285_),
    .Y(_4286_));
 sky130_fd_sc_hd__inv_6 _4486_ (.A(_4265_),
    .Y(_4287_));
 sky130_fd_sc_hd__clkinv_4 _4487_ (.A(\arbiter.master_sel[1][0] ),
    .Y(_4288_));
 sky130_fd_sc_hd__nand2_8 _4488_ (.A(_4288_),
    .B(\arbiter.master_sel[1][1] ),
    .Y(_4289_));
 sky130_fd_sc_hd__nand2_8 _4489_ (.A(\arbiter.master_sel[1][0] ),
    .B(\arbiter.master_sel[1][1] ),
    .Y(_0036_));
 sky130_fd_sc_hd__clkinv_4 _4490_ (.A(net748),
    .Y(_0037_));
 sky130_fd_sc_hd__nand2_8 _4491_ (.A(_0037_),
    .B(\arbiter.master_sel[1][0] ),
    .Y(_0038_));
 sky130_fd_sc_hd__nand2_8 _4492_ (.A(_4288_),
    .B(_0037_),
    .Y(_0039_));
 sky130_fd_sc_hd__o22a_1 _4493_ (.A1(net11),
    .A2(_0038_),
    .B1(_4150_),
    .B2(_0039_),
    .X(_0040_));
 sky130_fd_sc_hd__o221a_4 _4494_ (.A1(net74),
    .A2(_4289_),
    .B1(net138),
    .B2(_0036_),
    .C1(_0040_),
    .X(_0041_));
 sky130_fd_sc_hd__nor2_1 _4495_ (.A(_4287_),
    .B(_0041_),
    .Y(_0042_));
 sky130_fd_sc_hd__a31o_1 _4496_ (.A1(_4286_),
    .A2(_4185_),
    .A3(_0042_),
    .B1(_4260_),
    .X(_0043_));
 sky130_fd_sc_hd__inv_2 _4497_ (.A(_4235_),
    .Y(_0044_));
 sky130_fd_sc_hd__nand2_1 _4498_ (.A(_0043_),
    .B(_0044_),
    .Y(_0045_));
 sky130_fd_sc_hd__nand2_1 _4499_ (.A(_4261_),
    .B(_0045_),
    .Y(_0046_));
 sky130_fd_sc_hd__nand2_1 _4500_ (.A(_0046_),
    .B(net231),
    .Y(_0047_));
 sky130_fd_sc_hd__inv_2 _4501_ (.A(_0047_),
    .Y(_0048_));
 sky130_fd_sc_hd__and2_1 _4502_ (.A(_4247_),
    .B(\arbiter.crossbar[2] ),
    .X(_0049_));
 sky130_fd_sc_hd__nand3_1 _4503_ (.A(_0049_),
    .B(_4257_),
    .C(_4251_),
    .Y(_0050_));
 sky130_fd_sc_hd__nand2_1 _4504_ (.A(_4206_),
    .B(_4211_),
    .Y(_0051_));
 sky130_fd_sc_hd__inv_2 _4505_ (.A(_0051_),
    .Y(_0052_));
 sky130_fd_sc_hd__nand2_1 _4506_ (.A(_0050_),
    .B(_0052_),
    .Y(_0053_));
 sky130_fd_sc_hd__nor2_1 _4507_ (.A(_4272_),
    .B(_0041_),
    .Y(_0054_));
 sky130_fd_sc_hd__a31o_1 _4508_ (.A1(_4286_),
    .A2(_4185_),
    .A3(_0054_),
    .B1(_0052_),
    .X(_0055_));
 sky130_fd_sc_hd__buf_8 _4509_ (.A(_0044_),
    .X(_0056_));
 sky130_fd_sc_hd__nand2_1 _4510_ (.A(_0055_),
    .B(_0056_),
    .Y(_0057_));
 sky130_fd_sc_hd__nand2_1 _4511_ (.A(_0053_),
    .B(_0057_),
    .Y(_0058_));
 sky130_fd_sc_hd__nand2_1 _4512_ (.A(_0058_),
    .B(net291),
    .Y(_0059_));
 sky130_fd_sc_hd__a21boi_1 _4513_ (.A1(_4255_),
    .A2(_4220_),
    .B1_N(_4212_),
    .Y(_0060_));
 sky130_fd_sc_hd__nand3_1 _4514_ (.A(_0049_),
    .B(_0060_),
    .C(_4251_),
    .Y(_0061_));
 sky130_fd_sc_hd__nand2_1 _4515_ (.A(_4215_),
    .B(_4219_),
    .Y(_0062_));
 sky130_fd_sc_hd__inv_2 _4516_ (.A(_0062_),
    .Y(_0063_));
 sky130_fd_sc_hd__nand2_1 _4517_ (.A(_0061_),
    .B(_0063_),
    .Y(_0064_));
 sky130_fd_sc_hd__nor2_1 _4518_ (.A(_4271_),
    .B(_0041_),
    .Y(_0065_));
 sky130_fd_sc_hd__a31o_1 _4519_ (.A1(_4286_),
    .A2(_4185_),
    .A3(_0065_),
    .B1(_0063_),
    .X(_0066_));
 sky130_fd_sc_hd__nand2_1 _4520_ (.A(_0066_),
    .B(_0056_),
    .Y(_0067_));
 sky130_fd_sc_hd__nand2_2 _4521_ (.A(_0064_),
    .B(_0067_),
    .Y(_0068_));
 sky130_fd_sc_hd__nand2_1 _4522_ (.A(_0068_),
    .B(net328),
    .Y(_0069_));
 sky130_fd_sc_hd__nand2_1 _4523_ (.A(_0059_),
    .B(_0069_),
    .Y(_0070_));
 sky130_fd_sc_hd__nor2_1 _4524_ (.A(_0048_),
    .B(_0070_),
    .Y(_0071_));
 sky130_fd_sc_hd__nand3_1 _4525_ (.A(_4248_),
    .B(_0060_),
    .C(_4251_),
    .Y(_0072_));
 sky130_fd_sc_hd__nand2_1 _4526_ (.A(_4226_),
    .B(_4229_),
    .Y(_0073_));
 sky130_fd_sc_hd__inv_2 _4527_ (.A(_0073_),
    .Y(_0074_));
 sky130_fd_sc_hd__nand2_1 _4528_ (.A(_0072_),
    .B(_0074_),
    .Y(_0075_));
 sky130_fd_sc_hd__nor2_1 _4529_ (.A(_4263_),
    .B(_0041_),
    .Y(_0076_));
 sky130_fd_sc_hd__a31o_1 _4530_ (.A1(_4286_),
    .A2(_4185_),
    .A3(_0076_),
    .B1(_0074_),
    .X(_0077_));
 sky130_fd_sc_hd__nand2_1 _4531_ (.A(_0077_),
    .B(_0056_),
    .Y(_0078_));
 sky130_fd_sc_hd__nand2_2 _4532_ (.A(_0075_),
    .B(_0078_),
    .Y(_0079_));
 sky130_fd_sc_hd__a21oi_1 _4533_ (.A1(_0079_),
    .A2(_4107_),
    .B1(_4239_),
    .Y(_0080_));
 sky130_fd_sc_hd__nand2_1 _4534_ (.A(_0071_),
    .B(_0080_),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _4535_ (.A(_0081_),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_6 _4536_ (.A(_4239_),
    .Y(_0083_));
 sky130_fd_sc_hd__nor2_1 _4537_ (.A(net762),
    .B(_0083_),
    .Y(_0084_));
 sky130_fd_sc_hd__inv_2 _4538_ (.A(_0084_),
    .Y(_0085_));
 sky130_fd_sc_hd__o21a_1 _4539_ (.A1(_4242_),
    .A2(_0082_),
    .B1(_0085_),
    .X(_0086_));
 sky130_fd_sc_hd__inv_2 _4540_ (.A(_0086_),
    .Y(_0025_));
 sky130_fd_sc_hd__nand2_1 _4541_ (.A(_0079_),
    .B(_4107_),
    .Y(_0087_));
 sky130_fd_sc_hd__buf_8 _4542_ (.A(\arbiter.slave_sel[2][0] ),
    .X(_0088_));
 sky130_fd_sc_hd__inv_2 _4543_ (.A(_0088_),
    .Y(_0089_));
 sky130_fd_sc_hd__buf_8 _4544_ (.A(_0089_),
    .X(_0090_));
 sky130_fd_sc_hd__nand2_1 _4545_ (.A(_0087_),
    .B(_0090_),
    .Y(_0091_));
 sky130_fd_sc_hd__nand2_1 _4546_ (.A(_0091_),
    .B(_0047_),
    .Y(_0092_));
 sky130_fd_sc_hd__a21boi_1 _4547_ (.A1(_0092_),
    .A2(_0069_),
    .B1_N(_0059_),
    .Y(_0093_));
 sky130_fd_sc_hd__inv_2 _4548_ (.A(net734),
    .Y(_0094_));
 sky130_fd_sc_hd__inv_2 _4549_ (.A(_0070_),
    .Y(_0095_));
 sky130_fd_sc_hd__inv_6 _4550_ (.A(net745),
    .Y(_0096_));
 sky130_fd_sc_hd__nand3_1 _4551_ (.A(_0087_),
    .B(_0047_),
    .C(_0096_),
    .Y(_0097_));
 sky130_fd_sc_hd__nand2_1 _4552_ (.A(_0095_),
    .B(_0097_),
    .Y(_0098_));
 sky130_fd_sc_hd__nor2_1 _4553_ (.A(_0094_),
    .B(_0098_),
    .Y(_0099_));
 sky130_fd_sc_hd__and2_1 _4554_ (.A(_0087_),
    .B(net762),
    .X(_0100_));
 sky130_fd_sc_hd__o21ai_2 _4555_ (.A1(_0080_),
    .A2(_0100_),
    .B1(_0071_),
    .Y(_0101_));
 sky130_fd_sc_hd__nand3_1 _4556_ (.A(_0093_),
    .B(_0099_),
    .C(_0101_),
    .Y(_0102_));
 sky130_fd_sc_hd__nand2_1 _4557_ (.A(_0102_),
    .B(_0079_),
    .Y(_0103_));
 sky130_fd_sc_hd__inv_2 _4558_ (.A(net291),
    .Y(_0104_));
 sky130_fd_sc_hd__nor2_2 _4559_ (.A(_0088_),
    .B(\arbiter.slave_sel[2][1] ),
    .Y(_0105_));
 sky130_fd_sc_hd__inv_2 _4560_ (.A(_4107_),
    .Y(_0106_));
 sky130_fd_sc_hd__nand2_8 _4561_ (.A(_0088_),
    .B(\arbiter.slave_sel[2][1] ),
    .Y(_0107_));
 sky130_fd_sc_hd__inv_8 _4562_ (.A(_0107_),
    .Y(_0108_));
 sky130_fd_sc_hd__nor2_2 _4563_ (.A(\arbiter.slave_sel[2][1] ),
    .B(_0089_),
    .Y(_0109_));
 sky130_fd_sc_hd__inv_2 _4564_ (.A(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__nor2_8 _4565_ (.A(_0088_),
    .B(_0096_),
    .Y(_0111_));
 sky130_fd_sc_hd__inv_2 _4566_ (.A(net333),
    .Y(_0112_));
 sky130_fd_sc_hd__nor2_1 _4567_ (.A(_0112_),
    .B(_0107_),
    .Y(_0113_));
 sky130_fd_sc_hd__a22o_1 _4568_ (.A1(_0105_),
    .A2(net326),
    .B1(_0109_),
    .B2(net328),
    .X(_0114_));
 sky130_fd_sc_hd__a211o_1 _4569_ (.A1(net330),
    .A2(_0111_),
    .B1(_0113_),
    .C1(_0114_),
    .X(_0115_));
 sky130_fd_sc_hd__or3_1 _4570_ (.A(net231),
    .B(_0088_),
    .C(_0096_),
    .X(_0116_));
 sky130_fd_sc_hd__o21ai_1 _4571_ (.A1(_0110_),
    .A2(_0115_),
    .B1(_0116_),
    .Y(_0117_));
 sky130_fd_sc_hd__a221o_4 _4572_ (.A1(_0104_),
    .A2(_0105_),
    .B1(_0106_),
    .B2(_0108_),
    .C1(_0117_),
    .X(_0118_));
 sky130_fd_sc_hd__buf_4 _4573_ (.A(net776),
    .X(_0119_));
 sky130_fd_sc_hd__inv_2 _4574_ (.A(net754),
    .Y(_0120_));
 sky130_fd_sc_hd__nor2_4 _4575_ (.A(_0119_),
    .B(_0120_),
    .Y(_0121_));
 sky130_fd_sc_hd__clkinv_8 _4576_ (.A(_0121_),
    .Y(_0122_));
 sky130_fd_sc_hd__nand2_8 _4577_ (.A(_0119_),
    .B(\arbiter.master_sel[2][1] ),
    .Y(_0123_));
 sky130_fd_sc_hd__inv_2 _4578_ (.A(net11),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _4579_ (.A(_0119_),
    .Y(_0125_));
 sky130_fd_sc_hd__nor2_8 _4580_ (.A(\arbiter.master_sel[2][1] ),
    .B(_0125_),
    .Y(_0126_));
 sky130_fd_sc_hd__nor2_1 _4581_ (.A(_0119_),
    .B(\arbiter.master_sel[2][1] ),
    .Y(_0127_));
 sky130_fd_sc_hd__clkinv_4 _4582_ (.A(_0127_),
    .Y(_0128_));
 sky130_fd_sc_hd__nor2_1 _4583_ (.A(_4150_),
    .B(_0128_),
    .Y(_0129_));
 sky130_fd_sc_hd__a21oi_1 _4584_ (.A1(_0124_),
    .A2(_0126_),
    .B1(_0129_),
    .Y(_0130_));
 sky130_fd_sc_hd__o221a_4 _4585_ (.A1(net74),
    .A2(_0122_),
    .B1(net138),
    .B2(_0123_),
    .C1(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__nor2_1 _4586_ (.A(_0085_),
    .B(_0131_),
    .Y(_0132_));
 sky130_fd_sc_hd__a31o_1 _4587_ (.A1(_0118_),
    .A2(_0108_),
    .A3(_0132_),
    .B1(_0079_),
    .X(_0133_));
 sky130_fd_sc_hd__inv_4 _4588_ (.A(_4241_),
    .Y(_0134_));
 sky130_fd_sc_hd__nand2_1 _4589_ (.A(_0133_),
    .B(_0134_),
    .Y(_0135_));
 sky130_fd_sc_hd__nand2_1 _4590_ (.A(_0103_),
    .B(_0135_),
    .Y(_0136_));
 sky130_fd_sc_hd__nand2_1 _4591_ (.A(_0136_),
    .B(_4107_),
    .Y(_0137_));
 sky130_fd_sc_hd__inv_12 _4592_ (.A(net753),
    .Y(_0138_));
 sky130_fd_sc_hd__nand2_1 _4593_ (.A(_0137_),
    .B(_0138_),
    .Y(_0139_));
 sky130_fd_sc_hd__a21oi_1 _4594_ (.A1(_0095_),
    .A2(_0097_),
    .B1(_0094_),
    .Y(_0140_));
 sky130_fd_sc_hd__nand3_1 _4595_ (.A(_0140_),
    .B(_0093_),
    .C(_0101_),
    .Y(_0141_));
 sky130_fd_sc_hd__nand2_1 _4596_ (.A(_0141_),
    .B(_0068_),
    .Y(_0142_));
 sky130_fd_sc_hd__buf_12 _4597_ (.A(_0109_),
    .X(_0143_));
 sky130_fd_sc_hd__a31o_1 _4598_ (.A1(_0118_),
    .A2(_0143_),
    .A3(_0132_),
    .B1(_0068_),
    .X(_0144_));
 sky130_fd_sc_hd__nand2_1 _4599_ (.A(_0144_),
    .B(_0134_),
    .Y(_0145_));
 sky130_fd_sc_hd__nand2_1 _4600_ (.A(_0142_),
    .B(_0145_),
    .Y(_0146_));
 sky130_fd_sc_hd__nand2_1 _4601_ (.A(_0146_),
    .B(net328),
    .Y(_0147_));
 sky130_fd_sc_hd__nand2_1 _4602_ (.A(_0092_),
    .B(_0069_),
    .Y(_0148_));
 sky130_fd_sc_hd__nand2_1 _4603_ (.A(_0148_),
    .B(_0059_),
    .Y(_0149_));
 sky130_fd_sc_hd__nand3_1 _4604_ (.A(_0140_),
    .B(_0101_),
    .C(_0149_),
    .Y(_0150_));
 sky130_fd_sc_hd__nand2_1 _4605_ (.A(_0150_),
    .B(_0058_),
    .Y(_0151_));
 sky130_fd_sc_hd__inv_4 _4606_ (.A(_0105_),
    .Y(_0152_));
 sky130_fd_sc_hd__nand2_1 _4607_ (.A(_0118_),
    .B(_0132_),
    .Y(_0153_));
 sky130_fd_sc_hd__or2_1 _4608_ (.A(_0152_),
    .B(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__a31o_1 _4609_ (.A1(_0154_),
    .A2(_0057_),
    .A3(_0053_),
    .B1(_4241_),
    .X(_0155_));
 sky130_fd_sc_hd__nand2_1 _4610_ (.A(_0151_),
    .B(_0155_),
    .Y(_0156_));
 sky130_fd_sc_hd__nand2_1 _4611_ (.A(_0156_),
    .B(net291),
    .Y(_0157_));
 sky130_fd_sc_hd__nand3_1 _4612_ (.A(_0099_),
    .B(_0101_),
    .C(_0149_),
    .Y(_0158_));
 sky130_fd_sc_hd__nand2_1 _4613_ (.A(_0158_),
    .B(_0046_),
    .Y(_0159_));
 sky130_fd_sc_hd__clkinv_4 _4614_ (.A(_0111_),
    .Y(_0160_));
 sky130_fd_sc_hd__or2_1 _4615_ (.A(_0160_),
    .B(_0153_),
    .X(_0161_));
 sky130_fd_sc_hd__a31o_1 _4616_ (.A1(_0161_),
    .A2(_0045_),
    .A3(_4261_),
    .B1(_4241_),
    .X(_0162_));
 sky130_fd_sc_hd__nand2_1 _4617_ (.A(_0159_),
    .B(_0162_),
    .Y(_0163_));
 sky130_fd_sc_hd__nand2_1 _4618_ (.A(_0163_),
    .B(net231),
    .Y(_0164_));
 sky130_fd_sc_hd__nand3_1 _4619_ (.A(_0147_),
    .B(_0157_),
    .C(_0164_),
    .Y(_0165_));
 sky130_fd_sc_hd__clkinv_4 _4620_ (.A(net751),
    .Y(_0166_));
 sky130_fd_sc_hd__nor2_2 _4621_ (.A(net753),
    .B(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__buf_8 _4622_ (.A(_0167_),
    .X(_0168_));
 sky130_fd_sc_hd__nand2_1 _4623_ (.A(_0168_),
    .B(net740),
    .Y(_0169_));
 sky130_fd_sc_hd__o21bai_1 _4624_ (.A1(_0139_),
    .A2(_0165_),
    .B1_N(_0169_),
    .Y(_0170_));
 sky130_fd_sc_hd__nor2_1 _4625_ (.A(net751),
    .B(_0138_),
    .Y(_0171_));
 sky130_fd_sc_hd__inv_2 _4626_ (.A(_0171_),
    .Y(_0172_));
 sky130_fd_sc_hd__nand2_1 _4627_ (.A(_0170_),
    .B(_0172_),
    .Y(_0023_));
 sky130_fd_sc_hd__nand2_1 _4628_ (.A(_0023_),
    .B(net740),
    .Y(_0173_));
 sky130_fd_sc_hd__inv_2 _4629_ (.A(net740),
    .Y(_0174_));
 sky130_fd_sc_hd__and3_1 _4630_ (.A(_4243_),
    .B(_0094_),
    .C(_0174_),
    .X(_0175_));
 sky130_fd_sc_hd__inv_2 _4631_ (.A(_0175_),
    .Y(_0176_));
 sky130_fd_sc_hd__o2bb2a_1 _4632_ (.A1_N(\arbiter.crossbar[2] ),
    .A2_N(_0027_),
    .B1(_0094_),
    .B2(_0086_),
    .X(_0177_));
 sky130_fd_sc_hd__nand3_1 _4633_ (.A(_0173_),
    .B(_0176_),
    .C(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__or2_1 _4634_ (.A(_0176_),
    .B(_0021_),
    .X(_0179_));
 sky130_fd_sc_hd__nand2_2 _4635_ (.A(_0178_),
    .B(_0179_),
    .Y(_0180_));
 sky130_fd_sc_hd__nor2_1 _4636_ (.A(\arbiter.master_sel[3][0] ),
    .B(\arbiter.master_sel[3][1] ),
    .Y(_0181_));
 sky130_fd_sc_hd__clkinv_4 _4637_ (.A(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__clkinv_8 _4638_ (.A(\arbiter.master_sel[3][0] ),
    .Y(_0183_));
 sky130_fd_sc_hd__nor2_8 _4639_ (.A(\arbiter.master_sel[3][1] ),
    .B(_0183_),
    .Y(_0184_));
 sky130_fd_sc_hd__inv_8 _4640_ (.A(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__nand2_8 _4641_ (.A(\arbiter.master_sel[3][0] ),
    .B(\arbiter.master_sel[3][1] ),
    .Y(_0186_));
 sky130_fd_sc_hd__inv_2 _4642_ (.A(\arbiter.master_sel[3][1] ),
    .Y(_0187_));
 sky130_fd_sc_hd__nor2_1 _4643_ (.A(\arbiter.master_sel[3][0] ),
    .B(_0187_),
    .Y(_0188_));
 sky130_fd_sc_hd__inv_2 _4644_ (.A(_0188_),
    .Y(_0189_));
 sky130_fd_sc_hd__o22a_1 _4645_ (.A1(net138),
    .A2(_0186_),
    .B1(net74),
    .B2(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__o221a_4 _4646_ (.A1(_4150_),
    .A2(_0182_),
    .B1(net11),
    .B2(_0185_),
    .C1(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__nor2_8 _4647_ (.A(\arbiter.slave_sel[3][0] ),
    .B(\arbiter.slave_sel[3][1] ),
    .Y(_0192_));
 sky130_fd_sc_hd__nand2_8 _4648_ (.A(\arbiter.slave_sel[3][0] ),
    .B(\arbiter.slave_sel[3][1] ),
    .Y(_0193_));
 sky130_fd_sc_hd__inv_8 _4649_ (.A(_0193_),
    .Y(_0194_));
 sky130_fd_sc_hd__inv_2 _4650_ (.A(\arbiter.slave_sel[3][0] ),
    .Y(_0195_));
 sky130_fd_sc_hd__nor2_8 _4651_ (.A(\arbiter.slave_sel[3][1] ),
    .B(_0195_),
    .Y(_0196_));
 sky130_fd_sc_hd__inv_4 _4652_ (.A(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__buf_8 _4653_ (.A(\arbiter.slave_sel[3][0] ),
    .X(_0198_));
 sky130_fd_sc_hd__clkinv_4 _4654_ (.A(\arbiter.slave_sel[3][1] ),
    .Y(_0199_));
 sky130_fd_sc_hd__nor2_4 _4655_ (.A(_0198_),
    .B(_0199_),
    .Y(_0200_));
 sky130_fd_sc_hd__a22o_1 _4656_ (.A1(_0192_),
    .A2(net326),
    .B1(_0196_),
    .B2(net328),
    .X(_0201_));
 sky130_fd_sc_hd__a221o_1 _4657_ (.A1(net330),
    .A2(_0200_),
    .B1(net333),
    .B2(_0194_),
    .C1(_0201_),
    .X(_0202_));
 sky130_fd_sc_hd__or3_1 _4658_ (.A(net231),
    .B(_0198_),
    .C(_0199_),
    .X(_0203_));
 sky130_fd_sc_hd__o21ai_1 _4659_ (.A1(_0197_),
    .A2(_0202_),
    .B1(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__a221o_4 _4660_ (.A1(_0104_),
    .A2(_0192_),
    .B1(_0106_),
    .B2(_0194_),
    .C1(_0204_),
    .X(_0205_));
 sky130_fd_sc_hd__clkinv_4 _4661_ (.A(_0205_),
    .Y(_0206_));
 sky130_fd_sc_hd__or3_1 _4662_ (.A(_0172_),
    .B(_0191_),
    .C(_0206_),
    .X(_0207_));
 sky130_fd_sc_hd__inv_2 _4663_ (.A(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__clkbuf_16 _4664_ (.A(net753),
    .X(_0209_));
 sky130_fd_sc_hd__nor2_1 _4665_ (.A(net751),
    .B(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__nand2_1 _4666_ (.A(_0210_),
    .B(net740),
    .Y(_0211_));
 sky130_fd_sc_hd__nand2_1 _4667_ (.A(_4167_),
    .B(\arbiter.state[0][1] ),
    .Y(_0212_));
 sky130_fd_sc_hd__nor2_1 _4668_ (.A(_0212_),
    .B(_4175_),
    .Y(_0213_));
 sky130_fd_sc_hd__o21bai_1 _4669_ (.A1(_4168_),
    .A2(_4175_),
    .B1_N(_4110_),
    .Y(_0214_));
 sky130_fd_sc_hd__nor2_1 _4670_ (.A(_0213_),
    .B(_0214_),
    .Y(_0215_));
 sky130_fd_sc_hd__nand2_1 _4671_ (.A(_4174_),
    .B(_4153_),
    .Y(_0216_));
 sky130_fd_sc_hd__nand2_1 _4672_ (.A(_0216_),
    .B(_4172_),
    .Y(_0217_));
 sky130_fd_sc_hd__nand2_1 _4673_ (.A(_0217_),
    .B(_4170_),
    .Y(_0218_));
 sky130_fd_sc_hd__nand3_1 _4674_ (.A(_4172_),
    .B(_4174_),
    .C(_4156_),
    .Y(_0219_));
 sky130_fd_sc_hd__nand2_1 _4675_ (.A(_4170_),
    .B(_4167_),
    .Y(_0220_));
 sky130_fd_sc_hd__inv_2 _4676_ (.A(_0220_),
    .Y(_0221_));
 sky130_fd_sc_hd__nand2_1 _4677_ (.A(_0219_),
    .B(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__inv_2 _4678_ (.A(_0222_),
    .Y(_0223_));
 sky130_fd_sc_hd__a21oi_1 _4679_ (.A1(_0218_),
    .A2(_4167_),
    .B1(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__nand2_1 _4680_ (.A(_0215_),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__nand2_1 _4681_ (.A(_0225_),
    .B(_4166_),
    .Y(_0226_));
 sky130_fd_sc_hd__nand2_1 _4682_ (.A(_0226_),
    .B(_4162_),
    .Y(_0227_));
 sky130_fd_sc_hd__nand2_1 _4683_ (.A(_4149_),
    .B(_4108_),
    .Y(_0228_));
 sky130_fd_sc_hd__nand2_4 _4684_ (.A(_4152_),
    .B(_4157_),
    .Y(_0229_));
 sky130_fd_sc_hd__nor2_1 _4685_ (.A(_0228_),
    .B(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__nand2_1 _4686_ (.A(_4145_),
    .B(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__nand2_1 _4687_ (.A(_0231_),
    .B(net766),
    .Y(_0232_));
 sky130_fd_sc_hd__nand3_2 _4688_ (.A(_0227_),
    .B(_4150_),
    .C(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__nand2_1 _4689_ (.A(_0233_),
    .B(_4234_),
    .Y(_0234_));
 sky130_fd_sc_hd__inv_2 _4690_ (.A(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__nand2_1 _4691_ (.A(_0233_),
    .B(_4233_),
    .Y(_0236_));
 sky130_fd_sc_hd__inv_2 _4692_ (.A(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__nand2_1 _4693_ (.A(_0218_),
    .B(_4167_),
    .Y(_0238_));
 sky130_fd_sc_hd__nor2_1 _4694_ (.A(_0223_),
    .B(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__nand2_1 _4695_ (.A(_0215_),
    .B(_0239_),
    .Y(_0240_));
 sky130_fd_sc_hd__nand2_1 _4696_ (.A(_0240_),
    .B(_4169_),
    .Y(_0241_));
 sky130_fd_sc_hd__nand2_1 _4697_ (.A(_0241_),
    .B(_4162_),
    .Y(_0242_));
 sky130_fd_sc_hd__nand2_1 _4698_ (.A(_4147_),
    .B(_4108_),
    .Y(_0243_));
 sky130_fd_sc_hd__nor2_1 _4699_ (.A(_0243_),
    .B(_0229_),
    .Y(_0244_));
 sky130_fd_sc_hd__nand2_1 _4700_ (.A(_4145_),
    .B(_0244_),
    .Y(_0245_));
 sky130_fd_sc_hd__nand2_1 _4701_ (.A(_0245_),
    .B(\arbiter.master_handled[1] ),
    .Y(_0246_));
 sky130_fd_sc_hd__nand3_2 _4702_ (.A(_0242_),
    .B(net11),
    .C(_0246_),
    .Y(_0247_));
 sky130_fd_sc_hd__inv_2 _4703_ (.A(_0247_),
    .Y(_0248_));
 sky130_fd_sc_hd__a21oi_1 _4704_ (.A1(_0218_),
    .A2(_4167_),
    .B1(_0222_),
    .Y(_0249_));
 sky130_fd_sc_hd__nand2_1 _4705_ (.A(_0215_),
    .B(_0249_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand2_1 _4706_ (.A(_0250_),
    .B(_4171_),
    .Y(_0251_));
 sky130_fd_sc_hd__nand2_1 _4707_ (.A(_0251_),
    .B(_4162_),
    .Y(_0252_));
 sky130_fd_sc_hd__nand2_4 _4708_ (.A(_4153_),
    .B(\arbiter.master_sel[0][1] ),
    .Y(_0253_));
 sky130_fd_sc_hd__nor3_1 _4709_ (.A(\arbiter.state[0][0] ),
    .B(_0253_),
    .C(_0229_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand2_1 _4710_ (.A(_0254_),
    .B(_4145_),
    .Y(_0255_));
 sky130_fd_sc_hd__nand2_1 _4711_ (.A(_0255_),
    .B(net768),
    .Y(_0256_));
 sky130_fd_sc_hd__nand3_1 _4712_ (.A(_0252_),
    .B(_0256_),
    .C(net74),
    .Y(_0257_));
 sky130_fd_sc_hd__nor2_1 _4713_ (.A(_0222_),
    .B(_0238_),
    .Y(_0258_));
 sky130_fd_sc_hd__nand2_1 _4714_ (.A(_0215_),
    .B(_0258_),
    .Y(_0259_));
 sky130_fd_sc_hd__nand2_1 _4715_ (.A(_0259_),
    .B(_4173_),
    .Y(_0260_));
 sky130_fd_sc_hd__nand2_1 _4716_ (.A(_0260_),
    .B(_4162_),
    .Y(_0261_));
 sky130_fd_sc_hd__nand2_4 _4717_ (.A(\arbiter.master_sel[0][0] ),
    .B(\arbiter.master_sel[0][1] ),
    .Y(_0262_));
 sky130_fd_sc_hd__inv_6 _4718_ (.A(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__nand2_1 _4719_ (.A(_0263_),
    .B(_4108_),
    .Y(_0264_));
 sky130_fd_sc_hd__nor2_1 _4720_ (.A(_0264_),
    .B(_0229_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand2_1 _4721_ (.A(_4145_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__nand2_1 _4722_ (.A(_0266_),
    .B(\arbiter.master_handled[3] ),
    .Y(_0267_));
 sky130_fd_sc_hd__nand3_1 _4723_ (.A(_0261_),
    .B(net138),
    .C(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__nand2_1 _4724_ (.A(_0257_),
    .B(_0268_),
    .Y(_0269_));
 sky130_fd_sc_hd__nor2_1 _4725_ (.A(_0248_),
    .B(_0269_),
    .Y(_0270_));
 sky130_fd_sc_hd__o21ai_2 _4726_ (.A1(_0235_),
    .A2(_0237_),
    .B1(_0270_),
    .Y(_0271_));
 sky130_fd_sc_hd__nand3_1 _4727_ (.A(_0257_),
    .B(_0268_),
    .C(_0037_),
    .Y(_0272_));
 sky130_fd_sc_hd__nand2_1 _4728_ (.A(_0233_),
    .B(_0247_),
    .Y(_0273_));
 sky130_fd_sc_hd__inv_2 _4729_ (.A(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__a21oi_1 _4730_ (.A1(_0272_),
    .A2(_0274_),
    .B1(_4243_),
    .Y(_0275_));
 sky130_fd_sc_hd__nand2_1 _4731_ (.A(_0268_),
    .B(_4288_),
    .Y(_0276_));
 sky130_fd_sc_hd__nand2_1 _4732_ (.A(_0276_),
    .B(_0257_),
    .Y(_0277_));
 sky130_fd_sc_hd__nand2_1 _4733_ (.A(_0277_),
    .B(_0247_),
    .Y(_0278_));
 sky130_fd_sc_hd__nand2_1 _4734_ (.A(_0278_),
    .B(_0233_),
    .Y(_0279_));
 sky130_fd_sc_hd__nand3_1 _4735_ (.A(_0271_),
    .B(_0275_),
    .C(_0279_),
    .Y(_0280_));
 sky130_fd_sc_hd__nand2_1 _4736_ (.A(_0227_),
    .B(_0232_),
    .Y(_0281_));
 sky130_fd_sc_hd__inv_2 _4737_ (.A(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__nand2_1 _4738_ (.A(_0280_),
    .B(_0282_),
    .Y(_0283_));
 sky130_fd_sc_hd__inv_2 _4739_ (.A(_0041_),
    .Y(_0284_));
 sky130_fd_sc_hd__nor2_1 _4740_ (.A(\arbiter.state[1][0] ),
    .B(_0039_),
    .Y(_0285_));
 sky130_fd_sc_hd__a31o_1 _4741_ (.A1(_4286_),
    .A2(_0284_),
    .A3(_0285_),
    .B1(_0282_),
    .X(_0286_));
 sky130_fd_sc_hd__nor2_8 _4742_ (.A(net765),
    .B(_4233_),
    .Y(_0287_));
 sky130_fd_sc_hd__inv_6 _4743_ (.A(_0287_),
    .Y(_0288_));
 sky130_fd_sc_hd__nand2_1 _4744_ (.A(_0286_),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__nand2_1 _4745_ (.A(_0283_),
    .B(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__nand2_1 _4746_ (.A(_0290_),
    .B(_4150_),
    .Y(_0291_));
 sky130_fd_sc_hd__nand2_1 _4747_ (.A(_0291_),
    .B(_4239_),
    .Y(_0292_));
 sky130_fd_sc_hd__nand2_1 _4748_ (.A(_0291_),
    .B(_4240_),
    .Y(_0293_));
 sky130_fd_sc_hd__inv_2 _4749_ (.A(_0279_),
    .Y(_0294_));
 sky130_fd_sc_hd__nand3_1 _4750_ (.A(_0294_),
    .B(_0271_),
    .C(_0275_),
    .Y(_0295_));
 sky130_fd_sc_hd__and2_1 _4751_ (.A(_0242_),
    .B(_0246_),
    .X(_0296_));
 sky130_fd_sc_hd__nand2_1 _4752_ (.A(_0295_),
    .B(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__inv_2 _4753_ (.A(_0038_),
    .Y(_0298_));
 sky130_fd_sc_hd__nor2_1 _4754_ (.A(\arbiter.state[1][0] ),
    .B(_0041_),
    .Y(_0299_));
 sky130_fd_sc_hd__a31o_1 _4755_ (.A1(_4286_),
    .A2(_0298_),
    .A3(_0299_),
    .B1(_0296_),
    .X(_0300_));
 sky130_fd_sc_hd__nand2_1 _4756_ (.A(_0300_),
    .B(_0288_),
    .Y(_0301_));
 sky130_fd_sc_hd__nand2_1 _4757_ (.A(_0297_),
    .B(_0301_),
    .Y(_0302_));
 sky130_fd_sc_hd__nand2_1 _4758_ (.A(_0302_),
    .B(net11),
    .Y(_0303_));
 sky130_fd_sc_hd__nand2_1 _4759_ (.A(_0272_),
    .B(_0274_),
    .Y(_0304_));
 sky130_fd_sc_hd__nor2_1 _4760_ (.A(_4243_),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__nand3_1 _4761_ (.A(_0294_),
    .B(_0271_),
    .C(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__nand2_1 _4762_ (.A(_0261_),
    .B(_0267_),
    .Y(_0307_));
 sky130_fd_sc_hd__inv_2 _4763_ (.A(_0307_),
    .Y(_0308_));
 sky130_fd_sc_hd__nand2_1 _4764_ (.A(_0306_),
    .B(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__nor2_1 _4765_ (.A(\arbiter.state[1][0] ),
    .B(_0036_),
    .Y(_0310_));
 sky130_fd_sc_hd__a31o_1 _4766_ (.A1(_4286_),
    .A2(_0284_),
    .A3(_0310_),
    .B1(_0308_),
    .X(_0311_));
 sky130_fd_sc_hd__nand2_1 _4767_ (.A(_0311_),
    .B(_0288_),
    .Y(_0312_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(_0309_),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__nand2_1 _4769_ (.A(_0313_),
    .B(net138),
    .Y(_0314_));
 sky130_fd_sc_hd__nand3_1 _4770_ (.A(_0271_),
    .B(_0305_),
    .C(_0279_),
    .Y(_0315_));
 sky130_fd_sc_hd__nand2_1 _4771_ (.A(_0252_),
    .B(_0256_),
    .Y(_0316_));
 sky130_fd_sc_hd__inv_2 _4772_ (.A(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__nand2_1 _4773_ (.A(_0315_),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__inv_2 _4774_ (.A(_4289_),
    .Y(_0319_));
 sky130_fd_sc_hd__a31o_1 _4775_ (.A1(_4286_),
    .A2(_0319_),
    .A3(_0299_),
    .B1(_0317_),
    .X(_0320_));
 sky130_fd_sc_hd__nand2_1 _4776_ (.A(_0320_),
    .B(_0288_),
    .Y(_0321_));
 sky130_fd_sc_hd__nand2_1 _4777_ (.A(_0318_),
    .B(_0321_),
    .Y(_0322_));
 sky130_fd_sc_hd__nand2_1 _4778_ (.A(_0322_),
    .B(net74),
    .Y(_0323_));
 sky130_fd_sc_hd__nand3_2 _4779_ (.A(_0303_),
    .B(_0314_),
    .C(_0323_),
    .Y(_0324_));
 sky130_fd_sc_hd__a21oi_1 _4780_ (.A1(_0292_),
    .A2(_0293_),
    .B1(_0324_),
    .Y(_0325_));
 sky130_fd_sc_hd__nand2_1 _4781_ (.A(_0314_),
    .B(_0125_),
    .Y(_0326_));
 sky130_fd_sc_hd__nand2_1 _4782_ (.A(_0326_),
    .B(_0323_),
    .Y(_0327_));
 sky130_fd_sc_hd__nand2_1 _4783_ (.A(_0327_),
    .B(_0303_),
    .Y(_0328_));
 sky130_fd_sc_hd__nand2_1 _4784_ (.A(_0328_),
    .B(_0291_),
    .Y(_0329_));
 sky130_fd_sc_hd__nor2_1 _4785_ (.A(_0325_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__nand2_1 _4786_ (.A(_0303_),
    .B(_0291_),
    .Y(_0331_));
 sky130_fd_sc_hd__inv_2 _4787_ (.A(_0331_),
    .Y(_0332_));
 sky130_fd_sc_hd__nand3_1 _4788_ (.A(_0314_),
    .B(_0323_),
    .C(_0120_),
    .Y(_0333_));
 sky130_fd_sc_hd__nand2_1 _4789_ (.A(_0332_),
    .B(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__nor2_1 _4790_ (.A(_0094_),
    .B(_0334_),
    .Y(_0335_));
 sky130_fd_sc_hd__nand2_1 _4791_ (.A(_0330_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__nand2_1 _4792_ (.A(_0336_),
    .B(_0313_),
    .Y(_0337_));
 sky130_fd_sc_hd__inv_2 _4793_ (.A(_0131_),
    .Y(_0338_));
 sky130_fd_sc_hd__nor2_1 _4794_ (.A(net762),
    .B(_0123_),
    .Y(_0339_));
 sky130_fd_sc_hd__a31o_1 _4795_ (.A1(_0118_),
    .A2(_0338_),
    .A3(_0339_),
    .B1(_0313_),
    .X(_0340_));
 sky130_fd_sc_hd__nor2_1 _4796_ (.A(net762),
    .B(_4239_),
    .Y(_0341_));
 sky130_fd_sc_hd__inv_2 _4797_ (.A(_0341_),
    .Y(_0342_));
 sky130_fd_sc_hd__nand2_1 _4798_ (.A(_0340_),
    .B(_0342_),
    .Y(_0343_));
 sky130_fd_sc_hd__nand2_1 _4799_ (.A(_0337_),
    .B(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__nand2_1 _4800_ (.A(_0344_),
    .B(net138),
    .Y(_0345_));
 sky130_fd_sc_hd__a21oi_1 _4801_ (.A1(_0290_),
    .A2(_4150_),
    .B1(_0083_),
    .Y(_0346_));
 sky130_fd_sc_hd__inv_2 _4802_ (.A(_0293_),
    .Y(_0347_));
 sky130_fd_sc_hd__inv_2 _4803_ (.A(_0324_),
    .Y(_0348_));
 sky130_fd_sc_hd__o21ai_1 _4804_ (.A1(_0346_),
    .A2(_0347_),
    .B1(_0348_),
    .Y(_0349_));
 sky130_fd_sc_hd__nand3_1 _4805_ (.A(_0349_),
    .B(_0335_),
    .C(_0329_),
    .Y(_0350_));
 sky130_fd_sc_hd__nand2_1 _4806_ (.A(_0350_),
    .B(_0322_),
    .Y(_0351_));
 sky130_fd_sc_hd__a41o_1 _4807_ (.A1(_0118_),
    .A2(_4240_),
    .A3(_0121_),
    .A4(_0338_),
    .B1(_0322_),
    .X(_0352_));
 sky130_fd_sc_hd__nand2_1 _4808_ (.A(_0352_),
    .B(_0342_),
    .Y(_0353_));
 sky130_fd_sc_hd__nand2_1 _4809_ (.A(_0351_),
    .B(_0353_),
    .Y(_0354_));
 sky130_fd_sc_hd__nand2_1 _4810_ (.A(_0354_),
    .B(net74),
    .Y(_0355_));
 sky130_fd_sc_hd__nand2_1 _4811_ (.A(_0345_),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__a21oi_1 _4812_ (.A1(_0332_),
    .A2(_0333_),
    .B1(_0094_),
    .Y(_0357_));
 sky130_fd_sc_hd__nand3_1 _4813_ (.A(_0357_),
    .B(_0349_),
    .C(_0329_),
    .Y(_0358_));
 sky130_fd_sc_hd__nand2_1 _4814_ (.A(_0358_),
    .B(_0290_),
    .Y(_0359_));
 sky130_fd_sc_hd__a31o_1 _4815_ (.A1(_0118_),
    .A2(_4240_),
    .A3(_0129_),
    .B1(_0290_),
    .X(_0360_));
 sky130_fd_sc_hd__nand2_1 _4816_ (.A(_0360_),
    .B(_0342_),
    .Y(_0361_));
 sky130_fd_sc_hd__nand2_1 _4817_ (.A(_0359_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__nand2_1 _4818_ (.A(_0362_),
    .B(_4150_),
    .Y(_0363_));
 sky130_fd_sc_hd__nand3_1 _4819_ (.A(_0330_),
    .B(_0341_),
    .C(_0357_),
    .Y(_0364_));
 sky130_fd_sc_hd__inv_8 _4820_ (.A(_0126_),
    .Y(_0365_));
 sky130_fd_sc_hd__nor2_1 _4821_ (.A(_0341_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__a41o_1 _4822_ (.A1(_0118_),
    .A2(_4240_),
    .A3(_0338_),
    .A4(_0366_),
    .B1(_0302_),
    .X(_0367_));
 sky130_fd_sc_hd__nand3_1 _4823_ (.A(_0364_),
    .B(net11),
    .C(_0367_),
    .Y(_0368_));
 sky130_fd_sc_hd__nand3_1 _4824_ (.A(_0363_),
    .B(_0166_),
    .C(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__nor2_1 _4825_ (.A(_0356_),
    .B(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__nor2_1 _4826_ (.A(_0211_),
    .B(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__nor2_1 _4827_ (.A(_0208_),
    .B(_0371_),
    .Y(_0372_));
 sky130_fd_sc_hd__nand2_1 _4828_ (.A(_0137_),
    .B(net751),
    .Y(_0373_));
 sky130_fd_sc_hd__o21ai_1 _4829_ (.A1(_0373_),
    .A2(_0165_),
    .B1(net740),
    .Y(_0374_));
 sky130_fd_sc_hd__nand2_1 _4830_ (.A(_0374_),
    .B(_0168_),
    .Y(_0375_));
 sky130_fd_sc_hd__nand2_1 _4831_ (.A(_0372_),
    .B(net752),
    .Y(_0022_));
 sky130_fd_sc_hd__nand2_1 _4832_ (.A(_0022_),
    .B(net740),
    .Y(_0376_));
 sky130_fd_sc_hd__nand2_1 _4833_ (.A(_0270_),
    .B(_0235_),
    .Y(_0377_));
 sky130_fd_sc_hd__a21o_1 _4834_ (.A1(_4222_),
    .A2(_4250_),
    .B1(_4243_),
    .X(_0378_));
 sky130_fd_sc_hd__a32o_1 _4835_ (.A1(_4185_),
    .A2(_4286_),
    .A3(_0284_),
    .B1(_0378_),
    .B2(_4235_),
    .X(_0379_));
 sky130_fd_sc_hd__a31o_2 _4836_ (.A1(net743),
    .A2(_0287_),
    .A3(_0377_),
    .B1(_0379_),
    .X(_0026_));
 sky130_fd_sc_hd__nor2_1 _4837_ (.A(_0094_),
    .B(_0342_),
    .Y(_0380_));
 sky130_fd_sc_hd__o21a_1 _4838_ (.A1(_0293_),
    .A2(_0324_),
    .B1(_0380_),
    .X(_0381_));
 sky130_fd_sc_hd__nand2_1 _4839_ (.A(_0071_),
    .B(_0100_),
    .Y(_0382_));
 sky130_fd_sc_hd__a21o_1 _4840_ (.A1(_0382_),
    .A2(net734),
    .B1(_0134_),
    .X(_0383_));
 sky130_fd_sc_hd__nand2_1 _4841_ (.A(_0383_),
    .B(_0153_),
    .Y(_0384_));
 sky130_fd_sc_hd__nor2_2 _4842_ (.A(_0381_),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__o2bb2a_1 _4843_ (.A1_N(net743),
    .A2_N(_0026_),
    .B1(_0094_),
    .B2(_0385_),
    .X(_0386_));
 sky130_fd_sc_hd__nand2_1 _4844_ (.A(_0020_),
    .B(_0175_),
    .Y(_0387_));
 sky130_fd_sc_hd__nand3_4 _4845_ (.A(_0376_),
    .B(_0386_),
    .C(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__o21ai_1 _4846_ (.A1(_0180_),
    .A2(_0388_),
    .B1(net737),
    .Y(_0389_));
 sky130_fd_sc_hd__inv_4 _4847_ (.A(_0388_),
    .Y(_0390_));
 sky130_fd_sc_hd__inv_2 _4848_ (.A(_0180_),
    .Y(_0391_));
 sky130_fd_sc_hd__inv_2 _4849_ (.A(_0023_),
    .Y(_0392_));
 sky130_fd_sc_hd__nand3_1 _4850_ (.A(_0392_),
    .B(_0372_),
    .C(_0375_),
    .Y(_0393_));
 sky130_fd_sc_hd__nand2_1 _4851_ (.A(_0385_),
    .B(_0086_),
    .Y(_0394_));
 sky130_fd_sc_hd__nor2_1 _4852_ (.A(_0021_),
    .B(_0020_),
    .Y(_0395_));
 sky130_fd_sc_hd__nor2_1 _4853_ (.A(_0027_),
    .B(_0026_),
    .Y(_0396_));
 sky130_fd_sc_hd__nor2_1 _4854_ (.A(_0395_),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__nand2_1 _4855_ (.A(_0394_),
    .B(_0397_),
    .Y(_0398_));
 sky130_fd_sc_hd__inv_2 _4856_ (.A(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__nand2_1 _4857_ (.A(_0393_),
    .B(_0399_),
    .Y(_0400_));
 sky130_fd_sc_hd__inv_2 _4858_ (.A(_0395_),
    .Y(_0401_));
 sky130_fd_sc_hd__nand2_1 _4859_ (.A(_0400_),
    .B(_0401_),
    .Y(_0402_));
 sky130_fd_sc_hd__nand3_1 _4860_ (.A(_0390_),
    .B(_0391_),
    .C(_0402_),
    .Y(_0403_));
 sky130_fd_sc_hd__nand2_1 _4861_ (.A(net738),
    .B(_0403_),
    .Y(_0000_));
 sky130_fd_sc_hd__o21ai_1 _4862_ (.A1(_0180_),
    .A2(_0388_),
    .B1(net734),
    .Y(_0404_));
 sky130_fd_sc_hd__and3_1 _4863_ (.A(_0385_),
    .B(_0086_),
    .C(_0397_),
    .X(_0405_));
 sky130_fd_sc_hd__nand3_1 _4864_ (.A(_0390_),
    .B(_0391_),
    .C(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__nand2_1 _4865_ (.A(net735),
    .B(_0406_),
    .Y(_0001_));
 sky130_fd_sc_hd__inv_2 _4866_ (.A(_0385_),
    .Y(_0024_));
 sky130_fd_sc_hd__buf_8 _4867_ (.A(_0039_),
    .X(_0407_));
 sky130_fd_sc_hd__buf_8 _4868_ (.A(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__buf_8 _4869_ (.A(_0038_),
    .X(_0409_));
 sky130_fd_sc_hd__clkbuf_16 _4870_ (.A(_0409_),
    .X(_0410_));
 sky130_fd_sc_hd__buf_6 _4871_ (.A(_0036_),
    .X(_0411_));
 sky130_fd_sc_hd__buf_6 _4872_ (.A(_0411_),
    .X(_0412_));
 sky130_fd_sc_hd__buf_6 _4873_ (.A(_4289_),
    .X(_0413_));
 sky130_fd_sc_hd__buf_8 _4874_ (.A(_0413_),
    .X(_0414_));
 sky130_fd_sc_hd__o22a_1 _4875_ (.A1(net80),
    .A2(_0412_),
    .B1(net17),
    .B2(_0414_),
    .X(_0415_));
 sky130_fd_sc_hd__o221a_2 _4876_ (.A1(net1),
    .A2(_0408_),
    .B1(net181),
    .B2(_0410_),
    .C1(_0415_),
    .X(_0416_));
 sky130_fd_sc_hd__nor2_8 _4877_ (.A(_4105_),
    .B(_0056_),
    .Y(_0417_));
 sky130_fd_sc_hd__inv_8 _4878_ (.A(_0417_),
    .Y(_0418_));
 sky130_fd_sc_hd__nor2_8 _4879_ (.A(_4184_),
    .B(_4263_),
    .Y(_0419_));
 sky130_fd_sc_hd__inv_6 _4880_ (.A(_0419_),
    .Y(_0420_));
 sky130_fd_sc_hd__nand2_4 _4881_ (.A(_0418_),
    .B(_0420_),
    .Y(_0421_));
 sky130_fd_sc_hd__buf_6 _4882_ (.A(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__inv_2 _4883_ (.A(net1),
    .Y(_0423_));
 sky130_fd_sc_hd__inv_6 _4884_ (.A(_4149_),
    .Y(_0424_));
 sky130_fd_sc_hd__clkbuf_8 _4885_ (.A(_0424_),
    .X(_0425_));
 sky130_fd_sc_hd__clkbuf_16 _4886_ (.A(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__buf_8 _4887_ (.A(_0426_),
    .X(_0427_));
 sky130_fd_sc_hd__inv_2 _4888_ (.A(net181),
    .Y(_0428_));
 sky130_fd_sc_hd__inv_6 _4889_ (.A(_4147_),
    .Y(_0429_));
 sky130_fd_sc_hd__clkbuf_8 _4890_ (.A(_0429_),
    .X(_0430_));
 sky130_fd_sc_hd__buf_8 _4891_ (.A(_0430_),
    .X(_0431_));
 sky130_fd_sc_hd__buf_8 _4892_ (.A(_0263_),
    .X(_0432_));
 sky130_fd_sc_hd__buf_8 _4893_ (.A(_0432_),
    .X(_0433_));
 sky130_fd_sc_hd__inv_6 _4894_ (.A(_0253_),
    .Y(_0434_));
 sky130_fd_sc_hd__buf_8 _4895_ (.A(_0434_),
    .X(_0435_));
 sky130_fd_sc_hd__buf_12 _4896_ (.A(_0435_),
    .X(_0436_));
 sky130_fd_sc_hd__a22oi_1 _4897_ (.A1(_0433_),
    .A2(net80),
    .B1(_0436_),
    .B2(net17),
    .Y(_0437_));
 sky130_fd_sc_hd__o221a_2 _4898_ (.A1(_0423_),
    .A2(_0427_),
    .B1(_0428_),
    .B2(_0431_),
    .C1(_0437_),
    .X(_0438_));
 sky130_fd_sc_hd__inv_2 _4899_ (.A(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__inv_4 _4900_ (.A(_4112_),
    .Y(_0440_));
 sky130_fd_sc_hd__nor2_8 _4901_ (.A(_4105_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__inv_2 _4902_ (.A(_0441_),
    .Y(_0442_));
 sky130_fd_sc_hd__nor2_8 _4903_ (.A(_4158_),
    .B(_4223_),
    .Y(_0443_));
 sky130_fd_sc_hd__inv_2 _4904_ (.A(_0443_),
    .Y(_0444_));
 sky130_fd_sc_hd__nand2_1 _4905_ (.A(_0442_),
    .B(_0444_),
    .Y(_0445_));
 sky130_fd_sc_hd__inv_2 _4906_ (.A(_0445_),
    .Y(_0446_));
 sky130_fd_sc_hd__nor2_8 _4907_ (.A(_0421_),
    .B(_0446_),
    .Y(_0447_));
 sky130_fd_sc_hd__a22o_1 _4908_ (.A1(_0416_),
    .A2(_0422_),
    .B1(_0439_),
    .B2(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__buf_8 _4909_ (.A(_0128_),
    .X(_0449_));
 sky130_fd_sc_hd__buf_12 _4910_ (.A(_0449_),
    .X(_0450_));
 sky130_fd_sc_hd__clkbuf_16 _4911_ (.A(_0450_),
    .X(_0451_));
 sky130_fd_sc_hd__buf_8 _4912_ (.A(_0365_),
    .X(_0452_));
 sky130_fd_sc_hd__buf_8 _4913_ (.A(_0452_),
    .X(_0453_));
 sky130_fd_sc_hd__buf_8 _4914_ (.A(_0123_),
    .X(_0454_));
 sky130_fd_sc_hd__buf_8 _4915_ (.A(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__clkbuf_8 _4916_ (.A(_0122_),
    .X(_0456_));
 sky130_fd_sc_hd__buf_8 _4917_ (.A(_0456_),
    .X(_0457_));
 sky130_fd_sc_hd__o22a_1 _4918_ (.A1(net80),
    .A2(_0455_),
    .B1(net17),
    .B2(_0457_),
    .X(_0458_));
 sky130_fd_sc_hd__o221a_2 _4919_ (.A1(net1),
    .A2(_0451_),
    .B1(net181),
    .B2(_0453_),
    .C1(_0458_),
    .X(_0459_));
 sky130_fd_sc_hd__nor2_4 _4920_ (.A(_4105_),
    .B(_0134_),
    .Y(_0460_));
 sky130_fd_sc_hd__clkinv_4 _4921_ (.A(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__nor2_4 _4922_ (.A(_0083_),
    .B(_0107_),
    .Y(_0462_));
 sky130_fd_sc_hd__inv_2 _4923_ (.A(_0462_),
    .Y(_0463_));
 sky130_fd_sc_hd__nand2_2 _4924_ (.A(_0461_),
    .B(_0463_),
    .Y(_0464_));
 sky130_fd_sc_hd__buf_8 _4925_ (.A(_0464_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _4926_ (.A0(_0448_),
    .A1(_0459_),
    .S(_0465_),
    .X(_0466_));
 sky130_fd_sc_hd__clkbuf_16 _4927_ (.A(_0182_),
    .X(_0467_));
 sky130_fd_sc_hd__buf_8 _4928_ (.A(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__buf_12 _4929_ (.A(_0468_),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_16 _4930_ (.A(_0469_),
    .X(_0470_));
 sky130_fd_sc_hd__buf_8 _4931_ (.A(_0185_),
    .X(_0471_));
 sky130_fd_sc_hd__buf_8 _4932_ (.A(_0471_),
    .X(_0472_));
 sky130_fd_sc_hd__buf_12 _4933_ (.A(_0472_),
    .X(_0473_));
 sky130_fd_sc_hd__clkbuf_8 _4934_ (.A(_0186_),
    .X(_0474_));
 sky130_fd_sc_hd__buf_12 _4935_ (.A(_0474_),
    .X(_0475_));
 sky130_fd_sc_hd__buf_8 _4936_ (.A(_0475_),
    .X(_0476_));
 sky130_fd_sc_hd__clkbuf_8 _4937_ (.A(_0189_),
    .X(_0477_));
 sky130_fd_sc_hd__clkbuf_8 _4938_ (.A(_0477_),
    .X(_0478_));
 sky130_fd_sc_hd__buf_6 _4939_ (.A(_0478_),
    .X(_0479_));
 sky130_fd_sc_hd__buf_8 _4940_ (.A(_0479_),
    .X(_0480_));
 sky130_fd_sc_hd__o22a_1 _4941_ (.A1(net80),
    .A2(_0476_),
    .B1(net17),
    .B2(_0480_),
    .X(_0481_));
 sky130_fd_sc_hd__o221a_2 _4942_ (.A1(net1),
    .A2(_0470_),
    .B1(net181),
    .B2(_0473_),
    .C1(_0481_),
    .X(_0482_));
 sky130_fd_sc_hd__inv_6 _4943_ (.A(_0167_),
    .Y(_0483_));
 sky130_fd_sc_hd__nor2_2 _4944_ (.A(_4105_),
    .B(_0483_),
    .Y(_0484_));
 sky130_fd_sc_hd__inv_2 _4945_ (.A(_0484_),
    .Y(_0485_));
 sky130_fd_sc_hd__clkbuf_16 _4946_ (.A(_0193_),
    .X(_0486_));
 sky130_fd_sc_hd__nor2_4 _4947_ (.A(_0138_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__inv_2 _4948_ (.A(_0487_),
    .Y(_0488_));
 sky130_fd_sc_hd__nand2_4 _4949_ (.A(_0485_),
    .B(_0488_),
    .Y(_0489_));
 sky130_fd_sc_hd__clkbuf_8 _4950_ (.A(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__mux2_1 _4951_ (.A0(_0466_),
    .A1(_0482_),
    .S(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__buf_1 _4952_ (.A(_0491_),
    .X(net581));
 sky130_fd_sc_hd__buf_8 _4953_ (.A(_0039_),
    .X(_0492_));
 sky130_fd_sc_hd__o22a_1 _4954_ (.A1(net81),
    .A2(_0411_),
    .B1(net18),
    .B2(_0413_),
    .X(_0493_));
 sky130_fd_sc_hd__o221a_4 _4955_ (.A1(net112),
    .A2(_0492_),
    .B1(net182),
    .B2(_0409_),
    .C1(_0493_),
    .X(_0494_));
 sky130_fd_sc_hd__inv_2 _4956_ (.A(net112),
    .Y(_0495_));
 sky130_fd_sc_hd__inv_2 _4957_ (.A(net182),
    .Y(_0496_));
 sky130_fd_sc_hd__a22oi_1 _4958_ (.A1(_0432_),
    .A2(net81),
    .B1(_0435_),
    .B2(net18),
    .Y(_0497_));
 sky130_fd_sc_hd__o221a_2 _4959_ (.A1(_0495_),
    .A2(_0426_),
    .B1(_0496_),
    .B2(_0431_),
    .C1(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__inv_2 _4960_ (.A(_0498_),
    .Y(_0499_));
 sky130_fd_sc_hd__a22o_1 _4961_ (.A1(_0494_),
    .A2(_0422_),
    .B1(_0499_),
    .B2(_0447_),
    .X(_0500_));
 sky130_fd_sc_hd__o22a_1 _4962_ (.A1(net81),
    .A2(_0455_),
    .B1(net18),
    .B2(_0457_),
    .X(_0501_));
 sky130_fd_sc_hd__o221a_2 _4963_ (.A1(net112),
    .A2(_0451_),
    .B1(net182),
    .B2(_0453_),
    .C1(_0501_),
    .X(_0502_));
 sky130_fd_sc_hd__mux2_1 _4964_ (.A0(_0500_),
    .A1(_0502_),
    .S(_0465_),
    .X(_0503_));
 sky130_fd_sc_hd__o22a_1 _4965_ (.A1(net81),
    .A2(_0476_),
    .B1(net18),
    .B2(_0480_),
    .X(_0504_));
 sky130_fd_sc_hd__o221a_2 _4966_ (.A1(net112),
    .A2(_0470_),
    .B1(net182),
    .B2(_0473_),
    .C1(_0504_),
    .X(_0505_));
 sky130_fd_sc_hd__mux2_1 _4967_ (.A0(_0503_),
    .A1(_0505_),
    .S(_0490_),
    .X(_0506_));
 sky130_fd_sc_hd__buf_1 _4968_ (.A(_0506_),
    .X(net582));
 sky130_fd_sc_hd__o22a_1 _4969_ (.A1(net82),
    .A2(_0411_),
    .B1(net19),
    .B2(_0413_),
    .X(_0507_));
 sky130_fd_sc_hd__o221a_2 _4970_ (.A1(net151),
    .A2(_0407_),
    .B1(net183),
    .B2(_0409_),
    .C1(_0507_),
    .X(_0508_));
 sky130_fd_sc_hd__nand2_1 _4971_ (.A(_0508_),
    .B(_4272_),
    .Y(_0509_));
 sky130_fd_sc_hd__buf_8 _4972_ (.A(_4252_),
    .X(_0510_));
 sky130_fd_sc_hd__nand2_1 _4973_ (.A(_0509_),
    .B(_0510_),
    .Y(_0511_));
 sky130_fd_sc_hd__inv_2 _4974_ (.A(_0421_),
    .Y(_0512_));
 sky130_fd_sc_hd__inv_2 _4975_ (.A(net151),
    .Y(_0513_));
 sky130_fd_sc_hd__inv_2 _4976_ (.A(net183),
    .Y(_0514_));
 sky130_fd_sc_hd__nand2_1 _4977_ (.A(_4153_),
    .B(net19),
    .Y(_0515_));
 sky130_fd_sc_hd__nand2_1 _4978_ (.A(\arbiter.master_sel[0][0] ),
    .B(net82),
    .Y(_0516_));
 sky130_fd_sc_hd__a21o_1 _4979_ (.A1(_0515_),
    .A2(_0516_),
    .B1(_4156_),
    .X(_0517_));
 sky130_fd_sc_hd__o221a_1 _4980_ (.A1(_0513_),
    .A2(_0426_),
    .B1(_0514_),
    .B2(_0431_),
    .C1(_0517_),
    .X(_0518_));
 sky130_fd_sc_hd__inv_2 _4981_ (.A(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__inv_6 _4982_ (.A(_4204_),
    .Y(_0520_));
 sky130_fd_sc_hd__nand2_1 _4983_ (.A(_0519_),
    .B(_0520_),
    .Y(_0521_));
 sky130_fd_sc_hd__buf_6 _4984_ (.A(_4127_),
    .X(_0522_));
 sky130_fd_sc_hd__buf_8 _4985_ (.A(_0522_),
    .X(_0523_));
 sky130_fd_sc_hd__nand2_1 _4986_ (.A(_0521_),
    .B(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__nor2_2 _4987_ (.A(_4235_),
    .B(_0419_),
    .Y(_0525_));
 sky130_fd_sc_hd__a32o_1 _4988_ (.A1(_0519_),
    .A2(_0441_),
    .A3(_0525_),
    .B1(_0417_),
    .B2(_0508_),
    .X(_0526_));
 sky130_fd_sc_hd__a31o_1 _4989_ (.A1(_0512_),
    .A2(_0443_),
    .A3(_0524_),
    .B1(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__a31o_1 _4990_ (.A1(_4233_),
    .A2(_4268_),
    .A3(_0511_),
    .B1(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__o22a_1 _4991_ (.A1(net82),
    .A2(_0455_),
    .B1(net19),
    .B2(_0457_),
    .X(_0529_));
 sky130_fd_sc_hd__o221a_2 _4992_ (.A1(net151),
    .A2(_0451_),
    .B1(net183),
    .B2(_0453_),
    .C1(_0529_),
    .X(_0530_));
 sky130_fd_sc_hd__mux2_1 _4993_ (.A0(_0528_),
    .A1(_0530_),
    .S(_0465_),
    .X(_0531_));
 sky130_fd_sc_hd__o22a_1 _4994_ (.A1(net82),
    .A2(_0476_),
    .B1(net19),
    .B2(_0480_),
    .X(_0532_));
 sky130_fd_sc_hd__o221a_2 _4995_ (.A1(net151),
    .A2(_0470_),
    .B1(net183),
    .B2(_0473_),
    .C1(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__mux2_1 _4996_ (.A0(_0531_),
    .A1(_0533_),
    .S(_0490_),
    .X(_0534_));
 sky130_fd_sc_hd__buf_1 _4997_ (.A(_0534_),
    .X(net583));
 sky130_fd_sc_hd__buf_8 _4998_ (.A(_0465_),
    .X(_0535_));
 sky130_fd_sc_hd__o22a_1 _4999_ (.A1(net83),
    .A2(_0455_),
    .B1(net20),
    .B2(_0457_),
    .X(_0536_));
 sky130_fd_sc_hd__o221a_2 _5000_ (.A1(net185),
    .A2(_0453_),
    .B1(net162),
    .B2(_0451_),
    .C1(_0536_),
    .X(_0537_));
 sky130_fd_sc_hd__buf_12 _5001_ (.A(_4204_),
    .X(_0538_));
 sky130_fd_sc_hd__buf_12 _5002_ (.A(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__inv_2 _5003_ (.A(net185),
    .Y(_0540_));
 sky130_fd_sc_hd__inv_2 _5004_ (.A(net162),
    .Y(_0541_));
 sky130_fd_sc_hd__a22oi_1 _5005_ (.A1(_0432_),
    .A2(net83),
    .B1(_0435_),
    .B2(net20),
    .Y(_0542_));
 sky130_fd_sc_hd__o221a_2 _5006_ (.A1(_0540_),
    .A2(_0431_),
    .B1(_0541_),
    .B2(_0426_),
    .C1(_0542_),
    .X(_0543_));
 sky130_fd_sc_hd__nor2_1 _5007_ (.A(_0539_),
    .B(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__nand2_1 _5008_ (.A(_0544_),
    .B(_0523_),
    .Y(_0545_));
 sky130_fd_sc_hd__o21ai_1 _5009_ (.A1(_0523_),
    .A2(_0521_),
    .B1(_0545_),
    .Y(_0546_));
 sky130_fd_sc_hd__nand2_1 _5010_ (.A(_0546_),
    .B(_0443_),
    .Y(_0547_));
 sky130_fd_sc_hd__inv_2 _5011_ (.A(_0525_),
    .Y(_0548_));
 sky130_fd_sc_hd__nor2_1 _5012_ (.A(_0442_),
    .B(_0543_),
    .Y(_0549_));
 sky130_fd_sc_hd__nand2_4 _5013_ (.A(_4235_),
    .B(_4105_),
    .Y(_0550_));
 sky130_fd_sc_hd__o21ai_1 _5014_ (.A1(_0548_),
    .A2(_0549_),
    .B1(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__o22a_1 _5015_ (.A1(net83),
    .A2(_0411_),
    .B1(net20),
    .B2(_0413_),
    .X(_0552_));
 sky130_fd_sc_hd__o221a_2 _5016_ (.A1(net185),
    .A2(_0409_),
    .B1(net162),
    .B2(_0492_),
    .C1(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__nor2_1 _5017_ (.A(_0418_),
    .B(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__buf_8 _5018_ (.A(_4253_),
    .X(_0555_));
 sky130_fd_sc_hd__nand2_1 _5019_ (.A(_0553_),
    .B(_4272_),
    .Y(_0556_));
 sky130_fd_sc_hd__buf_8 _5020_ (.A(_0510_),
    .X(_0557_));
 sky130_fd_sc_hd__buf_8 _5021_ (.A(_0557_),
    .X(_0558_));
 sky130_fd_sc_hd__or2_1 _5022_ (.A(_0558_),
    .B(_0509_),
    .X(_0559_));
 sky130_fd_sc_hd__o21ai_1 _5023_ (.A1(_0555_),
    .A2(_0556_),
    .B1(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__nor2_1 _5024_ (.A(_0420_),
    .B(_0560_),
    .Y(_0561_));
 sky130_fd_sc_hd__a2111o_1 _5025_ (.A1(_0547_),
    .A2(_0551_),
    .B1(_0464_),
    .C1(_0554_),
    .D1(_0561_),
    .X(_0562_));
 sky130_fd_sc_hd__a21bo_1 _5026_ (.A1(_0535_),
    .A2(_0537_),
    .B1_N(_0562_),
    .X(_0563_));
 sky130_fd_sc_hd__o22a_1 _5027_ (.A1(net83),
    .A2(_0476_),
    .B1(net20),
    .B2(_0480_),
    .X(_0564_));
 sky130_fd_sc_hd__o221a_2 _5028_ (.A1(net185),
    .A2(_0473_),
    .B1(net162),
    .B2(_0470_),
    .C1(_0564_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_1 _5029_ (.A0(_0563_),
    .A1(_0565_),
    .S(_0490_),
    .X(_0566_));
 sky130_fd_sc_hd__buf_1 _5030_ (.A(_0566_),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_8 _5031_ (.A(_0490_),
    .X(_0567_));
 sky130_fd_sc_hd__o22a_1 _5032_ (.A1(net84),
    .A2(_0476_),
    .B1(net21),
    .B2(_0479_),
    .X(_0568_));
 sky130_fd_sc_hd__o221a_2 _5033_ (.A1(net173),
    .A2(_0470_),
    .B1(net186),
    .B2(_0473_),
    .C1(_0568_),
    .X(_0569_));
 sky130_fd_sc_hd__o22a_1 _5034_ (.A1(net84),
    .A2(_0455_),
    .B1(net21),
    .B2(_0456_),
    .X(_0570_));
 sky130_fd_sc_hd__o221a_4 _5035_ (.A1(net173),
    .A2(_0450_),
    .B1(net186),
    .B2(_0452_),
    .C1(_0570_),
    .X(_0571_));
 sky130_fd_sc_hd__clkbuf_16 _5036_ (.A(_0111_),
    .X(_0572_));
 sky130_fd_sc_hd__o22a_1 _5037_ (.A1(net85),
    .A2(_0455_),
    .B1(net22),
    .B2(_0456_),
    .X(_0573_));
 sky130_fd_sc_hd__o221a_4 _5038_ (.A1(net184),
    .A2(_0450_),
    .B1(net187),
    .B2(_0452_),
    .C1(_0573_),
    .X(_0574_));
 sky130_fd_sc_hd__o22a_1 _5039_ (.A1(net86),
    .A2(_0454_),
    .B1(net24),
    .B2(_0456_),
    .X(_0575_));
 sky130_fd_sc_hd__o221a_4 _5040_ (.A1(net195),
    .A2(_0450_),
    .B1(net188),
    .B2(_0452_),
    .C1(_0575_),
    .X(_0576_));
 sky130_fd_sc_hd__inv_2 _5041_ (.A(_0576_),
    .Y(_0577_));
 sky130_fd_sc_hd__nor2_1 _5042_ (.A(_0110_),
    .B(_0577_),
    .Y(_0578_));
 sky130_fd_sc_hd__a221o_1 _5043_ (.A1(_0571_),
    .A2(_0108_),
    .B1(_0572_),
    .B2(_0574_),
    .C1(_0578_),
    .X(_0579_));
 sky130_fd_sc_hd__o22a_1 _5044_ (.A1(net84),
    .A2(_0411_),
    .B1(net21),
    .B2(_0413_),
    .X(_0580_));
 sky130_fd_sc_hd__o221a_2 _5045_ (.A1(net173),
    .A2(_0492_),
    .B1(net186),
    .B2(_0409_),
    .C1(_0580_),
    .X(_0581_));
 sky130_fd_sc_hd__inv_2 _5046_ (.A(net173),
    .Y(_0582_));
 sky130_fd_sc_hd__inv_2 _5047_ (.A(net186),
    .Y(_0583_));
 sky130_fd_sc_hd__a22oi_1 _5048_ (.A1(_0432_),
    .A2(net84),
    .B1(_0435_),
    .B2(net21),
    .Y(_0584_));
 sky130_fd_sc_hd__o221a_1 _5049_ (.A1(_0582_),
    .A2(_0426_),
    .B1(_0583_),
    .B2(_0431_),
    .C1(_0584_),
    .X(_0585_));
 sky130_fd_sc_hd__inv_2 _5050_ (.A(_0585_),
    .Y(_0586_));
 sky130_fd_sc_hd__mux2_1 _5051_ (.A0(_0544_),
    .A1(_0586_),
    .S(_0523_),
    .X(_0587_));
 sky130_fd_sc_hd__clkbuf_16 _5052_ (.A(\arbiter.state[0][1] ),
    .X(_0588_));
 sky130_fd_sc_hd__buf_8 _5053_ (.A(_0588_),
    .X(_0589_));
 sky130_fd_sc_hd__inv_8 _5054_ (.A(_4223_),
    .Y(_0590_));
 sky130_fd_sc_hd__clkbuf_8 _5055_ (.A(_0442_),
    .X(_0591_));
 sky130_fd_sc_hd__buf_6 _5056_ (.A(_0512_),
    .X(_0592_));
 sky130_fd_sc_hd__o21ai_1 _5057_ (.A1(_0591_),
    .A2(_0585_),
    .B1(_0592_),
    .Y(_0593_));
 sky130_fd_sc_hd__a31o_1 _5058_ (.A1(_0587_),
    .A2(_0589_),
    .A3(_0590_),
    .B1(_0593_),
    .X(_0594_));
 sky130_fd_sc_hd__inv_2 _5059_ (.A(_0581_),
    .Y(_0595_));
 sky130_fd_sc_hd__or2_1 _5060_ (.A(_0557_),
    .B(_0556_),
    .X(_0596_));
 sky130_fd_sc_hd__o21ai_4 _5061_ (.A1(_0555_),
    .A2(_0595_),
    .B1(_0596_),
    .Y(_0597_));
 sky130_fd_sc_hd__or4_4 _5062_ (.A(_4184_),
    .B(_0555_),
    .C(_4245_),
    .D(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__o211a_1 _5063_ (.A1(_0418_),
    .A2(_0581_),
    .B1(_0594_),
    .C1(_0598_),
    .X(_0599_));
 sky130_fd_sc_hd__or2_1 _5064_ (.A(_0461_),
    .B(_0571_),
    .X(_0600_));
 sky130_fd_sc_hd__inv_4 _5065_ (.A(_0489_),
    .Y(_0601_));
 sky130_fd_sc_hd__and2_1 _5066_ (.A(_0600_),
    .B(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__o221a_1 _5067_ (.A1(_0463_),
    .A2(_0579_),
    .B1(_0535_),
    .B2(_0599_),
    .C1(_0602_),
    .X(_0603_));
 sky130_fd_sc_hd__a21o_1 _5068_ (.A1(_0567_),
    .A2(_0569_),
    .B1(_0603_),
    .X(net585));
 sky130_fd_sc_hd__buf_6 _5069_ (.A(_0592_),
    .X(_0604_));
 sky130_fd_sc_hd__inv_2 _5070_ (.A(net184),
    .Y(_0605_));
 sky130_fd_sc_hd__inv_2 _5071_ (.A(net187),
    .Y(_0606_));
 sky130_fd_sc_hd__a22oi_1 _5072_ (.A1(_0433_),
    .A2(net85),
    .B1(_0436_),
    .B2(net22),
    .Y(_0607_));
 sky130_fd_sc_hd__o221a_2 _5073_ (.A1(_0605_),
    .A2(_0426_),
    .B1(_0606_),
    .B2(_0431_),
    .C1(_0607_),
    .X(_0608_));
 sky130_fd_sc_hd__inv_2 _5074_ (.A(_0608_),
    .Y(_0609_));
 sky130_fd_sc_hd__nor2_1 _5075_ (.A(_0591_),
    .B(_0608_),
    .Y(_0610_));
 sky130_fd_sc_hd__a31o_1 _5076_ (.A1(_0609_),
    .A2(_0589_),
    .A3(_0590_),
    .B1(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__clkbuf_16 _5077_ (.A(_4265_),
    .X(_0612_));
 sky130_fd_sc_hd__buf_8 _5078_ (.A(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__clkbuf_16 _5079_ (.A(_4287_),
    .X(_0614_));
 sky130_fd_sc_hd__buf_8 _5080_ (.A(_0408_),
    .X(_0615_));
 sky130_fd_sc_hd__o22a_1 _5081_ (.A1(net86),
    .A2(_0412_),
    .B1(net24),
    .B2(_0414_),
    .X(_0616_));
 sky130_fd_sc_hd__o221ai_4 _5082_ (.A1(net195),
    .A2(_0615_),
    .B1(net188),
    .B2(_0410_),
    .C1(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__o22a_1 _5083_ (.A1(net87),
    .A2(_0412_),
    .B1(net25),
    .B2(_0414_),
    .X(_0618_));
 sky130_fd_sc_hd__o221ai_4 _5084_ (.A1(net206),
    .A2(_0408_),
    .B1(net189),
    .B2(_0410_),
    .C1(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__o22a_1 _5085_ (.A1(net85),
    .A2(_0412_),
    .B1(net22),
    .B2(_0414_),
    .X(_0620_));
 sky130_fd_sc_hd__o221a_2 _5086_ (.A1(net184),
    .A2(_0408_),
    .B1(net187),
    .B2(_0410_),
    .C1(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__nand2_1 _5087_ (.A(_0621_),
    .B(_4268_),
    .Y(_0622_));
 sky130_fd_sc_hd__o221a_1 _5088_ (.A1(_0614_),
    .A2(_0617_),
    .B1(_4271_),
    .B2(_0619_),
    .C1(_0622_),
    .X(_0623_));
 sky130_fd_sc_hd__buf_8 _5089_ (.A(_0038_),
    .X(_0624_));
 sky130_fd_sc_hd__buf_8 _5090_ (.A(_0411_),
    .X(_0625_));
 sky130_fd_sc_hd__buf_6 _5091_ (.A(_4289_),
    .X(_0626_));
 sky130_fd_sc_hd__o22a_1 _5092_ (.A1(net95),
    .A2(_0625_),
    .B1(net32),
    .B2(_0626_),
    .X(_0627_));
 sky130_fd_sc_hd__o221a_4 _5093_ (.A1(net56),
    .A2(_0492_),
    .B1(net197),
    .B2(_0624_),
    .C1(_0627_),
    .X(_0628_));
 sky130_fd_sc_hd__nand2_1 _5094_ (.A(_0628_),
    .B(_0613_),
    .Y(_0629_));
 sky130_fd_sc_hd__o21ai_1 _5095_ (.A1(_0613_),
    .A2(_0623_),
    .B1(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__buf_8 _5096_ (.A(_0419_),
    .X(_0631_));
 sky130_fd_sc_hd__buf_8 _5097_ (.A(_0417_),
    .X(_0632_));
 sky130_fd_sc_hd__buf_8 _5098_ (.A(_0465_),
    .X(_0633_));
 sky130_fd_sc_hd__a21o_1 _5099_ (.A1(_0621_),
    .A2(_0632_),
    .B1(_0633_),
    .X(_0634_));
 sky130_fd_sc_hd__a221o_1 _5100_ (.A1(_0604_),
    .A2(_0611_),
    .B1(_0630_),
    .B2(_0631_),
    .C1(_0634_),
    .X(_0635_));
 sky130_fd_sc_hd__buf_6 _5101_ (.A(_0601_),
    .X(_0636_));
 sky130_fd_sc_hd__buf_8 _5102_ (.A(_0449_),
    .X(_0637_));
 sky130_fd_sc_hd__o22a_1 _5103_ (.A1(net87),
    .A2(_0454_),
    .B1(net25),
    .B2(_0456_),
    .X(_0638_));
 sky130_fd_sc_hd__o221a_4 _5104_ (.A1(net206),
    .A2(_0637_),
    .B1(net189),
    .B2(_0452_),
    .C1(_0638_),
    .X(_0639_));
 sky130_fd_sc_hd__inv_2 _5105_ (.A(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__nor2_1 _5106_ (.A(_0110_),
    .B(_0640_),
    .Y(_0641_));
 sky130_fd_sc_hd__a221o_1 _5107_ (.A1(_0574_),
    .A2(_0108_),
    .B1(_0572_),
    .B2(_0576_),
    .C1(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__or2_1 _5108_ (.A(_0463_),
    .B(_0642_),
    .X(_0643_));
 sky130_fd_sc_hd__or2_1 _5109_ (.A(_0461_),
    .B(_0574_),
    .X(_0644_));
 sky130_fd_sc_hd__buf_4 _5110_ (.A(_0484_),
    .X(_0645_));
 sky130_fd_sc_hd__buf_12 _5111_ (.A(_0467_),
    .X(_0646_));
 sky130_fd_sc_hd__o22a_1 _5112_ (.A1(net85),
    .A2(_0475_),
    .B1(net22),
    .B2(_0479_),
    .X(_0647_));
 sky130_fd_sc_hd__o221a_4 _5113_ (.A1(net184),
    .A2(_0646_),
    .B1(net187),
    .B2(_0472_),
    .C1(_0647_),
    .X(_0648_));
 sky130_fd_sc_hd__o22a_1 _5114_ (.A1(net87),
    .A2(_0475_),
    .B1(net25),
    .B2(_0479_),
    .X(_0649_));
 sky130_fd_sc_hd__o221a_4 _5115_ (.A1(net206),
    .A2(_0646_),
    .B1(net189),
    .B2(_0472_),
    .C1(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__buf_12 _5116_ (.A(_0196_),
    .X(_0651_));
 sky130_fd_sc_hd__buf_12 _5117_ (.A(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__clkinv_4 _5118_ (.A(_0200_),
    .Y(_0653_));
 sky130_fd_sc_hd__clkbuf_16 _5119_ (.A(_0653_),
    .X(_0654_));
 sky130_fd_sc_hd__o22a_1 _5120_ (.A1(net86),
    .A2(_0474_),
    .B1(net24),
    .B2(_0478_),
    .X(_0655_));
 sky130_fd_sc_hd__o221a_4 _5121_ (.A1(net195),
    .A2(_0468_),
    .B1(net188),
    .B2(_0471_),
    .C1(_0655_),
    .X(_0656_));
 sky130_fd_sc_hd__inv_2 _5122_ (.A(_0656_),
    .Y(_0657_));
 sky130_fd_sc_hd__nor2_1 _5123_ (.A(_0654_),
    .B(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__a221o_1 _5124_ (.A1(_0650_),
    .A2(_0652_),
    .B1(_0194_),
    .B2(_0648_),
    .C1(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__clkbuf_8 _5125_ (.A(_0487_),
    .X(_0660_));
 sky130_fd_sc_hd__a22o_1 _5126_ (.A1(_0645_),
    .A2(_0648_),
    .B1(_0659_),
    .B2(_0660_),
    .X(_0661_));
 sky130_fd_sc_hd__a41o_2 _5127_ (.A1(_0635_),
    .A2(_0636_),
    .A3(_0643_),
    .A4(_0644_),
    .B1(_0661_),
    .X(net586));
 sky130_fd_sc_hd__inv_2 _5128_ (.A(_0447_),
    .Y(_0662_));
 sky130_fd_sc_hd__buf_8 _5129_ (.A(_4149_),
    .X(_0663_));
 sky130_fd_sc_hd__buf_8 _5130_ (.A(_4147_),
    .X(_0664_));
 sky130_fd_sc_hd__a22o_1 _5131_ (.A1(_0663_),
    .A2(net195),
    .B1(_0664_),
    .B2(net188),
    .X(_0665_));
 sky130_fd_sc_hd__a221oi_2 _5132_ (.A1(net24),
    .A2(_0436_),
    .B1(net86),
    .B2(_0433_),
    .C1(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__inv_2 _5133_ (.A(_0465_),
    .Y(_0667_));
 sky130_fd_sc_hd__buf_4 _5134_ (.A(_0667_),
    .X(_0668_));
 sky130_fd_sc_hd__o221ai_1 _5135_ (.A1(_0604_),
    .A2(_0617_),
    .B1(_0662_),
    .B2(net730),
    .C1(_0668_),
    .Y(_0669_));
 sky130_fd_sc_hd__clkbuf_8 _5136_ (.A(_0601_),
    .X(_0670_));
 sky130_fd_sc_hd__o21a_1 _5137_ (.A1(_0668_),
    .A2(_0576_),
    .B1(_0670_),
    .X(_0671_));
 sky130_fd_sc_hd__a22o_2 _5138_ (.A1(_0567_),
    .A2(_0656_),
    .B1(_0669_),
    .B2(_0671_),
    .X(net587));
 sky130_fd_sc_hd__inv_2 _5139_ (.A(net206),
    .Y(_0672_));
 sky130_fd_sc_hd__inv_2 _5140_ (.A(net189),
    .Y(_0673_));
 sky130_fd_sc_hd__a22oi_1 _5141_ (.A1(_0432_),
    .A2(net87),
    .B1(_0435_),
    .B2(net25),
    .Y(_0674_));
 sky130_fd_sc_hd__o221a_4 _5142_ (.A1(_0672_),
    .A2(_0426_),
    .B1(_0673_),
    .B2(_0431_),
    .C1(_0674_),
    .X(_0675_));
 sky130_fd_sc_hd__inv_2 _5143_ (.A(_0675_),
    .Y(_0676_));
 sky130_fd_sc_hd__clkbuf_8 _5144_ (.A(_0441_),
    .X(_0677_));
 sky130_fd_sc_hd__clkbuf_16 _5145_ (.A(_4223_),
    .X(_0678_));
 sky130_fd_sc_hd__nor2_1 _5146_ (.A(_0678_),
    .B(_0675_),
    .Y(_0679_));
 sky130_fd_sc_hd__a22o_1 _5147_ (.A1(_0676_),
    .A2(_0677_),
    .B1(_0679_),
    .B2(_0589_),
    .X(_0680_));
 sky130_fd_sc_hd__nand2_1 _5148_ (.A(_0680_),
    .B(_0604_),
    .Y(_0681_));
 sky130_fd_sc_hd__clkbuf_8 _5149_ (.A(_0667_),
    .X(_0682_));
 sky130_fd_sc_hd__inv_2 _5150_ (.A(_0619_),
    .Y(_0683_));
 sky130_fd_sc_hd__nand2_1 _5151_ (.A(_0683_),
    .B(_0422_),
    .Y(_0684_));
 sky130_fd_sc_hd__o21ai_1 _5152_ (.A1(_0682_),
    .A2(_0639_),
    .B1(_0601_),
    .Y(_0685_));
 sky130_fd_sc_hd__a31o_1 _5153_ (.A1(_0681_),
    .A2(_0682_),
    .A3(_0684_),
    .B1(_0685_),
    .X(_0686_));
 sky130_fd_sc_hd__a21bo_1 _5154_ (.A1(_0567_),
    .A2(_0650_),
    .B1_N(_0686_),
    .X(net588));
 sky130_fd_sc_hd__o22a_1 _5155_ (.A1(net88),
    .A2(_0186_),
    .B1(net26),
    .B2(_0477_),
    .X(_0687_));
 sky130_fd_sc_hd__o221a_4 _5156_ (.A1(net217),
    .A2(_0467_),
    .B1(net190),
    .B2(_0185_),
    .C1(_0687_),
    .X(_0688_));
 sky130_fd_sc_hd__inv_2 _5157_ (.A(_0192_),
    .Y(_0689_));
 sky130_fd_sc_hd__nand2_1 _5158_ (.A(_0688_),
    .B(_0689_),
    .Y(_0690_));
 sky130_fd_sc_hd__nand2_1 _5159_ (.A(_0688_),
    .B(_0645_),
    .Y(_0691_));
 sky130_fd_sc_hd__a22o_1 _5160_ (.A1(_0663_),
    .A2(net217),
    .B1(_0664_),
    .B2(net190),
    .X(_0692_));
 sky130_fd_sc_hd__a221o_4 _5161_ (.A1(net26),
    .A2(_0435_),
    .B1(net88),
    .B2(_0432_),
    .C1(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__buf_8 _5162_ (.A(_4186_),
    .X(_0694_));
 sky130_fd_sc_hd__a22o_1 _5163_ (.A1(_0694_),
    .A2(_0676_),
    .B1(_0693_),
    .B2(_0523_),
    .X(_0695_));
 sky130_fd_sc_hd__a22o_1 _5164_ (.A1(_0663_),
    .A2(net228),
    .B1(_0664_),
    .B2(net191),
    .X(_0696_));
 sky130_fd_sc_hd__a221oi_2 _5165_ (.A1(net90),
    .A2(_0432_),
    .B1(net27),
    .B2(_0435_),
    .C1(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__inv_2 _5166_ (.A(_0697_),
    .Y(_0698_));
 sky130_fd_sc_hd__a22o_1 _5167_ (.A1(_0663_),
    .A2(net12),
    .B1(_4147_),
    .B2(net192),
    .X(_0699_));
 sky130_fd_sc_hd__a221oi_4 _5168_ (.A1(net28),
    .A2(_0435_),
    .B1(net91),
    .B2(_0432_),
    .C1(_0699_),
    .Y(_0700_));
 sky130_fd_sc_hd__inv_2 _5169_ (.A(_0700_),
    .Y(_0701_));
 sky130_fd_sc_hd__a22o_1 _5170_ (.A1(_0698_),
    .A2(_0694_),
    .B1(_0523_),
    .B2(_0701_),
    .X(_0702_));
 sky130_fd_sc_hd__nor2_8 _5171_ (.A(_4204_),
    .B(_0590_),
    .Y(_0703_));
 sky130_fd_sc_hd__buf_6 _5172_ (.A(_0703_),
    .X(_0704_));
 sky130_fd_sc_hd__mux2_1 _5173_ (.A0(_0695_),
    .A1(_0702_),
    .S(_0704_),
    .X(_0705_));
 sky130_fd_sc_hd__buf_6 _5174_ (.A(_0443_),
    .X(_0706_));
 sky130_fd_sc_hd__a22o_1 _5175_ (.A1(_0677_),
    .A2(_0693_),
    .B1(_0705_),
    .B2(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__nand2_1 _5176_ (.A(_0707_),
    .B(_0604_),
    .Y(_0708_));
 sky130_fd_sc_hd__o22a_1 _5177_ (.A1(net90),
    .A2(_0411_),
    .B1(net27),
    .B2(_0413_),
    .X(_0709_));
 sky130_fd_sc_hd__o221a_4 _5178_ (.A1(net228),
    .A2(_0492_),
    .B1(net191),
    .B2(_0409_),
    .C1(_0709_),
    .X(_0710_));
 sky130_fd_sc_hd__o22a_1 _5179_ (.A1(net91),
    .A2(_0625_),
    .B1(net28),
    .B2(_0626_),
    .X(_0711_));
 sky130_fd_sc_hd__o221a_4 _5180_ (.A1(net12),
    .A2(_0408_),
    .B1(net192),
    .B2(_0624_),
    .C1(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__a22o_1 _5181_ (.A1(_0710_),
    .A2(_0613_),
    .B1(_0558_),
    .B2(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__o22a_1 _5182_ (.A1(net88),
    .A2(_0411_),
    .B1(net26),
    .B2(_0413_),
    .X(_0714_));
 sky130_fd_sc_hd__o221a_4 _5183_ (.A1(net217),
    .A2(_0492_),
    .B1(net190),
    .B2(_0409_),
    .C1(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__a22o_1 _5184_ (.A1(_0683_),
    .A2(_0613_),
    .B1(_0715_),
    .B2(_0558_),
    .X(_0716_));
 sky130_fd_sc_hd__nor2_4 _5185_ (.A(_4268_),
    .B(_4278_),
    .Y(_0717_));
 sky130_fd_sc_hd__inv_6 _5186_ (.A(_0717_),
    .Y(_0718_));
 sky130_fd_sc_hd__buf_8 _5187_ (.A(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__mux2_2 _5188_ (.A0(_0713_),
    .A1(_0716_),
    .S(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__nand2_1 _5189_ (.A(_0720_),
    .B(_0631_),
    .Y(_0721_));
 sky130_fd_sc_hd__nand2_1 _5190_ (.A(_0715_),
    .B(_0632_),
    .Y(_0722_));
 sky130_fd_sc_hd__buf_8 _5191_ (.A(_0365_),
    .X(_0723_));
 sky130_fd_sc_hd__clkbuf_8 _5192_ (.A(_0123_),
    .X(_0724_));
 sky130_fd_sc_hd__clkbuf_8 _5193_ (.A(_0122_),
    .X(_0725_));
 sky130_fd_sc_hd__o22a_1 _5194_ (.A1(net88),
    .A2(_0724_),
    .B1(net26),
    .B2(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__o221a_4 _5195_ (.A1(net217),
    .A2(_0637_),
    .B1(net190),
    .B2(_0723_),
    .C1(_0726_),
    .X(_0727_));
 sky130_fd_sc_hd__inv_2 _5196_ (.A(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__buf_8 _5197_ (.A(_0111_),
    .X(_0729_));
 sky130_fd_sc_hd__buf_6 _5198_ (.A(_0088_),
    .X(_0730_));
 sky130_fd_sc_hd__a22o_1 _5199_ (.A1(_0639_),
    .A2(_0729_),
    .B1(_0730_),
    .B2(_0727_),
    .X(_0731_));
 sky130_fd_sc_hd__inv_2 _5200_ (.A(_0731_),
    .Y(_0732_));
 sky130_fd_sc_hd__a221o_1 _5201_ (.A1(_0460_),
    .A2(_0728_),
    .B1(_0732_),
    .B2(_0462_),
    .C1(_0489_),
    .X(_0733_));
 sky130_fd_sc_hd__a41o_1 _5202_ (.A1(_0708_),
    .A2(_0682_),
    .A3(_0721_),
    .A4(_0722_),
    .B1(_0733_),
    .X(_0734_));
 sky130_fd_sc_hd__o211ai_4 _5203_ (.A1(_0488_),
    .A2(_0690_),
    .B1(_0691_),
    .C1(_0734_),
    .Y(net589));
 sky130_fd_sc_hd__o22a_1 _5204_ (.A1(net90),
    .A2(_0186_),
    .B1(net27),
    .B2(_0189_),
    .X(_0735_));
 sky130_fd_sc_hd__o221a_4 _5205_ (.A1(net228),
    .A2(_0182_),
    .B1(net191),
    .B2(_0185_),
    .C1(_0735_),
    .X(_0736_));
 sky130_fd_sc_hd__a22o_1 _5206_ (.A1(_0710_),
    .A2(_0422_),
    .B1(_0698_),
    .B2(_0447_),
    .X(_0737_));
 sky130_fd_sc_hd__o22a_1 _5207_ (.A1(net90),
    .A2(_0724_),
    .B1(net27),
    .B2(_0725_),
    .X(_0738_));
 sky130_fd_sc_hd__o221a_4 _5208_ (.A1(net228),
    .A2(_0637_),
    .B1(net191),
    .B2(_0723_),
    .C1(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_1 _5209_ (.A0(_0737_),
    .A1(_0739_),
    .S(_0633_),
    .X(_0740_));
 sky130_fd_sc_hd__buf_12 _5210_ (.A(_0192_),
    .X(_0741_));
 sky130_fd_sc_hd__inv_2 _5211_ (.A(_0736_),
    .Y(_0742_));
 sky130_fd_sc_hd__nor2_1 _5212_ (.A(_0741_),
    .B(_0742_),
    .Y(_0743_));
 sky130_fd_sc_hd__and3_2 _5213_ (.A(_0743_),
    .B(_0209_),
    .C(_0194_),
    .X(_0744_));
 sky130_fd_sc_hd__a221o_1 _5214_ (.A1(_0645_),
    .A2(_0736_),
    .B1(_0740_),
    .B2(_0636_),
    .C1(_0744_),
    .X(net591));
 sky130_fd_sc_hd__o22a_1 _5215_ (.A1(net91),
    .A2(_0474_),
    .B1(net28),
    .B2(_0478_),
    .X(_0745_));
 sky130_fd_sc_hd__o221a_4 _5216_ (.A1(net12),
    .A2(_0468_),
    .B1(net192),
    .B2(_0471_),
    .C1(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__a22o_1 _5217_ (.A1(_0677_),
    .A2(_0701_),
    .B1(_0702_),
    .B2(_0706_),
    .X(_0747_));
 sky130_fd_sc_hd__inv_2 _5218_ (.A(_0712_),
    .Y(_0748_));
 sky130_fd_sc_hd__nor2_1 _5219_ (.A(_0604_),
    .B(_0748_),
    .Y(_0749_));
 sky130_fd_sc_hd__a211o_1 _5220_ (.A1(_0747_),
    .A2(_0604_),
    .B1(_0535_),
    .C1(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__o22a_1 _5221_ (.A1(net91),
    .A2(_0454_),
    .B1(net28),
    .B2(_0725_),
    .X(_0751_));
 sky130_fd_sc_hd__o221a_4 _5222_ (.A1(net12),
    .A2(_0637_),
    .B1(net192),
    .B2(_0723_),
    .C1(_0751_),
    .X(_0752_));
 sky130_fd_sc_hd__o22a_1 _5223_ (.A1(net92),
    .A2(_0724_),
    .B1(net29),
    .B2(_0725_),
    .X(_0753_));
 sky130_fd_sc_hd__o221a_4 _5224_ (.A1(net193),
    .A2(_0723_),
    .B1(net23),
    .B2(_0450_),
    .C1(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__o22a_1 _5225_ (.A1(net93),
    .A2(_0454_),
    .B1(net30),
    .B2(_0456_),
    .X(_0755_));
 sky130_fd_sc_hd__o221a_4 _5226_ (.A1(net34),
    .A2(_0450_),
    .B1(net194),
    .B2(_0452_),
    .C1(_0755_),
    .X(_0756_));
 sky130_fd_sc_hd__a22o_1 _5227_ (.A1(_0754_),
    .A2(_0729_),
    .B1(_0730_),
    .B2(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__a22o_1 _5228_ (.A1(_0739_),
    .A2(_0729_),
    .B1(_0730_),
    .B2(_0752_),
    .X(_0758_));
 sky130_fd_sc_hd__clkbuf_16 _5229_ (.A(_0105_),
    .X(_0759_));
 sky130_fd_sc_hd__nor2_2 _5230_ (.A(_0759_),
    .B(_0108_),
    .Y(_0760_));
 sky130_fd_sc_hd__inv_6 _5231_ (.A(_0760_),
    .Y(_0761_));
 sky130_fd_sc_hd__mux2_1 _5232_ (.A0(_0757_),
    .A1(_0758_),
    .S(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__o221a_1 _5233_ (.A1(_0461_),
    .A2(_0752_),
    .B1(_0463_),
    .B2(_0762_),
    .C1(_0670_),
    .X(_0763_));
 sky130_fd_sc_hd__a22o_2 _5234_ (.A1(_0567_),
    .A2(_0746_),
    .B1(_0750_),
    .B2(_0763_),
    .X(net592));
 sky130_fd_sc_hd__o22a_1 _5235_ (.A1(net92),
    .A2(_0186_),
    .B1(net29),
    .B2(_0477_),
    .X(_0764_));
 sky130_fd_sc_hd__o221a_4 _5236_ (.A1(net193),
    .A2(_0185_),
    .B1(net23),
    .B2(_0467_),
    .C1(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__clkbuf_16 _5237_ (.A(_0200_),
    .X(_0766_));
 sky130_fd_sc_hd__clkbuf_16 _5238_ (.A(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__and2_1 _5239_ (.A(_0765_),
    .B(_0689_),
    .X(_0768_));
 sky130_fd_sc_hd__clkbuf_8 _5240_ (.A(_0198_),
    .X(_0769_));
 sky130_fd_sc_hd__a22o_1 _5241_ (.A1(_0767_),
    .A2(_0746_),
    .B1(_0768_),
    .B2(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__clkbuf_8 _5242_ (.A(_0730_),
    .X(_0771_));
 sky130_fd_sc_hd__o22a_1 _5243_ (.A1(net94),
    .A2(_0724_),
    .B1(net31),
    .B2(_0725_),
    .X(_0772_));
 sky130_fd_sc_hd__o221a_4 _5244_ (.A1(net45),
    .A2(_0637_),
    .B1(net196),
    .B2(_0723_),
    .C1(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__a22o_1 _5245_ (.A1(_0756_),
    .A2(_0572_),
    .B1(_0771_),
    .B2(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__a22o_1 _5246_ (.A1(_0752_),
    .A2(_0729_),
    .B1(_0771_),
    .B2(_0754_),
    .X(_0775_));
 sky130_fd_sc_hd__mux2_1 _5247_ (.A0(_0774_),
    .A1(_0775_),
    .S(_0761_),
    .X(_0776_));
 sky130_fd_sc_hd__inv_2 _5248_ (.A(_0754_),
    .Y(_0777_));
 sky130_fd_sc_hd__nand2_1 _5249_ (.A(_0777_),
    .B(_0460_),
    .Y(_0778_));
 sky130_fd_sc_hd__o22a_1 _5250_ (.A1(net92),
    .A2(_0412_),
    .B1(net29),
    .B2(_0626_),
    .X(_0779_));
 sky130_fd_sc_hd__o221a_4 _5251_ (.A1(net193),
    .A2(_0624_),
    .B1(net23),
    .B2(_0408_),
    .C1(_0779_),
    .X(_0780_));
 sky130_fd_sc_hd__buf_8 _5252_ (.A(_0717_),
    .X(_0781_));
 sky130_fd_sc_hd__a22o_1 _5253_ (.A1(_0712_),
    .A2(_0612_),
    .B1(_0557_),
    .B2(_0780_),
    .X(_0782_));
 sky130_fd_sc_hd__o22a_1 _5254_ (.A1(net94),
    .A2(_0625_),
    .B1(net31),
    .B2(_0413_),
    .X(_0783_));
 sky130_fd_sc_hd__o221a_4 _5255_ (.A1(net45),
    .A2(_0492_),
    .B1(net196),
    .B2(_0624_),
    .C1(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__buf_8 _5256_ (.A(_4272_),
    .X(_0785_));
 sky130_fd_sc_hd__nand2_1 _5257_ (.A(_0784_),
    .B(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__o22a_1 _5258_ (.A1(net93),
    .A2(_0625_),
    .B1(net30),
    .B2(_0626_),
    .X(_0787_));
 sky130_fd_sc_hd__o221a_4 _5259_ (.A1(net34),
    .A2(_0492_),
    .B1(net194),
    .B2(_0624_),
    .C1(_0787_),
    .X(_0788_));
 sky130_fd_sc_hd__nand2_1 _5260_ (.A(_0788_),
    .B(_0785_),
    .Y(_0789_));
 sky130_fd_sc_hd__mux2_1 _5261_ (.A0(_0786_),
    .A1(_0789_),
    .S(_4253_),
    .X(_0790_));
 sky130_fd_sc_hd__nand2_1 _5262_ (.A(_0790_),
    .B(_0781_),
    .Y(_0791_));
 sky130_fd_sc_hd__o21ai_1 _5263_ (.A1(_0781_),
    .A2(_0782_),
    .B1(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__inv_2 _5264_ (.A(_0792_),
    .Y(_0793_));
 sky130_fd_sc_hd__inv_2 _5265_ (.A(net193),
    .Y(_0794_));
 sky130_fd_sc_hd__inv_2 _5266_ (.A(net23),
    .Y(_0795_));
 sky130_fd_sc_hd__a22oi_1 _5267_ (.A1(_0432_),
    .A2(net92),
    .B1(_0435_),
    .B2(net29),
    .Y(_0796_));
 sky130_fd_sc_hd__o221a_4 _5268_ (.A1(_0794_),
    .A2(_0430_),
    .B1(_0795_),
    .B2(_0425_),
    .C1(_0796_),
    .X(_0797_));
 sky130_fd_sc_hd__o21ai_1 _5269_ (.A1(_0591_),
    .A2(_0797_),
    .B1(_0525_),
    .Y(_0798_));
 sky130_fd_sc_hd__buf_8 _5270_ (.A(_4114_),
    .X(_0799_));
 sky130_fd_sc_hd__buf_8 _5271_ (.A(_0799_),
    .X(_0800_));
 sky130_fd_sc_hd__inv_2 _5272_ (.A(net45),
    .Y(_0801_));
 sky130_fd_sc_hd__inv_2 _5273_ (.A(net196),
    .Y(_0802_));
 sky130_fd_sc_hd__buf_6 _5274_ (.A(_0263_),
    .X(_0803_));
 sky130_fd_sc_hd__clkbuf_8 _5275_ (.A(_0434_),
    .X(_0804_));
 sky130_fd_sc_hd__a22oi_2 _5276_ (.A1(_0803_),
    .A2(net94),
    .B1(_0804_),
    .B2(net31),
    .Y(_0805_));
 sky130_fd_sc_hd__o221a_2 _5277_ (.A1(_0801_),
    .A2(_0424_),
    .B1(_0802_),
    .B2(_0429_),
    .C1(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__a22o_1 _5278_ (.A1(_0663_),
    .A2(net34),
    .B1(_0664_),
    .B2(net194),
    .X(_0807_));
 sky130_fd_sc_hd__a221o_4 _5279_ (.A1(net30),
    .A2(_0435_),
    .B1(net93),
    .B2(_0432_),
    .C1(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__nand2_1 _5280_ (.A(_0808_),
    .B(_0694_),
    .Y(_0809_));
 sky130_fd_sc_hd__o21ai_1 _5281_ (.A1(_0800_),
    .A2(_0806_),
    .B1(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__nand2_1 _5282_ (.A(_0701_),
    .B(_0694_),
    .Y(_0811_));
 sky130_fd_sc_hd__o21ai_1 _5283_ (.A1(_0800_),
    .A2(_0797_),
    .B1(_0811_),
    .Y(_0812_));
 sky130_fd_sc_hd__inv_4 _5284_ (.A(_0703_),
    .Y(_0813_));
 sky130_fd_sc_hd__mux2_1 _5285_ (.A0(_0810_),
    .A1(_0812_),
    .S(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__a22o_1 _5286_ (.A1(_0550_),
    .A2(_0798_),
    .B1(_0814_),
    .B2(_0706_),
    .X(_0815_));
 sky130_fd_sc_hd__o221ai_4 _5287_ (.A1(_0418_),
    .A2(_0780_),
    .B1(_0420_),
    .B2(_0793_),
    .C1(_0815_),
    .Y(_0816_));
 sky130_fd_sc_hd__nand2_1 _5288_ (.A(_0816_),
    .B(_0682_),
    .Y(_0817_));
 sky130_fd_sc_hd__o2111a_1 _5289_ (.A1(_0463_),
    .A2(_0776_),
    .B1(_0601_),
    .C1(_0778_),
    .D1(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__a221o_2 _5290_ (.A1(_0645_),
    .A2(_0765_),
    .B1(_0660_),
    .B2(_0770_),
    .C1(_0818_),
    .X(net593));
 sky130_fd_sc_hd__inv_2 _5291_ (.A(_0797_),
    .Y(_0819_));
 sky130_fd_sc_hd__nand2_1 _5292_ (.A(_0819_),
    .B(_0694_),
    .Y(_0820_));
 sky130_fd_sc_hd__a21bo_1 _5293_ (.A1(_0808_),
    .A2(_0523_),
    .B1_N(_0820_),
    .X(_0821_));
 sky130_fd_sc_hd__inv_2 _5294_ (.A(net56),
    .Y(_0822_));
 sky130_fd_sc_hd__inv_2 _5295_ (.A(net197),
    .Y(_0823_));
 sky130_fd_sc_hd__a22oi_1 _5296_ (.A1(_0803_),
    .A2(net95),
    .B1(_0435_),
    .B2(net32),
    .Y(_0824_));
 sky130_fd_sc_hd__o221a_2 _5297_ (.A1(_0822_),
    .A2(_0425_),
    .B1(_0823_),
    .B2(_0430_),
    .C1(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__inv_2 _5298_ (.A(_0806_),
    .Y(_0826_));
 sky130_fd_sc_hd__nand2_1 _5299_ (.A(_0826_),
    .B(_0694_),
    .Y(_0827_));
 sky130_fd_sc_hd__o21ai_1 _5300_ (.A1(_0800_),
    .A2(_0825_),
    .B1(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__or2_1 _5301_ (.A(_0813_),
    .B(_0828_),
    .X(_0829_));
 sky130_fd_sc_hd__o21ai_1 _5302_ (.A1(_0704_),
    .A2(_0821_),
    .B1(_0829_),
    .Y(_0830_));
 sky130_fd_sc_hd__inv_2 _5303_ (.A(_0830_),
    .Y(_0831_));
 sky130_fd_sc_hd__a22o_1 _5304_ (.A1(_0677_),
    .A2(_0808_),
    .B1(_0831_),
    .B2(_0706_),
    .X(_0832_));
 sky130_fd_sc_hd__buf_8 _5305_ (.A(_0781_),
    .X(_0833_));
 sky130_fd_sc_hd__a22o_1 _5306_ (.A1(_0780_),
    .A2(_0613_),
    .B1(_0558_),
    .B2(_0788_),
    .X(_0834_));
 sky130_fd_sc_hd__a22o_1 _5307_ (.A1(_0784_),
    .A2(_0612_),
    .B1(_0557_),
    .B2(_0628_),
    .X(_0835_));
 sky130_fd_sc_hd__or2_1 _5308_ (.A(_0718_),
    .B(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__o21ai_1 _5309_ (.A1(_0833_),
    .A2(_0834_),
    .B1(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__inv_2 _5310_ (.A(_0837_),
    .Y(_0838_));
 sky130_fd_sc_hd__a22o_1 _5311_ (.A1(_0632_),
    .A2(_0788_),
    .B1(_0838_),
    .B2(_0631_),
    .X(_0839_));
 sky130_fd_sc_hd__a211o_1 _5312_ (.A1(_0832_),
    .A2(_0604_),
    .B1(_0535_),
    .C1(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__clkbuf_8 _5313_ (.A(_0760_),
    .X(_0841_));
 sky130_fd_sc_hd__o22a_1 _5314_ (.A1(net95),
    .A2(_0724_),
    .B1(net32),
    .B2(_0725_),
    .X(_0842_));
 sky130_fd_sc_hd__o221a_4 _5315_ (.A1(net56),
    .A2(_0637_),
    .B1(net197),
    .B2(_0723_),
    .C1(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__buf_6 _5316_ (.A(_0152_),
    .X(_0844_));
 sky130_fd_sc_hd__nand2_1 _5317_ (.A(_0843_),
    .B(_0844_),
    .Y(_0845_));
 sky130_fd_sc_hd__nand2_1 _5318_ (.A(_0773_),
    .B(_0844_),
    .Y(_0846_));
 sky130_fd_sc_hd__mux2_1 _5319_ (.A0(_0845_),
    .A1(_0846_),
    .S(_0090_),
    .X(_0847_));
 sky130_fd_sc_hd__nand2_1 _5320_ (.A(_0847_),
    .B(_0841_),
    .Y(_0848_));
 sky130_fd_sc_hd__o21ai_2 _5321_ (.A1(_0841_),
    .A2(_0757_),
    .B1(_0848_),
    .Y(_0849_));
 sky130_fd_sc_hd__nand2_1 _5322_ (.A(_0849_),
    .B(_0462_),
    .Y(_0850_));
 sky130_fd_sc_hd__inv_2 _5323_ (.A(_0756_),
    .Y(_0851_));
 sky130_fd_sc_hd__nand2_1 _5324_ (.A(_0851_),
    .B(_0460_),
    .Y(_0852_));
 sky130_fd_sc_hd__o22a_1 _5325_ (.A1(net93),
    .A2(_0186_),
    .B1(net30),
    .B2(_0477_),
    .X(_0853_));
 sky130_fd_sc_hd__o221a_4 _5326_ (.A1(net34),
    .A2(_0467_),
    .B1(net194),
    .B2(_0185_),
    .C1(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__clkbuf_16 _5327_ (.A(_0195_),
    .X(_0855_));
 sky130_fd_sc_hd__nand2_1 _5328_ (.A(_0854_),
    .B(_0689_),
    .Y(_0856_));
 sky130_fd_sc_hd__nand2_1 _5329_ (.A(_0768_),
    .B(_0855_),
    .Y(_0857_));
 sky130_fd_sc_hd__o21ai_2 _5330_ (.A1(_0855_),
    .A2(_0856_),
    .B1(_0857_),
    .Y(_0858_));
 sky130_fd_sc_hd__a22o_1 _5331_ (.A1(_0645_),
    .A2(_0854_),
    .B1(_0858_),
    .B2(_0660_),
    .X(_0859_));
 sky130_fd_sc_hd__a41o_2 _5332_ (.A1(_0840_),
    .A2(_0636_),
    .A3(_0850_),
    .A4(_0852_),
    .B1(_0859_),
    .X(net594));
 sky130_fd_sc_hd__nor2_1 _5333_ (.A(_0591_),
    .B(_0806_),
    .Y(_0860_));
 sky130_fd_sc_hd__o21ai_1 _5334_ (.A1(_0548_),
    .A2(_0860_),
    .B1(_0550_),
    .Y(_0861_));
 sky130_fd_sc_hd__buf_6 _5335_ (.A(_0813_),
    .X(_0862_));
 sky130_fd_sc_hd__inv_2 _5336_ (.A(_0825_),
    .Y(_0863_));
 sky130_fd_sc_hd__inv_2 _5337_ (.A(net67),
    .Y(_0864_));
 sky130_fd_sc_hd__inv_2 _5338_ (.A(net198),
    .Y(_0865_));
 sky130_fd_sc_hd__a22oi_2 _5339_ (.A1(_0263_),
    .A2(net96),
    .B1(_0434_),
    .B2(net33),
    .Y(_0866_));
 sky130_fd_sc_hd__o221a_2 _5340_ (.A1(_0864_),
    .A2(_0424_),
    .B1(_0865_),
    .B2(_0429_),
    .C1(_0866_),
    .X(_0867_));
 sky130_fd_sc_hd__nor2_1 _5341_ (.A(_4204_),
    .B(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__a22o_1 _5342_ (.A1(_0863_),
    .A2(_0694_),
    .B1(_0868_),
    .B2(_0522_),
    .X(_0869_));
 sky130_fd_sc_hd__or2_1 _5343_ (.A(_0704_),
    .B(_0810_),
    .X(_0870_));
 sky130_fd_sc_hd__o21ai_1 _5344_ (.A1(_0862_),
    .A2(_0869_),
    .B1(_0870_),
    .Y(_0871_));
 sky130_fd_sc_hd__inv_2 _5345_ (.A(_0871_),
    .Y(_0872_));
 sky130_fd_sc_hd__nand2_1 _5346_ (.A(_0872_),
    .B(_0706_),
    .Y(_0873_));
 sky130_fd_sc_hd__a2bb2o_1 _5347_ (.A1_N(_0604_),
    .A2_N(_0784_),
    .B1(_0861_),
    .B2(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__nand2_1 _5348_ (.A(_0874_),
    .B(_0668_),
    .Y(_0875_));
 sky130_fd_sc_hd__o22a_1 _5349_ (.A1(net96),
    .A2(_0724_),
    .B1(net33),
    .B2(_0725_),
    .X(_0876_));
 sky130_fd_sc_hd__o221a_4 _5350_ (.A1(net67),
    .A2(_0637_),
    .B1(net198),
    .B2(_0723_),
    .C1(_0876_),
    .X(_0877_));
 sky130_fd_sc_hd__a22o_1 _5351_ (.A1(_0877_),
    .A2(_0730_),
    .B1(_0729_),
    .B2(_0843_),
    .X(_0878_));
 sky130_fd_sc_hd__inv_2 _5352_ (.A(_0878_),
    .Y(_0879_));
 sky130_fd_sc_hd__nand2_2 _5353_ (.A(_0879_),
    .B(_0841_),
    .Y(_0880_));
 sky130_fd_sc_hd__o21ai_2 _5354_ (.A1(_0841_),
    .A2(_0774_),
    .B1(_0880_),
    .Y(_0881_));
 sky130_fd_sc_hd__nand2_1 _5355_ (.A(_0881_),
    .B(_0462_),
    .Y(_0882_));
 sky130_fd_sc_hd__or2_1 _5356_ (.A(_0461_),
    .B(_0773_),
    .X(_0883_));
 sky130_fd_sc_hd__o22a_1 _5357_ (.A1(net94),
    .A2(_0474_),
    .B1(net31),
    .B2(_0478_),
    .X(_0884_));
 sky130_fd_sc_hd__o221a_4 _5358_ (.A1(net45),
    .A2(_0468_),
    .B1(net196),
    .B2(_0471_),
    .C1(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__nor2_4 _5359_ (.A(_0192_),
    .B(_0194_),
    .Y(_0886_));
 sky130_fd_sc_hd__buf_6 _5360_ (.A(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__buf_8 _5361_ (.A(_0689_),
    .X(_0888_));
 sky130_fd_sc_hd__nand2_1 _5362_ (.A(_0885_),
    .B(_0888_),
    .Y(_0889_));
 sky130_fd_sc_hd__or2_1 _5363_ (.A(_0198_),
    .B(_0856_),
    .X(_0890_));
 sky130_fd_sc_hd__o21ai_1 _5364_ (.A1(_0855_),
    .A2(_0889_),
    .B1(_0890_),
    .Y(_0891_));
 sky130_fd_sc_hd__o22a_1 _5365_ (.A1(net96),
    .A2(_0186_),
    .B1(net33),
    .B2(_0477_),
    .X(_0892_));
 sky130_fd_sc_hd__o221a_4 _5366_ (.A1(net67),
    .A2(_0467_),
    .B1(net198),
    .B2(_0185_),
    .C1(_0892_),
    .X(_0893_));
 sky130_fd_sc_hd__nand2_1 _5367_ (.A(_0893_),
    .B(_0888_),
    .Y(_0894_));
 sky130_fd_sc_hd__o22a_1 _5368_ (.A1(net95),
    .A2(_0474_),
    .B1(net32),
    .B2(_0477_),
    .X(_0895_));
 sky130_fd_sc_hd__o221a_4 _5369_ (.A1(net56),
    .A2(_0467_),
    .B1(net197),
    .B2(_0471_),
    .C1(_0895_),
    .X(_0896_));
 sky130_fd_sc_hd__nand2_1 _5370_ (.A(_0896_),
    .B(_0888_),
    .Y(_0897_));
 sky130_fd_sc_hd__mux2_1 _5371_ (.A0(_0894_),
    .A1(_0897_),
    .S(_0855_),
    .X(_0898_));
 sky130_fd_sc_hd__nand2_1 _5372_ (.A(_0898_),
    .B(_0886_),
    .Y(_0899_));
 sky130_fd_sc_hd__o21ai_1 _5373_ (.A1(_0887_),
    .A2(_0891_),
    .B1(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__inv_2 _5374_ (.A(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__a22o_1 _5375_ (.A1(_0645_),
    .A2(_0885_),
    .B1(_0901_),
    .B2(_0660_),
    .X(_0902_));
 sky130_fd_sc_hd__a41o_2 _5376_ (.A1(_0875_),
    .A2(_0636_),
    .A3(_0882_),
    .A4(_0883_),
    .B1(_0902_),
    .X(net595));
 sky130_fd_sc_hd__o22a_1 _5377_ (.A1(net97),
    .A2(_0036_),
    .B1(net35),
    .B2(_4289_),
    .X(_0903_));
 sky130_fd_sc_hd__o221a_4 _5378_ (.A1(net78),
    .A2(_0407_),
    .B1(net199),
    .B2(_0409_),
    .C1(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__o22a_1 _5379_ (.A1(net96),
    .A2(_0412_),
    .B1(net33),
    .B2(_0414_),
    .X(_0905_));
 sky130_fd_sc_hd__o221a_2 _5380_ (.A1(net67),
    .A2(_0408_),
    .B1(net198),
    .B2(_0410_),
    .C1(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__a221o_1 _5381_ (.A1(_0904_),
    .A2(_0558_),
    .B1(_0906_),
    .B2(_0613_),
    .C1(_0718_),
    .X(_0907_));
 sky130_fd_sc_hd__o21ai_1 _5382_ (.A1(_0833_),
    .A2(_0835_),
    .B1(_0907_),
    .Y(_0908_));
 sky130_fd_sc_hd__inv_2 _5383_ (.A(_0908_),
    .Y(_0909_));
 sky130_fd_sc_hd__clkbuf_16 _5384_ (.A(_4204_),
    .X(_0910_));
 sky130_fd_sc_hd__inv_2 _5385_ (.A(net78),
    .Y(_0911_));
 sky130_fd_sc_hd__inv_2 _5386_ (.A(net199),
    .Y(_0912_));
 sky130_fd_sc_hd__a22oi_1 _5387_ (.A1(_0803_),
    .A2(net97),
    .B1(_0804_),
    .B2(net35),
    .Y(_0913_));
 sky130_fd_sc_hd__o221a_4 _5388_ (.A1(_0911_),
    .A2(_0424_),
    .B1(_0912_),
    .B2(_0430_),
    .C1(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__nor2_1 _5389_ (.A(_0910_),
    .B(_0914_),
    .Y(_0915_));
 sky130_fd_sc_hd__nand2_1 _5390_ (.A(_0868_),
    .B(_0799_),
    .Y(_0916_));
 sky130_fd_sc_hd__inv_2 _5391_ (.A(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__a211o_1 _5392_ (.A1(_0522_),
    .A2(_0915_),
    .B1(_0813_),
    .C1(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__o21ai_1 _5393_ (.A1(_0703_),
    .A2(_0828_),
    .B1(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__inv_2 _5394_ (.A(_0919_),
    .Y(_0920_));
 sky130_fd_sc_hd__a221o_1 _5395_ (.A1(_0677_),
    .A2(_0863_),
    .B1(_0920_),
    .B2(_0706_),
    .C1(_0422_),
    .X(_0921_));
 sky130_fd_sc_hd__o221a_1 _5396_ (.A1(_0418_),
    .A2(_0628_),
    .B1(_0420_),
    .B2(_0909_),
    .C1(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__or2_1 _5397_ (.A(_0535_),
    .B(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__o21a_1 _5398_ (.A1(_0668_),
    .A2(_0843_),
    .B1(_0670_),
    .X(_0924_));
 sky130_fd_sc_hd__a22o_1 _5399_ (.A1(_0567_),
    .A2(_0896_),
    .B1(_0923_),
    .B2(_0924_),
    .X(net596));
 sky130_fd_sc_hd__inv_2 _5400_ (.A(_0906_),
    .Y(_0925_));
 sky130_fd_sc_hd__inv_2 _5401_ (.A(net89),
    .Y(_0926_));
 sky130_fd_sc_hd__inv_2 _5402_ (.A(net200),
    .Y(_0927_));
 sky130_fd_sc_hd__a22oi_1 _5403_ (.A1(_0803_),
    .A2(net98),
    .B1(_0804_),
    .B2(net36),
    .Y(_0928_));
 sky130_fd_sc_hd__o221a_2 _5404_ (.A1(_0926_),
    .A2(_0424_),
    .B1(_0927_),
    .B2(_0429_),
    .C1(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__nor2_1 _5405_ (.A(_0910_),
    .B(_0929_),
    .Y(_0930_));
 sky130_fd_sc_hd__mux2_2 _5406_ (.A0(_0930_),
    .A1(_0915_),
    .S(_4114_),
    .X(_0931_));
 sky130_fd_sc_hd__mux2_1 _5407_ (.A0(_0869_),
    .A1(_0931_),
    .S(_0703_),
    .X(_0932_));
 sky130_fd_sc_hd__nand2_1 _5408_ (.A(_0932_),
    .B(_0706_),
    .Y(_0933_));
 sky130_fd_sc_hd__nor2_1 _5409_ (.A(_0591_),
    .B(_0867_),
    .Y(_0934_));
 sky130_fd_sc_hd__o21ai_1 _5410_ (.A1(_0548_),
    .A2(_0934_),
    .B1(_0550_),
    .Y(_0935_));
 sky130_fd_sc_hd__a22o_1 _5411_ (.A1(_0422_),
    .A2(_0925_),
    .B1(_0933_),
    .B2(_0935_),
    .X(_0936_));
 sky130_fd_sc_hd__nand2_1 _5412_ (.A(_0936_),
    .B(_0668_),
    .Y(_0937_));
 sky130_fd_sc_hd__o21a_1 _5413_ (.A1(_0668_),
    .A2(_0877_),
    .B1(_0670_),
    .X(_0938_));
 sky130_fd_sc_hd__a22o_1 _5414_ (.A1(_0567_),
    .A2(_0893_),
    .B1(_0937_),
    .B2(_0938_),
    .X(net597));
 sky130_fd_sc_hd__o22a_1 _5415_ (.A1(net97),
    .A2(_0475_),
    .B1(net35),
    .B2(_0479_),
    .X(_0939_));
 sky130_fd_sc_hd__o221a_4 _5416_ (.A1(net78),
    .A2(_0646_),
    .B1(net199),
    .B2(_0472_),
    .C1(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__o22a_1 _5417_ (.A1(net99),
    .A2(_0036_),
    .B1(net37),
    .B2(_4289_),
    .X(_0941_));
 sky130_fd_sc_hd__o221a_4 _5418_ (.A1(net100),
    .A2(_0407_),
    .B1(net201),
    .B2(_0038_),
    .C1(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__o22a_1 _5419_ (.A1(net98),
    .A2(_0036_),
    .B1(net36),
    .B2(_4289_),
    .X(_0943_));
 sky130_fd_sc_hd__o221a_4 _5420_ (.A1(net89),
    .A2(_0407_),
    .B1(net200),
    .B2(_0038_),
    .C1(_0943_),
    .X(_0944_));
 sky130_fd_sc_hd__a22o_1 _5421_ (.A1(_0942_),
    .A2(_0510_),
    .B1(_4265_),
    .B2(_0944_),
    .X(_0945_));
 sky130_fd_sc_hd__and3_1 _5422_ (.A(_0904_),
    .B(_0558_),
    .C(\arbiter.slave_sel[1][1] ),
    .X(_0946_));
 sky130_fd_sc_hd__a21o_1 _5423_ (.A1(_0945_),
    .A2(_0833_),
    .B1(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__inv_2 _5424_ (.A(_0914_),
    .Y(_0948_));
 sky130_fd_sc_hd__or3_1 _5425_ (.A(_0800_),
    .B(_4119_),
    .C(_0914_),
    .X(_0949_));
 sky130_fd_sc_hd__inv_2 _5426_ (.A(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__a22o_1 _5427_ (.A1(_0677_),
    .A2(_0948_),
    .B1(_0950_),
    .B2(_0589_),
    .X(_0951_));
 sky130_fd_sc_hd__a21o_1 _5428_ (.A1(_0904_),
    .A2(_0632_),
    .B1(_0633_),
    .X(_0952_));
 sky130_fd_sc_hd__a221o_2 _5429_ (.A1(_0631_),
    .A2(_0947_),
    .B1(_0951_),
    .B2(_0604_),
    .C1(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__o22a_1 _5430_ (.A1(net97),
    .A2(_0724_),
    .B1(net35),
    .B2(_0725_),
    .X(_0954_));
 sky130_fd_sc_hd__o221a_4 _5431_ (.A1(net78),
    .A2(_0637_),
    .B1(net199),
    .B2(_0723_),
    .C1(_0954_),
    .X(_0955_));
 sky130_fd_sc_hd__o21a_1 _5432_ (.A1(_0668_),
    .A2(_0955_),
    .B1(_0670_),
    .X(_0956_));
 sky130_fd_sc_hd__a22o_1 _5433_ (.A1(_0567_),
    .A2(_0940_),
    .B1(_0953_),
    .B2(_0956_),
    .X(net598));
 sky130_fd_sc_hd__inv_2 _5434_ (.A(_0929_),
    .Y(_0957_));
 sky130_fd_sc_hd__inv_2 _5435_ (.A(net202),
    .Y(_0958_));
 sky130_fd_sc_hd__inv_2 _5436_ (.A(net111),
    .Y(_0959_));
 sky130_fd_sc_hd__a22oi_1 _5437_ (.A1(_0263_),
    .A2(net101),
    .B1(_0804_),
    .B2(net38),
    .Y(_0960_));
 sky130_fd_sc_hd__o221a_2 _5438_ (.A1(_0958_),
    .A2(_0429_),
    .B1(_0959_),
    .B2(_0425_),
    .C1(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__nor2_1 _5439_ (.A(_0910_),
    .B(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__inv_2 _5440_ (.A(net100),
    .Y(_0963_));
 sky130_fd_sc_hd__inv_2 _5441_ (.A(net201),
    .Y(_0964_));
 sky130_fd_sc_hd__a22oi_1 _5442_ (.A1(_0803_),
    .A2(net99),
    .B1(_0804_),
    .B2(net37),
    .Y(_0965_));
 sky130_fd_sc_hd__o221a_2 _5443_ (.A1(_0963_),
    .A2(_0425_),
    .B1(_0964_),
    .B2(_0430_),
    .C1(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__nor2_1 _5444_ (.A(_0910_),
    .B(_0966_),
    .Y(_0967_));
 sky130_fd_sc_hd__mux2_1 _5445_ (.A0(_0962_),
    .A1(_0967_),
    .S(_0799_),
    .X(_0968_));
 sky130_fd_sc_hd__mux2_1 _5446_ (.A0(_0931_),
    .A1(_0968_),
    .S(_0703_),
    .X(_0969_));
 sky130_fd_sc_hd__a22o_1 _5447_ (.A1(_0441_),
    .A2(_0957_),
    .B1(_0969_),
    .B2(_0443_),
    .X(_0970_));
 sky130_fd_sc_hd__a22o_1 _5448_ (.A1(_0904_),
    .A2(_4265_),
    .B1(_0510_),
    .B2(_0944_),
    .X(_0971_));
 sky130_fd_sc_hd__o22a_1 _5449_ (.A1(net101),
    .A2(_0036_),
    .B1(net38),
    .B2(_4289_),
    .X(_0972_));
 sky130_fd_sc_hd__o221a_4 _5450_ (.A1(net202),
    .A2(_0038_),
    .B1(net111),
    .B2(_0407_),
    .C1(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__a22o_1 _5451_ (.A1(_0942_),
    .A2(_4265_),
    .B1(_0510_),
    .B2(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__mux2_1 _5452_ (.A0(_0971_),
    .A1(_0974_),
    .S(_0717_),
    .X(_0975_));
 sky130_fd_sc_hd__inv_2 _5453_ (.A(_0975_),
    .Y(_0976_));
 sky130_fd_sc_hd__nor2_1 _5454_ (.A(_0420_),
    .B(_0976_),
    .Y(_0977_));
 sky130_fd_sc_hd__a221o_1 _5455_ (.A1(_0417_),
    .A2(_0944_),
    .B1(_0970_),
    .B2(_0592_),
    .C1(_0977_),
    .X(_0978_));
 sky130_fd_sc_hd__o22a_1 _5456_ (.A1(net98),
    .A2(_0123_),
    .B1(net36),
    .B2(_0122_),
    .X(_0979_));
 sky130_fd_sc_hd__o221a_4 _5457_ (.A1(net89),
    .A2(_0449_),
    .B1(net200),
    .B2(_0365_),
    .C1(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__mux2_2 _5458_ (.A0(_0978_),
    .A1(_0980_),
    .S(_0465_),
    .X(_0981_));
 sky130_fd_sc_hd__o22a_1 _5459_ (.A1(net98),
    .A2(_0476_),
    .B1(net36),
    .B2(_0479_),
    .X(_0982_));
 sky130_fd_sc_hd__o221a_4 _5460_ (.A1(net89),
    .A2(_0470_),
    .B1(net200),
    .B2(_0472_),
    .C1(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__mux2_1 _5461_ (.A0(_0981_),
    .A1(_0983_),
    .S(_0490_),
    .X(_0984_));
 sky130_fd_sc_hd__buf_1 _5462_ (.A(_0984_),
    .X(net599));
 sky130_fd_sc_hd__o22a_1 _5463_ (.A1(net99),
    .A2(_0475_),
    .B1(net37),
    .B2(_0479_),
    .X(_0985_));
 sky130_fd_sc_hd__o221a_4 _5464_ (.A1(net100),
    .A2(_0469_),
    .B1(net201),
    .B2(_0472_),
    .C1(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__inv_2 _5465_ (.A(_0942_),
    .Y(_0987_));
 sky130_fd_sc_hd__inv_2 _5466_ (.A(_0945_),
    .Y(_0988_));
 sky130_fd_sc_hd__o22a_1 _5467_ (.A1(net102),
    .A2(_0036_),
    .B1(net39),
    .B2(_4289_),
    .X(_0989_));
 sky130_fd_sc_hd__o221a_4 _5468_ (.A1(net123),
    .A2(_0407_),
    .B1(net203),
    .B2(_0038_),
    .C1(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__a22o_1 _5469_ (.A1(_0973_),
    .A2(_4265_),
    .B1(_0510_),
    .B2(_0990_),
    .X(_0991_));
 sky130_fd_sc_hd__inv_2 _5470_ (.A(_0991_),
    .Y(_0992_));
 sky130_fd_sc_hd__mux2_2 _5471_ (.A0(_0988_),
    .A1(_0992_),
    .S(_0717_),
    .X(_0993_));
 sky130_fd_sc_hd__o22a_1 _5472_ (.A1(net107),
    .A2(_0625_),
    .B1(net44),
    .B2(_0626_),
    .X(_0994_));
 sky130_fd_sc_hd__o221a_4 _5473_ (.A1(net146),
    .A2(_0408_),
    .B1(net209),
    .B2(_0624_),
    .C1(_0994_),
    .X(_0995_));
 sky130_fd_sc_hd__o22a_1 _5474_ (.A1(net108),
    .A2(_0625_),
    .B1(net46),
    .B2(_0626_),
    .X(_0996_));
 sky130_fd_sc_hd__o221a_4 _5475_ (.A1(net147),
    .A2(_0492_),
    .B1(net210),
    .B2(_0624_),
    .C1(_0996_),
    .X(_0997_));
 sky130_fd_sc_hd__a22o_1 _5476_ (.A1(_0995_),
    .A2(_0612_),
    .B1(_0557_),
    .B2(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__o22a_1 _5477_ (.A1(net109),
    .A2(_0036_),
    .B1(net47),
    .B2(_4289_),
    .X(_0999_));
 sky130_fd_sc_hd__o221a_4 _5478_ (.A1(net211),
    .A2(_0038_),
    .B1(net148),
    .B2(_0407_),
    .C1(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__o22a_1 _5479_ (.A1(net110),
    .A2(_0036_),
    .B1(net48),
    .B2(_4289_),
    .X(_1001_));
 sky130_fd_sc_hd__o221a_2 _5480_ (.A1(net149),
    .A2(_0407_),
    .B1(net212),
    .B2(_0038_),
    .C1(_1001_),
    .X(_1002_));
 sky130_fd_sc_hd__a22o_1 _5481_ (.A1(_1000_),
    .A2(_4265_),
    .B1(_0510_),
    .B2(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__or2_1 _5482_ (.A(_0718_),
    .B(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__o21ai_4 _5483_ (.A1(_0781_),
    .A2(_0998_),
    .B1(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__mux2_1 _5484_ (.A0(_0993_),
    .A1(_1005_),
    .S(_0613_),
    .X(_1006_));
 sky130_fd_sc_hd__buf_8 _5485_ (.A(_4158_),
    .X(_1007_));
 sky130_fd_sc_hd__mux2_1 _5486_ (.A0(_0930_),
    .A1(_0967_),
    .S(_0523_),
    .X(_1008_));
 sky130_fd_sc_hd__nand2_1 _5487_ (.A(_1008_),
    .B(_0862_),
    .Y(_1009_));
 sky130_fd_sc_hd__o221a_1 _5488_ (.A1(_0591_),
    .A2(_0966_),
    .B1(_1007_),
    .B2(_1009_),
    .C1(_0592_),
    .X(_1010_));
 sky130_fd_sc_hd__a221o_2 _5489_ (.A1(_0632_),
    .A2(_0987_),
    .B1(_1006_),
    .B2(_0631_),
    .C1(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__nand2_1 _5490_ (.A(_1011_),
    .B(_0668_),
    .Y(_1012_));
 sky130_fd_sc_hd__o22a_1 _5491_ (.A1(net99),
    .A2(_0123_),
    .B1(net37),
    .B2(_0122_),
    .X(_1013_));
 sky130_fd_sc_hd__o221a_4 _5492_ (.A1(net100),
    .A2(_0449_),
    .B1(net201),
    .B2(_0365_),
    .C1(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__o21a_1 _5493_ (.A1(_0668_),
    .A2(_1014_),
    .B1(_0670_),
    .X(_1015_));
 sky130_fd_sc_hd__a22o_2 _5494_ (.A1(_0567_),
    .A2(_0986_),
    .B1(_1012_),
    .B2(_1015_),
    .X(net600));
 sky130_fd_sc_hd__o22a_1 _5495_ (.A1(net101),
    .A2(_0476_),
    .B1(net38),
    .B2(_0479_),
    .X(_1016_));
 sky130_fd_sc_hd__o221a_4 _5496_ (.A1(net202),
    .A2(_0473_),
    .B1(net111),
    .B2(_0470_),
    .C1(_1016_),
    .X(_1017_));
 sky130_fd_sc_hd__o22a_1 _5497_ (.A1(net101),
    .A2(_0123_),
    .B1(net38),
    .B2(_0122_),
    .X(_1018_));
 sky130_fd_sc_hd__o221a_4 _5498_ (.A1(net202),
    .A2(_0365_),
    .B1(net111),
    .B2(_0449_),
    .C1(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__o22a_1 _5499_ (.A1(net103),
    .A2(_0411_),
    .B1(net40),
    .B2(_0413_),
    .X(_1020_));
 sky130_fd_sc_hd__o221a_4 _5500_ (.A1(net134),
    .A2(_0492_),
    .B1(net204),
    .B2(_0409_),
    .C1(_1020_),
    .X(_1021_));
 sky130_fd_sc_hd__a22o_1 _5501_ (.A1(_0990_),
    .A2(_0612_),
    .B1(_0510_),
    .B2(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__mux2_1 _5502_ (.A0(_1022_),
    .A1(_0974_),
    .S(_0718_),
    .X(_1023_));
 sky130_fd_sc_hd__a221o_1 _5503_ (.A1(_0632_),
    .A2(_0973_),
    .B1(_1023_),
    .B2(_0631_),
    .C1(_0633_),
    .X(_1024_));
 sky130_fd_sc_hd__inv_2 _5504_ (.A(_0961_),
    .Y(_1025_));
 sky130_fd_sc_hd__inv_2 _5505_ (.A(net134),
    .Y(_1026_));
 sky130_fd_sc_hd__inv_2 _5506_ (.A(net204),
    .Y(_1027_));
 sky130_fd_sc_hd__a22oi_1 _5507_ (.A1(_0432_),
    .A2(net103),
    .B1(_0435_),
    .B2(net40),
    .Y(_1028_));
 sky130_fd_sc_hd__o221a_2 _5508_ (.A1(_1026_),
    .A2(_0425_),
    .B1(_1027_),
    .B2(_0430_),
    .C1(_1028_),
    .X(_1029_));
 sky130_fd_sc_hd__nor2_1 _5509_ (.A(_0538_),
    .B(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__inv_2 _5510_ (.A(net123),
    .Y(_1031_));
 sky130_fd_sc_hd__inv_2 _5511_ (.A(net203),
    .Y(_1032_));
 sky130_fd_sc_hd__a22oi_1 _5512_ (.A1(_0803_),
    .A2(net102),
    .B1(_0435_),
    .B2(net39),
    .Y(_1033_));
 sky130_fd_sc_hd__o221a_4 _5513_ (.A1(_1031_),
    .A2(_0425_),
    .B1(_1032_),
    .B2(_0430_),
    .C1(_1033_),
    .X(_1034_));
 sky130_fd_sc_hd__nor2_1 _5514_ (.A(_0538_),
    .B(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__mux2_1 _5515_ (.A0(_1030_),
    .A1(_1035_),
    .S(_0799_),
    .X(_1036_));
 sky130_fd_sc_hd__or2_1 _5516_ (.A(_0813_),
    .B(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__o21ai_1 _5517_ (.A1(_0704_),
    .A2(_0968_),
    .B1(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__inv_2 _5518_ (.A(net149),
    .Y(_1039_));
 sky130_fd_sc_hd__inv_2 _5519_ (.A(net212),
    .Y(_1040_));
 sky130_fd_sc_hd__a22oi_1 _5520_ (.A1(_0263_),
    .A2(net110),
    .B1(_0434_),
    .B2(net48),
    .Y(_1041_));
 sky130_fd_sc_hd__o221a_2 _5521_ (.A1(_1039_),
    .A2(_0424_),
    .B1(_1040_),
    .B2(_0429_),
    .C1(_1041_),
    .X(_1042_));
 sky130_fd_sc_hd__nor2_1 _5522_ (.A(_4204_),
    .B(_1042_),
    .Y(_1043_));
 sky130_fd_sc_hd__nand2_1 _5523_ (.A(_1043_),
    .B(_0799_),
    .Y(_1044_));
 sky130_fd_sc_hd__o21ai_1 _5524_ (.A1(_0800_),
    .A2(_1038_),
    .B1(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__a22o_1 _5525_ (.A1(_0677_),
    .A2(_1025_),
    .B1(_1045_),
    .B2(_0706_),
    .X(_1046_));
 sky130_fd_sc_hd__and2_1 _5526_ (.A(_1046_),
    .B(_0604_),
    .X(_1047_));
 sky130_fd_sc_hd__o221a_1 _5527_ (.A1(_0682_),
    .A2(_1019_),
    .B1(_1024_),
    .B2(_1047_),
    .C1(_0636_),
    .X(_1048_));
 sky130_fd_sc_hd__a21o_2 _5528_ (.A1(_0567_),
    .A2(_1017_),
    .B1(_1048_),
    .X(net602));
 sky130_fd_sc_hd__o22a_1 _5529_ (.A1(net102),
    .A2(_0476_),
    .B1(net39),
    .B2(_0480_),
    .X(_1049_));
 sky130_fd_sc_hd__o221a_4 _5530_ (.A1(net123),
    .A2(_0470_),
    .B1(net203),
    .B2(_0473_),
    .C1(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__o22a_1 _5531_ (.A1(net104),
    .A2(_0625_),
    .B1(net41),
    .B2(_0626_),
    .X(_1051_));
 sky130_fd_sc_hd__o221a_4 _5532_ (.A1(net143),
    .A2(_0408_),
    .B1(net205),
    .B2(_0624_),
    .C1(_1051_),
    .X(_1052_));
 sky130_fd_sc_hd__a22o_1 _5533_ (.A1(_1021_),
    .A2(_0612_),
    .B1(_0557_),
    .B2(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__inv_2 _5534_ (.A(_1053_),
    .Y(_1054_));
 sky130_fd_sc_hd__mux2_2 _5535_ (.A0(_1054_),
    .A1(_0992_),
    .S(_0719_),
    .X(_1055_));
 sky130_fd_sc_hd__o2bb2a_1 _5536_ (.A1_N(_0631_),
    .A2_N(_1055_),
    .B1(_0418_),
    .B2(_0990_),
    .X(_1056_));
 sky130_fd_sc_hd__nand2_1 _5537_ (.A(_0962_),
    .B(_0799_),
    .Y(_1057_));
 sky130_fd_sc_hd__inv_2 _5538_ (.A(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__a21o_1 _5539_ (.A1(_0523_),
    .A2(_1035_),
    .B1(_1058_),
    .X(_1059_));
 sky130_fd_sc_hd__o21ai_1 _5540_ (.A1(_0591_),
    .A2(_1034_),
    .B1(_0604_),
    .Y(_1060_));
 sky130_fd_sc_hd__a31o_1 _5541_ (.A1(_1059_),
    .A2(_0589_),
    .A3(_0862_),
    .B1(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__a21o_1 _5542_ (.A1(_1056_),
    .A2(_1061_),
    .B1(_0535_),
    .X(_1062_));
 sky130_fd_sc_hd__o22a_1 _5543_ (.A1(net102),
    .A2(_0123_),
    .B1(net39),
    .B2(_0122_),
    .X(_1063_));
 sky130_fd_sc_hd__o221a_4 _5544_ (.A1(net123),
    .A2(_0449_),
    .B1(net203),
    .B2(_0365_),
    .C1(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__o21a_1 _5545_ (.A1(_0668_),
    .A2(_1064_),
    .B1(_0670_),
    .X(_1065_));
 sky130_fd_sc_hd__a22o_2 _5546_ (.A1(_0567_),
    .A2(_1050_),
    .B1(_1062_),
    .B2(_1065_),
    .X(net603));
 sky130_fd_sc_hd__o22a_1 _5547_ (.A1(net103),
    .A2(_0476_),
    .B1(net40),
    .B2(_0480_),
    .X(_1066_));
 sky130_fd_sc_hd__o221a_4 _5548_ (.A1(net134),
    .A2(_0470_),
    .B1(net204),
    .B2(_0473_),
    .C1(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__inv_2 _5549_ (.A(_1029_),
    .Y(_1068_));
 sky130_fd_sc_hd__a32o_1 _5550_ (.A1(_1036_),
    .A2(_0589_),
    .A3(_0862_),
    .B1(_0677_),
    .B2(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__o22a_1 _5551_ (.A1(net105),
    .A2(_0625_),
    .B1(net42),
    .B2(_0626_),
    .X(_1070_));
 sky130_fd_sc_hd__o221a_4 _5552_ (.A1(net144),
    .A2(_0492_),
    .B1(net207),
    .B2(_0624_),
    .C1(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__a22o_1 _5553_ (.A1(_1052_),
    .A2(_0612_),
    .B1(_0557_),
    .B2(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__mux2_1 _5554_ (.A0(_1022_),
    .A1(_1072_),
    .S(_0781_),
    .X(_1073_));
 sky130_fd_sc_hd__a22o_1 _5555_ (.A1(_0632_),
    .A2(_1021_),
    .B1(_1073_),
    .B2(_0631_),
    .X(_1074_));
 sky130_fd_sc_hd__a211o_1 _5556_ (.A1(_1069_),
    .A2(_0604_),
    .B1(_0535_),
    .C1(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__o22a_1 _5557_ (.A1(net103),
    .A2(_0123_),
    .B1(net40),
    .B2(_0122_),
    .X(_1076_));
 sky130_fd_sc_hd__o221a_4 _5558_ (.A1(net134),
    .A2(_0449_),
    .B1(net204),
    .B2(_0365_),
    .C1(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__a22o_1 _5559_ (.A1(_1077_),
    .A2(_0088_),
    .B1(_0111_),
    .B2(_1064_),
    .X(_1078_));
 sky130_fd_sc_hd__inv_2 _5560_ (.A(_1078_),
    .Y(_1079_));
 sky130_fd_sc_hd__o22a_1 _5561_ (.A1(net104),
    .A2(_0724_),
    .B1(net41),
    .B2(_0122_),
    .X(_1080_));
 sky130_fd_sc_hd__o221a_4 _5562_ (.A1(net143),
    .A2(_0449_),
    .B1(net205),
    .B2(_0365_),
    .C1(_1080_),
    .X(_1081_));
 sky130_fd_sc_hd__o22a_1 _5563_ (.A1(net105),
    .A2(_0724_),
    .B1(net42),
    .B2(_0725_),
    .X(_1082_));
 sky130_fd_sc_hd__o221a_4 _5564_ (.A1(net144),
    .A2(_0449_),
    .B1(net207),
    .B2(_0723_),
    .C1(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__a22o_1 _5565_ (.A1(_1081_),
    .A2(_0111_),
    .B1(_0730_),
    .B2(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__nor2_1 _5566_ (.A(_0761_),
    .B(_1084_),
    .Y(_1085_));
 sky130_fd_sc_hd__a21o_1 _5567_ (.A1(_0761_),
    .A2(_1079_),
    .B1(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__inv_2 _5568_ (.A(_1086_),
    .Y(_1087_));
 sky130_fd_sc_hd__o221a_1 _5569_ (.A1(_0461_),
    .A2(_1077_),
    .B1(_0463_),
    .B2(_1087_),
    .C1(_0670_),
    .X(_1088_));
 sky130_fd_sc_hd__a22o_2 _5570_ (.A1(_0567_),
    .A2(_1067_),
    .B1(_1075_),
    .B2(_1088_),
    .X(net604));
 sky130_fd_sc_hd__o22a_1 _5571_ (.A1(net106),
    .A2(_0625_),
    .B1(net43),
    .B2(_0626_),
    .X(_1089_));
 sky130_fd_sc_hd__o221a_4 _5572_ (.A1(net145),
    .A2(_0492_),
    .B1(net208),
    .B2(_0624_),
    .C1(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__a22o_1 _5573_ (.A1(_1071_),
    .A2(_0612_),
    .B1(_0557_),
    .B2(_1090_),
    .X(_1091_));
 sky130_fd_sc_hd__mux2_1 _5574_ (.A0(_1091_),
    .A1(_1053_),
    .S(_0718_),
    .X(_1092_));
 sky130_fd_sc_hd__inv_2 _5575_ (.A(net143),
    .Y(_1093_));
 sky130_fd_sc_hd__inv_2 _5576_ (.A(net205),
    .Y(_1094_));
 sky130_fd_sc_hd__a22oi_1 _5577_ (.A1(_0803_),
    .A2(net104),
    .B1(_0804_),
    .B2(net41),
    .Y(_1095_));
 sky130_fd_sc_hd__o221a_2 _5578_ (.A1(_1093_),
    .A2(_0425_),
    .B1(_1094_),
    .B2(_0430_),
    .C1(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__nor2_1 _5579_ (.A(_0910_),
    .B(_1096_),
    .Y(_1097_));
 sky130_fd_sc_hd__mux2_2 _5580_ (.A0(_1097_),
    .A1(_1030_),
    .S(_0799_),
    .X(_1098_));
 sky130_fd_sc_hd__inv_2 _5581_ (.A(_1096_),
    .Y(_1099_));
 sky130_fd_sc_hd__a32o_1 _5582_ (.A1(_1098_),
    .A2(_0588_),
    .A3(_0862_),
    .B1(_0441_),
    .B2(_1099_),
    .X(_1100_));
 sky130_fd_sc_hd__inv_2 _5583_ (.A(_1052_),
    .Y(_1101_));
 sky130_fd_sc_hd__nor2_1 _5584_ (.A(_0418_),
    .B(_1101_),
    .Y(_1102_));
 sky130_fd_sc_hd__a221o_2 _5585_ (.A1(_0419_),
    .A2(_1092_),
    .B1(_1100_),
    .B2(_0592_),
    .C1(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__mux2_1 _5586_ (.A0(_1103_),
    .A1(_1081_),
    .S(_0465_),
    .X(_1104_));
 sky130_fd_sc_hd__o22a_1 _5587_ (.A1(net104),
    .A2(_0475_),
    .B1(net41),
    .B2(_0479_),
    .X(_1105_));
 sky130_fd_sc_hd__o221a_4 _5588_ (.A1(net143),
    .A2(_0646_),
    .B1(net205),
    .B2(_0472_),
    .C1(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__mux2_1 _5589_ (.A0(_1104_),
    .A1(_1106_),
    .S(_0490_),
    .X(_1107_));
 sky130_fd_sc_hd__buf_1 _5590_ (.A(_1107_),
    .X(net605));
 sky130_fd_sc_hd__inv_2 _5591_ (.A(net144),
    .Y(_1108_));
 sky130_fd_sc_hd__inv_2 _5592_ (.A(net207),
    .Y(_1109_));
 sky130_fd_sc_hd__a22oi_1 _5593_ (.A1(_0432_),
    .A2(net105),
    .B1(_0435_),
    .B2(net42),
    .Y(_1110_));
 sky130_fd_sc_hd__o221a_2 _5594_ (.A1(_1108_),
    .A2(_0425_),
    .B1(_1109_),
    .B2(_0430_),
    .C1(_1110_),
    .X(_1111_));
 sky130_fd_sc_hd__inv_2 _5595_ (.A(_1111_),
    .Y(_1112_));
 sky130_fd_sc_hd__inv_2 _5596_ (.A(net146),
    .Y(_1113_));
 sky130_fd_sc_hd__inv_2 _5597_ (.A(net209),
    .Y(_1114_));
 sky130_fd_sc_hd__a22oi_1 _5598_ (.A1(_0263_),
    .A2(net107),
    .B1(_0434_),
    .B2(net44),
    .Y(_1115_));
 sky130_fd_sc_hd__o221a_2 _5599_ (.A1(_1113_),
    .A2(_0424_),
    .B1(_1114_),
    .B2(_0429_),
    .C1(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__inv_2 _5600_ (.A(_1116_),
    .Y(_1117_));
 sky130_fd_sc_hd__inv_2 _5601_ (.A(net145),
    .Y(_1118_));
 sky130_fd_sc_hd__inv_2 _5602_ (.A(net208),
    .Y(_1119_));
 sky130_fd_sc_hd__a22oi_1 _5603_ (.A1(_0263_),
    .A2(net106),
    .B1(_0804_),
    .B2(net43),
    .Y(_1120_));
 sky130_fd_sc_hd__o221a_2 _5604_ (.A1(_1118_),
    .A2(_0424_),
    .B1(_1119_),
    .B2(_0429_),
    .C1(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__nor2_1 _5605_ (.A(_4204_),
    .B(_1121_),
    .Y(_1122_));
 sky130_fd_sc_hd__nand2_1 _5606_ (.A(_1122_),
    .B(_0799_),
    .Y(_1123_));
 sky130_fd_sc_hd__inv_2 _5607_ (.A(_1123_),
    .Y(_1124_));
 sky130_fd_sc_hd__a31o_1 _5608_ (.A1(_1117_),
    .A2(_0522_),
    .A3(_0520_),
    .B1(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__nor2_1 _5609_ (.A(_0538_),
    .B(_1111_),
    .Y(_1126_));
 sky130_fd_sc_hd__nand2_1 _5610_ (.A(_1097_),
    .B(_0799_),
    .Y(_1127_));
 sky130_fd_sc_hd__inv_2 _5611_ (.A(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__a21o_1 _5612_ (.A1(_0523_),
    .A2(_1126_),
    .B1(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__or2_1 _5613_ (.A(_0704_),
    .B(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__o21ai_1 _5614_ (.A1(_0862_),
    .A2(_1125_),
    .B1(_1130_),
    .Y(_1131_));
 sky130_fd_sc_hd__clkinv_4 _5615_ (.A(_4186_),
    .Y(_1132_));
 sky130_fd_sc_hd__buf_8 _5616_ (.A(_1132_),
    .X(_1133_));
 sky130_fd_sc_hd__nand2_1 _5617_ (.A(_1131_),
    .B(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__a22o_1 _5618_ (.A1(_0677_),
    .A2(_1112_),
    .B1(_1134_),
    .B2(_0706_),
    .X(_1135_));
 sky130_fd_sc_hd__a22o_1 _5619_ (.A1(_1090_),
    .A2(_0612_),
    .B1(_0557_),
    .B2(_0995_),
    .X(_1136_));
 sky130_fd_sc_hd__mux2_1 _5620_ (.A0(_1136_),
    .A1(_1072_),
    .S(_0719_),
    .X(_1137_));
 sky130_fd_sc_hd__a22o_1 _5621_ (.A1(_0632_),
    .A2(_1071_),
    .B1(_1137_),
    .B2(_0631_),
    .X(_1138_));
 sky130_fd_sc_hd__a211o_1 _5622_ (.A1(_1135_),
    .A2(_0604_),
    .B1(_0535_),
    .C1(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__o22a_1 _5623_ (.A1(net107),
    .A2(_0123_),
    .B1(net44),
    .B2(_0122_),
    .X(_1140_));
 sky130_fd_sc_hd__o221a_4 _5624_ (.A1(net146),
    .A2(_0449_),
    .B1(net209),
    .B2(_0365_),
    .C1(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__inv_2 _5625_ (.A(_1141_),
    .Y(_1142_));
 sky130_fd_sc_hd__o22a_1 _5626_ (.A1(net106),
    .A2(_0724_),
    .B1(net43),
    .B2(_0725_),
    .X(_1143_));
 sky130_fd_sc_hd__o221a_4 _5627_ (.A1(net145),
    .A2(_0449_),
    .B1(net208),
    .B2(_0723_),
    .C1(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__nand2_1 _5628_ (.A(_1144_),
    .B(_0111_),
    .Y(_1145_));
 sky130_fd_sc_hd__o21ai_1 _5629_ (.A1(_0090_),
    .A2(_1142_),
    .B1(_1145_),
    .Y(_1146_));
 sky130_fd_sc_hd__inv_2 _5630_ (.A(_1146_),
    .Y(_1147_));
 sky130_fd_sc_hd__nand2_1 _5631_ (.A(_1147_),
    .B(_0841_),
    .Y(_1148_));
 sky130_fd_sc_hd__o21ai_1 _5632_ (.A1(_0841_),
    .A2(_1084_),
    .B1(_1148_),
    .Y(_1149_));
 sky130_fd_sc_hd__nand2_1 _5633_ (.A(_1149_),
    .B(_0462_),
    .Y(_1150_));
 sky130_fd_sc_hd__or2_1 _5634_ (.A(_0461_),
    .B(_1083_),
    .X(_1151_));
 sky130_fd_sc_hd__o22a_1 _5635_ (.A1(net105),
    .A2(_0474_),
    .B1(net42),
    .B2(_0478_),
    .X(_1152_));
 sky130_fd_sc_hd__o221a_4 _5636_ (.A1(net144),
    .A2(_0468_),
    .B1(net207),
    .B2(_0471_),
    .C1(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__o22a_1 _5637_ (.A1(net107),
    .A2(_0474_),
    .B1(net44),
    .B2(_0478_),
    .X(_1154_));
 sky130_fd_sc_hd__o221a_4 _5638_ (.A1(net146),
    .A2(_0468_),
    .B1(net209),
    .B2(_0471_),
    .C1(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__nand2_1 _5639_ (.A(_1155_),
    .B(_0888_),
    .Y(_1156_));
 sky130_fd_sc_hd__o22a_1 _5640_ (.A1(net106),
    .A2(_0474_),
    .B1(net43),
    .B2(_0478_),
    .X(_1157_));
 sky130_fd_sc_hd__o221a_4 _5641_ (.A1(net145),
    .A2(_0468_),
    .B1(net208),
    .B2(_0471_),
    .C1(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__nand2_1 _5642_ (.A(_1158_),
    .B(_0888_),
    .Y(_1159_));
 sky130_fd_sc_hd__mux2_1 _5643_ (.A0(_1156_),
    .A1(_1159_),
    .S(_0855_),
    .X(_1160_));
 sky130_fd_sc_hd__inv_2 _5644_ (.A(_1153_),
    .Y(_1161_));
 sky130_fd_sc_hd__nand2_1 _5645_ (.A(_1106_),
    .B(_0767_),
    .Y(_1162_));
 sky130_fd_sc_hd__o21ai_1 _5646_ (.A1(_0855_),
    .A2(_1161_),
    .B1(_1162_),
    .Y(_1163_));
 sky130_fd_sc_hd__nor2_1 _5647_ (.A(_0887_),
    .B(_1163_),
    .Y(_1164_));
 sky130_fd_sc_hd__a21oi_2 _5648_ (.A1(_1160_),
    .A2(_0887_),
    .B1(_1164_),
    .Y(_1165_));
 sky130_fd_sc_hd__a22o_1 _5649_ (.A1(_0645_),
    .A2(_1153_),
    .B1(_1165_),
    .B2(_0660_),
    .X(_1166_));
 sky130_fd_sc_hd__a41o_2 _5650_ (.A1(_1139_),
    .A2(_0636_),
    .A3(_1150_),
    .A4(_1151_),
    .B1(_1166_),
    .X(net606));
 sky130_fd_sc_hd__a22o_1 _5651_ (.A1(_1153_),
    .A2(_0767_),
    .B1(_0769_),
    .B2(_1158_),
    .X(_1167_));
 sky130_fd_sc_hd__o22a_1 _5652_ (.A1(net108),
    .A2(_0474_),
    .B1(net46),
    .B2(_0478_),
    .X(_1168_));
 sky130_fd_sc_hd__o221a_4 _5653_ (.A1(net147),
    .A2(_0468_),
    .B1(net210),
    .B2(_0471_),
    .C1(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__inv_2 _5654_ (.A(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__nand2_2 _5655_ (.A(_1155_),
    .B(_0767_),
    .Y(_1171_));
 sky130_fd_sc_hd__o21ai_2 _5656_ (.A1(_0855_),
    .A2(_1170_),
    .B1(_1171_),
    .Y(_1172_));
 sky130_fd_sc_hd__mux2_1 _5657_ (.A0(_1167_),
    .A1(_1172_),
    .S(_0886_),
    .X(_1173_));
 sky130_fd_sc_hd__inv_2 _5658_ (.A(_1121_),
    .Y(_1174_));
 sky130_fd_sc_hd__nand2_1 _5659_ (.A(_1090_),
    .B(_4106_),
    .Y(_1175_));
 sky130_fd_sc_hd__nand2_1 _5660_ (.A(_1175_),
    .B(_4235_),
    .Y(_1176_));
 sky130_fd_sc_hd__inv_2 _5661_ (.A(net147),
    .Y(_1177_));
 sky130_fd_sc_hd__inv_2 _5662_ (.A(net210),
    .Y(_1178_));
 sky130_fd_sc_hd__a22oi_1 _5663_ (.A1(_0803_),
    .A2(net108),
    .B1(_0804_),
    .B2(net46),
    .Y(_1179_));
 sky130_fd_sc_hd__o221a_2 _5664_ (.A1(_1177_),
    .A2(_0424_),
    .B1(_1178_),
    .B2(_0429_),
    .C1(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__nor2_1 _5665_ (.A(_0910_),
    .B(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__or3_1 _5666_ (.A(_4127_),
    .B(_4119_),
    .C(_1116_),
    .X(_1182_));
 sky130_fd_sc_hd__inv_2 _5667_ (.A(_1182_),
    .Y(_1183_));
 sky130_fd_sc_hd__a21o_1 _5668_ (.A1(_0522_),
    .A2(_1181_),
    .B1(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__mux2_1 _5669_ (.A0(_1122_),
    .A1(_1126_),
    .S(_0800_),
    .X(_1185_));
 sky130_fd_sc_hd__or2_1 _5670_ (.A(_0704_),
    .B(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__o21ai_1 _5671_ (.A1(_0862_),
    .A2(_1184_),
    .B1(_1186_),
    .Y(_1187_));
 sky130_fd_sc_hd__nor2_1 _5672_ (.A(_0444_),
    .B(_1187_),
    .Y(_1188_));
 sky130_fd_sc_hd__a221o_1 _5673_ (.A1(_0677_),
    .A2(_1174_),
    .B1(_0548_),
    .B2(_1176_),
    .C1(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__or2_1 _5674_ (.A(_0718_),
    .B(_0998_),
    .X(_1190_));
 sky130_fd_sc_hd__o21ai_1 _5675_ (.A1(_0833_),
    .A2(_1091_),
    .B1(_1190_),
    .Y(_1191_));
 sky130_fd_sc_hd__o21ai_1 _5676_ (.A1(_0555_),
    .A2(_1191_),
    .B1(_0631_),
    .Y(_1192_));
 sky130_fd_sc_hd__a21oi_1 _5677_ (.A1(_1175_),
    .A2(_0632_),
    .B1(_0633_),
    .Y(_1193_));
 sky130_fd_sc_hd__a32o_1 _5678_ (.A1(_1189_),
    .A2(_1192_),
    .A3(_1193_),
    .B1(_0535_),
    .B2(_1144_),
    .X(_1194_));
 sky130_fd_sc_hd__and2_1 _5679_ (.A(_1158_),
    .B(_0484_),
    .X(_1195_));
 sky130_fd_sc_hd__a221o_2 _5680_ (.A1(_0660_),
    .A2(_1173_),
    .B1(_1194_),
    .B2(_0636_),
    .C1(_1195_),
    .X(net607));
 sky130_fd_sc_hd__inv_2 _5681_ (.A(_1000_),
    .Y(_1196_));
 sky130_fd_sc_hd__nand2_1 _5682_ (.A(_0997_),
    .B(_0613_),
    .Y(_1197_));
 sky130_fd_sc_hd__o21ai_1 _5683_ (.A1(_0555_),
    .A2(_1196_),
    .B1(_1197_),
    .Y(_1198_));
 sky130_fd_sc_hd__mux2_1 _5684_ (.A0(_1136_),
    .A1(_1198_),
    .S(_0781_),
    .X(_1199_));
 sky130_fd_sc_hd__inv_2 _5685_ (.A(net211),
    .Y(_1200_));
 sky130_fd_sc_hd__inv_2 _5686_ (.A(net148),
    .Y(_1201_));
 sky130_fd_sc_hd__a22oi_1 _5687_ (.A1(_0263_),
    .A2(net109),
    .B1(_0434_),
    .B2(net47),
    .Y(_1202_));
 sky130_fd_sc_hd__o221a_2 _5688_ (.A1(_1200_),
    .A2(_0429_),
    .B1(_1201_),
    .B2(_0424_),
    .C1(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__nor2_1 _5689_ (.A(_4204_),
    .B(_1203_),
    .Y(_1204_));
 sky130_fd_sc_hd__nand2_1 _5690_ (.A(_1181_),
    .B(_0799_),
    .Y(_1205_));
 sky130_fd_sc_hd__inv_2 _5691_ (.A(_1205_),
    .Y(_1206_));
 sky130_fd_sc_hd__a21o_1 _5692_ (.A1(_0522_),
    .A2(_1204_),
    .B1(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__mux2_1 _5693_ (.A0(_1125_),
    .A1(_1207_),
    .S(_0703_),
    .X(_1208_));
 sky130_fd_sc_hd__a221o_1 _5694_ (.A1(_0677_),
    .A2(_1117_),
    .B1(_1208_),
    .B2(_0706_),
    .C1(_0422_),
    .X(_1209_));
 sky130_fd_sc_hd__o221a_1 _5695_ (.A1(_0418_),
    .A2(_0995_),
    .B1(_0420_),
    .B2(_1199_),
    .C1(_1209_),
    .X(_1210_));
 sky130_fd_sc_hd__or2_1 _5696_ (.A(_0535_),
    .B(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__o22a_1 _5697_ (.A1(net108),
    .A2(_0454_),
    .B1(net46),
    .B2(_0456_),
    .X(_1212_));
 sky130_fd_sc_hd__o221a_4 _5698_ (.A1(net147),
    .A2(_0450_),
    .B1(net210),
    .B2(_0452_),
    .C1(_1212_),
    .X(_1213_));
 sky130_fd_sc_hd__o22a_1 _5699_ (.A1(net109),
    .A2(_0454_),
    .B1(net47),
    .B2(_0456_),
    .X(_1214_));
 sky130_fd_sc_hd__o221a_4 _5700_ (.A1(net211),
    .A2(_0452_),
    .B1(net148),
    .B2(_0450_),
    .C1(_1214_),
    .X(_1215_));
 sky130_fd_sc_hd__a22o_1 _5701_ (.A1(_1213_),
    .A2(_0729_),
    .B1(_0730_),
    .B2(_1215_),
    .X(_1216_));
 sky130_fd_sc_hd__nand2_1 _5702_ (.A(_1147_),
    .B(_0761_),
    .Y(_1217_));
 sky130_fd_sc_hd__o21ai_1 _5703_ (.A1(_0761_),
    .A2(_1216_),
    .B1(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__inv_2 _5704_ (.A(_1218_),
    .Y(_1219_));
 sky130_fd_sc_hd__o221a_1 _5705_ (.A1(_0461_),
    .A2(_1141_),
    .B1(_0463_),
    .B2(_1219_),
    .C1(_0670_),
    .X(_1220_));
 sky130_fd_sc_hd__a22o_2 _5706_ (.A1(_0567_),
    .A2(_1155_),
    .B1(_1211_),
    .B2(_1220_),
    .X(net608));
 sky130_fd_sc_hd__inv_2 _5707_ (.A(_1005_),
    .Y(_1221_));
 sky130_fd_sc_hd__a221o_1 _5708_ (.A1(_0417_),
    .A2(_0997_),
    .B1(_1221_),
    .B2(_0419_),
    .C1(_0465_),
    .X(_1222_));
 sky130_fd_sc_hd__inv_2 _5709_ (.A(_1180_),
    .Y(_1223_));
 sky130_fd_sc_hd__mux2_1 _5710_ (.A0(_1204_),
    .A1(_1043_),
    .S(_4127_),
    .X(_1224_));
 sky130_fd_sc_hd__or2_1 _5711_ (.A(_0813_),
    .B(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__o21ai_1 _5712_ (.A1(_0703_),
    .A2(_1184_),
    .B1(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__inv_2 _5713_ (.A(_1226_),
    .Y(_1227_));
 sky130_fd_sc_hd__a22o_1 _5714_ (.A1(_0677_),
    .A2(_1223_),
    .B1(_1227_),
    .B2(_0443_),
    .X(_1228_));
 sky130_fd_sc_hd__and2_1 _5715_ (.A(_1228_),
    .B(_0592_),
    .X(_1229_));
 sky130_fd_sc_hd__o221a_1 _5716_ (.A1(_0667_),
    .A2(_1213_),
    .B1(_1222_),
    .B2(_1229_),
    .C1(_0670_),
    .X(_1230_));
 sky130_fd_sc_hd__a221o_1 _5717_ (.A1(_0645_),
    .A2(_1169_),
    .B1(_0660_),
    .B2(_1172_),
    .C1(_1230_),
    .X(net609));
 sky130_fd_sc_hd__o22a_1 _5718_ (.A1(net109),
    .A2(_0186_),
    .B1(net47),
    .B2(_0477_),
    .X(_1231_));
 sky130_fd_sc_hd__o221a_4 _5719_ (.A1(net211),
    .A2(_0185_),
    .B1(net148),
    .B2(_0467_),
    .C1(_1231_),
    .X(_1232_));
 sky130_fd_sc_hd__a22o_1 _5720_ (.A1(_1169_),
    .A2(_0766_),
    .B1(_0769_),
    .B2(_1232_),
    .X(_1233_));
 sky130_fd_sc_hd__a21o_1 _5721_ (.A1(_1000_),
    .A2(_4106_),
    .B1(_0056_),
    .X(_1234_));
 sky130_fd_sc_hd__inv_2 _5722_ (.A(net150),
    .Y(_1235_));
 sky130_fd_sc_hd__inv_2 _5723_ (.A(net213),
    .Y(_1236_));
 sky130_fd_sc_hd__a22oi_1 _5724_ (.A1(_0263_),
    .A2(net113),
    .B1(_0434_),
    .B2(net49),
    .Y(_1237_));
 sky130_fd_sc_hd__o221a_2 _5725_ (.A1(_1235_),
    .A2(_0424_),
    .B1(_1236_),
    .B2(_0429_),
    .C1(_1237_),
    .X(_1238_));
 sky130_fd_sc_hd__nor2_1 _5726_ (.A(_4204_),
    .B(_1238_),
    .Y(_1239_));
 sky130_fd_sc_hd__inv_2 _5727_ (.A(_1044_),
    .Y(_1240_));
 sky130_fd_sc_hd__a21o_1 _5728_ (.A1(_0523_),
    .A2(_1239_),
    .B1(_1240_),
    .X(_1241_));
 sky130_fd_sc_hd__mux2_1 _5729_ (.A0(_1241_),
    .A1(_1207_),
    .S(_0862_),
    .X(_1242_));
 sky130_fd_sc_hd__nor2_1 _5730_ (.A(_0591_),
    .B(_1203_),
    .Y(_1243_));
 sky130_fd_sc_hd__a221o_1 _5731_ (.A1(_0548_),
    .A2(_1234_),
    .B1(_1242_),
    .B2(_0706_),
    .C1(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__o22a_1 _5732_ (.A1(net113),
    .A2(_0036_),
    .B1(net49),
    .B2(_4289_),
    .X(_1245_));
 sky130_fd_sc_hd__o221a_4 _5733_ (.A1(net150),
    .A2(_0407_),
    .B1(net213),
    .B2(_0038_),
    .C1(_1245_),
    .X(_1246_));
 sky130_fd_sc_hd__a22o_1 _5734_ (.A1(_1002_),
    .A2(_0612_),
    .B1(_0557_),
    .B2(_1246_),
    .X(_1247_));
 sky130_fd_sc_hd__or2_1 _5735_ (.A(_0833_),
    .B(_1198_),
    .X(_1248_));
 sky130_fd_sc_hd__o21ai_1 _5736_ (.A1(_0719_),
    .A2(_1247_),
    .B1(_1248_),
    .Y(_1249_));
 sky130_fd_sc_hd__nand2_1 _5737_ (.A(_1249_),
    .B(_0631_),
    .Y(_1250_));
 sky130_fd_sc_hd__or3_1 _5738_ (.A(_4105_),
    .B(_0056_),
    .C(_1000_),
    .X(_1251_));
 sky130_fd_sc_hd__a31o_2 _5739_ (.A1(_1244_),
    .A2(_1250_),
    .A3(_1251_),
    .B1(_0535_),
    .X(_1252_));
 sky130_fd_sc_hd__o21a_1 _5740_ (.A1(_0682_),
    .A2(_1215_),
    .B1(_0601_),
    .X(_1253_));
 sky130_fd_sc_hd__and2_1 _5741_ (.A(_1232_),
    .B(_0484_),
    .X(_1254_));
 sky130_fd_sc_hd__a221o_2 _5742_ (.A1(_0660_),
    .A2(_1233_),
    .B1(_1252_),
    .B2(_1253_),
    .C1(_1254_),
    .X(net610));
 sky130_fd_sc_hd__o22a_1 _5743_ (.A1(net110),
    .A2(_0186_),
    .B1(net48),
    .B2(_0477_),
    .X(_1255_));
 sky130_fd_sc_hd__o221a_4 _5744_ (.A1(net149),
    .A2(_0467_),
    .B1(net212),
    .B2(_0185_),
    .C1(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__inv_2 _5745_ (.A(_1042_),
    .Y(_1257_));
 sky130_fd_sc_hd__a22o_1 _5746_ (.A1(_4149_),
    .A2(net152),
    .B1(_4147_),
    .B2(net214),
    .X(_1258_));
 sky130_fd_sc_hd__a221oi_4 _5747_ (.A1(net50),
    .A2(_0434_),
    .B1(net114),
    .B2(_0803_),
    .C1(_1258_),
    .Y(_1259_));
 sky130_fd_sc_hd__inv_2 _5748_ (.A(_1259_),
    .Y(_1260_));
 sky130_fd_sc_hd__nand2_1 _5749_ (.A(_1239_),
    .B(_4114_),
    .Y(_1261_));
 sky130_fd_sc_hd__inv_2 _5750_ (.A(_1261_),
    .Y(_1262_));
 sky130_fd_sc_hd__a31o_1 _5751_ (.A1(_1260_),
    .A2(_4127_),
    .A3(_0520_),
    .B1(_1262_),
    .X(_1263_));
 sky130_fd_sc_hd__or2_1 _5752_ (.A(_0703_),
    .B(_1224_),
    .X(_1264_));
 sky130_fd_sc_hd__o21ai_1 _5753_ (.A1(_0813_),
    .A2(_1263_),
    .B1(_1264_),
    .Y(_1265_));
 sky130_fd_sc_hd__inv_2 _5754_ (.A(_1265_),
    .Y(_1266_));
 sky130_fd_sc_hd__a22o_1 _5755_ (.A1(_0441_),
    .A2(_1257_),
    .B1(_1266_),
    .B2(_0443_),
    .X(_1267_));
 sky130_fd_sc_hd__o22a_1 _5756_ (.A1(net114),
    .A2(_0411_),
    .B1(net50),
    .B2(_0413_),
    .X(_1268_));
 sky130_fd_sc_hd__o221a_4 _5757_ (.A1(net152),
    .A2(_0407_),
    .B1(net214),
    .B2(_0038_),
    .C1(_1268_),
    .X(_1269_));
 sky130_fd_sc_hd__a22o_1 _5758_ (.A1(_1246_),
    .A2(_4265_),
    .B1(_0510_),
    .B2(_1269_),
    .X(_1270_));
 sky130_fd_sc_hd__inv_2 _5759_ (.A(_1270_),
    .Y(_1271_));
 sky130_fd_sc_hd__nand2_1 _5760_ (.A(_1271_),
    .B(_0781_),
    .Y(_1272_));
 sky130_fd_sc_hd__o21ai_2 _5761_ (.A1(_0781_),
    .A2(_1003_),
    .B1(_1272_),
    .Y(_1273_));
 sky130_fd_sc_hd__nor2_1 _5762_ (.A(_0420_),
    .B(_1273_),
    .Y(_1274_));
 sky130_fd_sc_hd__a221o_1 _5763_ (.A1(_0417_),
    .A2(_1002_),
    .B1(_1267_),
    .B2(_0592_),
    .C1(_1274_),
    .X(_1275_));
 sky130_fd_sc_hd__o22a_1 _5764_ (.A1(net110),
    .A2(_0123_),
    .B1(net48),
    .B2(_0122_),
    .X(_1276_));
 sky130_fd_sc_hd__o221a_4 _5765_ (.A1(net149),
    .A2(_0449_),
    .B1(net212),
    .B2(_0365_),
    .C1(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__mux2_2 _5766_ (.A0(_1275_),
    .A1(_1277_),
    .S(_0633_),
    .X(_1278_));
 sky130_fd_sc_hd__inv_2 _5767_ (.A(_0886_),
    .Y(_1279_));
 sky130_fd_sc_hd__buf_4 _5768_ (.A(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__o22a_1 _5769_ (.A1(net113),
    .A2(_0186_),
    .B1(net49),
    .B2(_0477_),
    .X(_1281_));
 sky130_fd_sc_hd__o221a_4 _5770_ (.A1(net150),
    .A2(_0467_),
    .B1(net213),
    .B2(_0185_),
    .C1(_1281_),
    .X(_1282_));
 sky130_fd_sc_hd__o22a_1 _5771_ (.A1(net114),
    .A2(_0186_),
    .B1(net50),
    .B2(_0477_),
    .X(_1283_));
 sky130_fd_sc_hd__o221a_4 _5772_ (.A1(net152),
    .A2(_0467_),
    .B1(net214),
    .B2(_0185_),
    .C1(_1283_),
    .X(_1284_));
 sky130_fd_sc_hd__a22o_1 _5773_ (.A1(_1282_),
    .A2(_0766_),
    .B1(_0198_),
    .B2(_1284_),
    .X(_1285_));
 sky130_fd_sc_hd__inv_2 _5774_ (.A(_1285_),
    .Y(_1286_));
 sky130_fd_sc_hd__a22o_1 _5775_ (.A1(_1232_),
    .A2(_0766_),
    .B1(_0198_),
    .B2(_1256_),
    .X(_1287_));
 sky130_fd_sc_hd__nand2_1 _5776_ (.A(_1287_),
    .B(_1280_),
    .Y(_1288_));
 sky130_fd_sc_hd__o21ai_1 _5777_ (.A1(_1280_),
    .A2(_1286_),
    .B1(_1288_),
    .Y(_1289_));
 sky130_fd_sc_hd__and2_1 _5778_ (.A(_1289_),
    .B(_0487_),
    .X(_1290_));
 sky130_fd_sc_hd__a221o_2 _5779_ (.A1(_0645_),
    .A2(_1256_),
    .B1(_1278_),
    .B2(_0636_),
    .C1(_1290_),
    .X(net611));
 sky130_fd_sc_hd__buf_8 _5780_ (.A(_4263_),
    .X(_1291_));
 sky130_fd_sc_hd__nand2_1 _5781_ (.A(_1247_),
    .B(_0718_),
    .Y(_1292_));
 sky130_fd_sc_hd__nand2_1 _5782_ (.A(_1292_),
    .B(_4233_),
    .Y(_1293_));
 sky130_fd_sc_hd__inv_2 _5783_ (.A(_1238_),
    .Y(_1294_));
 sky130_fd_sc_hd__a22o_1 _5784_ (.A1(_0441_),
    .A2(_1294_),
    .B1(_1293_),
    .B2(_0288_),
    .X(_1295_));
 sky130_fd_sc_hd__a32o_1 _5785_ (.A1(_0589_),
    .A2(_0862_),
    .A3(_1241_),
    .B1(_1295_),
    .B2(_0550_),
    .X(_1296_));
 sky130_fd_sc_hd__o221a_2 _5786_ (.A1(_1291_),
    .A2(_1293_),
    .B1(_0418_),
    .B2(_1246_),
    .C1(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__o22a_1 _5787_ (.A1(net114),
    .A2(_0454_),
    .B1(net50),
    .B2(_0456_),
    .X(_1298_));
 sky130_fd_sc_hd__o221a_4 _5788_ (.A1(net152),
    .A2(_0637_),
    .B1(net214),
    .B2(_0452_),
    .C1(_1298_),
    .X(_1299_));
 sky130_fd_sc_hd__o22a_1 _5789_ (.A1(net115),
    .A2(_0724_),
    .B1(net51),
    .B2(_0725_),
    .X(_1300_));
 sky130_fd_sc_hd__o221a_4 _5790_ (.A1(net153),
    .A2(_0637_),
    .B1(net215),
    .B2(_0723_),
    .C1(_1300_),
    .X(_1301_));
 sky130_fd_sc_hd__a22o_1 _5791_ (.A1(_1299_),
    .A2(_0572_),
    .B1(_0771_),
    .B2(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__o22a_1 _5792_ (.A1(net113),
    .A2(_0724_),
    .B1(net49),
    .B2(_0725_),
    .X(_1303_));
 sky130_fd_sc_hd__o221a_4 _5793_ (.A1(net150),
    .A2(_0449_),
    .B1(net213),
    .B2(_0723_),
    .C1(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__a22o_1 _5794_ (.A1(_1277_),
    .A2(_0111_),
    .B1(_0730_),
    .B2(_1304_),
    .X(_1305_));
 sky130_fd_sc_hd__inv_2 _5795_ (.A(_1305_),
    .Y(_1306_));
 sky130_fd_sc_hd__nand2_1 _5796_ (.A(_1306_),
    .B(_0761_),
    .Y(_1307_));
 sky130_fd_sc_hd__o21ai_2 _5797_ (.A1(_0761_),
    .A2(_1302_),
    .B1(_1307_),
    .Y(_1308_));
 sky130_fd_sc_hd__nand2_1 _5798_ (.A(_1308_),
    .B(_0462_),
    .Y(_1309_));
 sky130_fd_sc_hd__inv_2 _5799_ (.A(_1304_),
    .Y(_1310_));
 sky130_fd_sc_hd__nand2_1 _5800_ (.A(_1310_),
    .B(_0460_),
    .Y(_1311_));
 sky130_fd_sc_hd__o2111a_1 _5801_ (.A1(_0535_),
    .A2(_1297_),
    .B1(_0670_),
    .C1(_1309_),
    .D1(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__a21o_1 _5802_ (.A1(_0567_),
    .A2(_1282_),
    .B1(_1312_),
    .X(net614));
 sky130_fd_sc_hd__inv_2 _5803_ (.A(_1269_),
    .Y(_1313_));
 sky130_fd_sc_hd__inv_2 _5804_ (.A(net154),
    .Y(_1314_));
 sky130_fd_sc_hd__inv_2 _5805_ (.A(net216),
    .Y(_1315_));
 sky130_fd_sc_hd__a22oi_1 _5806_ (.A1(_0803_),
    .A2(net116),
    .B1(_0804_),
    .B2(net52),
    .Y(_1316_));
 sky130_fd_sc_hd__o221a_2 _5807_ (.A1(_1314_),
    .A2(_0425_),
    .B1(_1315_),
    .B2(_0430_),
    .C1(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__nor2_1 _5808_ (.A(_0910_),
    .B(_1317_),
    .Y(_1318_));
 sky130_fd_sc_hd__inv_2 _5809_ (.A(net153),
    .Y(_1319_));
 sky130_fd_sc_hd__inv_2 _5810_ (.A(net215),
    .Y(_1320_));
 sky130_fd_sc_hd__a22oi_1 _5811_ (.A1(_0803_),
    .A2(net115),
    .B1(_0804_),
    .B2(net51),
    .Y(_1321_));
 sky130_fd_sc_hd__o221a_2 _5812_ (.A1(_1319_),
    .A2(_0425_),
    .B1(_1320_),
    .B2(_0430_),
    .C1(_1321_),
    .X(_1322_));
 sky130_fd_sc_hd__nor2_1 _5813_ (.A(_0910_),
    .B(_1322_),
    .Y(_1323_));
 sky130_fd_sc_hd__mux2_2 _5814_ (.A0(_1318_),
    .A1(_1323_),
    .S(_0799_),
    .X(_1324_));
 sky130_fd_sc_hd__mux2_1 _5815_ (.A0(_1263_),
    .A1(_1324_),
    .S(_0704_),
    .X(_1325_));
 sky130_fd_sc_hd__nand2_1 _5816_ (.A(_1325_),
    .B(_0706_),
    .Y(_1326_));
 sky130_fd_sc_hd__nor2_1 _5817_ (.A(_0591_),
    .B(_1259_),
    .Y(_1327_));
 sky130_fd_sc_hd__o21ai_1 _5818_ (.A1(_0548_),
    .A2(_1327_),
    .B1(_0550_),
    .Y(_1328_));
 sky130_fd_sc_hd__a22o_1 _5819_ (.A1(_0422_),
    .A2(_1313_),
    .B1(_1326_),
    .B2(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__nand2_1 _5820_ (.A(_1329_),
    .B(_0668_),
    .Y(_1330_));
 sky130_fd_sc_hd__o21a_1 _5821_ (.A1(_0668_),
    .A2(_1299_),
    .B1(_0670_),
    .X(_1331_));
 sky130_fd_sc_hd__a22o_2 _5822_ (.A1(_0567_),
    .A2(_1284_),
    .B1(_1330_),
    .B2(_1331_),
    .X(net615));
 sky130_fd_sc_hd__o22a_1 _5823_ (.A1(net115),
    .A2(_0186_),
    .B1(net51),
    .B2(_0477_),
    .X(_1332_));
 sky130_fd_sc_hd__o221a_4 _5824_ (.A1(net153),
    .A2(_0467_),
    .B1(net215),
    .B2(_0185_),
    .C1(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__o22a_1 _5825_ (.A1(net115),
    .A2(_0036_),
    .B1(net51),
    .B2(_4289_),
    .X(_1334_));
 sky130_fd_sc_hd__o221a_4 _5826_ (.A1(net153),
    .A2(_0039_),
    .B1(net215),
    .B2(_0038_),
    .C1(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__nand2_1 _5827_ (.A(_1335_),
    .B(_4106_),
    .Y(_1336_));
 sky130_fd_sc_hd__nand2_1 _5828_ (.A(_1336_),
    .B(_4235_),
    .Y(_1337_));
 sky130_fd_sc_hd__or3_1 _5829_ (.A(_4127_),
    .B(_4119_),
    .C(_1259_),
    .X(_1338_));
 sky130_fd_sc_hd__inv_2 _5830_ (.A(_1338_),
    .Y(_1339_));
 sky130_fd_sc_hd__a21oi_1 _5831_ (.A1(_0523_),
    .A2(_1323_),
    .B1(_1339_),
    .Y(_1340_));
 sky130_fd_sc_hd__nor2_1 _5832_ (.A(_0704_),
    .B(_1340_),
    .Y(_1341_));
 sky130_fd_sc_hd__nor2_1 _5833_ (.A(_0591_),
    .B(_1322_),
    .Y(_1342_));
 sky130_fd_sc_hd__a221o_1 _5834_ (.A1(_0548_),
    .A2(_1337_),
    .B1(_1341_),
    .B2(_0589_),
    .C1(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__o22a_1 _5835_ (.A1(net117),
    .A2(_0036_),
    .B1(net53),
    .B2(_4289_),
    .X(_1344_));
 sky130_fd_sc_hd__o221a_4 _5836_ (.A1(net155),
    .A2(_0039_),
    .B1(net218),
    .B2(_0038_),
    .C1(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__o22a_1 _5837_ (.A1(net116),
    .A2(_0036_),
    .B1(net52),
    .B2(_4289_),
    .X(_1346_));
 sky130_fd_sc_hd__o221a_4 _5838_ (.A1(net154),
    .A2(_0407_),
    .B1(net216),
    .B2(_0038_),
    .C1(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__a22o_1 _5839_ (.A1(_1345_),
    .A2(_0558_),
    .B1(_0613_),
    .B2(_1347_),
    .X(_1348_));
 sky130_fd_sc_hd__a22o_1 _5840_ (.A1(_1335_),
    .A2(_0510_),
    .B1(_0612_),
    .B2(_1269_),
    .X(_1349_));
 sky130_fd_sc_hd__inv_2 _5841_ (.A(_1349_),
    .Y(_1350_));
 sky130_fd_sc_hd__nand2_1 _5842_ (.A(_1350_),
    .B(_0719_),
    .Y(_1351_));
 sky130_fd_sc_hd__o21ai_2 _5843_ (.A1(_0719_),
    .A2(_1348_),
    .B1(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__nand2_1 _5844_ (.A(_1352_),
    .B(_0631_),
    .Y(_1353_));
 sky130_fd_sc_hd__nand2_1 _5845_ (.A(_1336_),
    .B(_0632_),
    .Y(_1354_));
 sky130_fd_sc_hd__a31o_2 _5846_ (.A1(_1343_),
    .A2(_1353_),
    .A3(_1354_),
    .B1(_0535_),
    .X(_1355_));
 sky130_fd_sc_hd__o21a_1 _5847_ (.A1(_0682_),
    .A2(_1301_),
    .B1(_0601_),
    .X(_1356_));
 sky130_fd_sc_hd__a22o_1 _5848_ (.A1(_1284_),
    .A2(_0766_),
    .B1(_0198_),
    .B2(_1333_),
    .X(_1357_));
 sky130_fd_sc_hd__inv_2 _5849_ (.A(_1357_),
    .Y(_1358_));
 sky130_fd_sc_hd__nor2_1 _5850_ (.A(_0488_),
    .B(_1358_),
    .Y(_1359_));
 sky130_fd_sc_hd__a221o_2 _5851_ (.A1(_0645_),
    .A2(_1333_),
    .B1(_1355_),
    .B2(_1356_),
    .C1(_1359_),
    .X(net616));
 sky130_fd_sc_hd__o22a_1 _5852_ (.A1(net116),
    .A2(_0474_),
    .B1(net52),
    .B2(_0478_),
    .X(_1360_));
 sky130_fd_sc_hd__o221a_4 _5853_ (.A1(net154),
    .A2(_0468_),
    .B1(net216),
    .B2(_0471_),
    .C1(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__a22o_1 _5854_ (.A1(_1335_),
    .A2(_4265_),
    .B1(_0510_),
    .B2(_1347_),
    .X(_1362_));
 sky130_fd_sc_hd__inv_2 _5855_ (.A(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__nand2_1 _5856_ (.A(_1363_),
    .B(_0718_),
    .Y(_1364_));
 sky130_fd_sc_hd__inv_2 _5857_ (.A(_1345_),
    .Y(_1365_));
 sky130_fd_sc_hd__o22a_1 _5858_ (.A1(net118),
    .A2(_0411_),
    .B1(net54),
    .B2(_0413_),
    .X(_1366_));
 sky130_fd_sc_hd__o221a_4 _5859_ (.A1(net156),
    .A2(_0407_),
    .B1(net219),
    .B2(_0409_),
    .C1(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__nand2_1 _5860_ (.A(_1367_),
    .B(_4272_),
    .Y(_1368_));
 sky130_fd_sc_hd__o22a_1 _5861_ (.A1(_4287_),
    .A2(_1365_),
    .B1(_4253_),
    .B2(_1368_),
    .X(_1369_));
 sky130_fd_sc_hd__nand2_1 _5862_ (.A(_1369_),
    .B(_0781_),
    .Y(_1370_));
 sky130_fd_sc_hd__nand2_1 _5863_ (.A(_1364_),
    .B(_1370_),
    .Y(_1371_));
 sky130_fd_sc_hd__inv_2 _5864_ (.A(_1371_),
    .Y(_1372_));
 sky130_fd_sc_hd__inv_2 _5865_ (.A(_1317_),
    .Y(_1373_));
 sky130_fd_sc_hd__inv_2 _5866_ (.A(net156),
    .Y(_1374_));
 sky130_fd_sc_hd__inv_2 _5867_ (.A(net219),
    .Y(_1375_));
 sky130_fd_sc_hd__a22oi_1 _5868_ (.A1(_0803_),
    .A2(net118),
    .B1(_0804_),
    .B2(net54),
    .Y(_1376_));
 sky130_fd_sc_hd__o221a_2 _5869_ (.A1(_1374_),
    .A2(_0425_),
    .B1(_1375_),
    .B2(_0430_),
    .C1(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__nor2_1 _5870_ (.A(_0910_),
    .B(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__inv_2 _5871_ (.A(net155),
    .Y(_1379_));
 sky130_fd_sc_hd__inv_2 _5872_ (.A(net218),
    .Y(_1380_));
 sky130_fd_sc_hd__a22oi_1 _5873_ (.A1(_0803_),
    .A2(net117),
    .B1(_0804_),
    .B2(net53),
    .Y(_1381_));
 sky130_fd_sc_hd__o221a_2 _5874_ (.A1(_1379_),
    .A2(_0425_),
    .B1(_1380_),
    .B2(_0430_),
    .C1(_1381_),
    .X(_1382_));
 sky130_fd_sc_hd__nor2_1 _5875_ (.A(_0910_),
    .B(_1382_),
    .Y(_1383_));
 sky130_fd_sc_hd__mux2_1 _5876_ (.A0(_1378_),
    .A1(_1383_),
    .S(_0799_),
    .X(_1384_));
 sky130_fd_sc_hd__mux2_1 _5877_ (.A0(_1384_),
    .A1(_1324_),
    .S(_0813_),
    .X(_1385_));
 sky130_fd_sc_hd__a22o_1 _5878_ (.A1(_0441_),
    .A2(_1373_),
    .B1(_1385_),
    .B2(_0443_),
    .X(_1386_));
 sky130_fd_sc_hd__and2_1 _5879_ (.A(_1347_),
    .B(_0417_),
    .X(_1387_));
 sky130_fd_sc_hd__a221o_2 _5880_ (.A1(_0419_),
    .A2(_1372_),
    .B1(_1386_),
    .B2(_0592_),
    .C1(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__o22a_1 _5881_ (.A1(net116),
    .A2(_0724_),
    .B1(net52),
    .B2(_0725_),
    .X(_1389_));
 sky130_fd_sc_hd__o221a_4 _5882_ (.A1(net154),
    .A2(_0637_),
    .B1(net216),
    .B2(_0723_),
    .C1(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__mux2_1 _5883_ (.A0(_1388_),
    .A1(_1390_),
    .S(_0633_),
    .X(_1391_));
 sky130_fd_sc_hd__o22a_1 _5884_ (.A1(net117),
    .A2(_0186_),
    .B1(net53),
    .B2(_0477_),
    .X(_1392_));
 sky130_fd_sc_hd__o221a_4 _5885_ (.A1(net155),
    .A2(_0467_),
    .B1(net218),
    .B2(_0185_),
    .C1(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__o22a_1 _5886_ (.A1(net118),
    .A2(_0186_),
    .B1(net54),
    .B2(_0477_),
    .X(_1394_));
 sky130_fd_sc_hd__o221a_4 _5887_ (.A1(net156),
    .A2(_0467_),
    .B1(net219),
    .B2(_0185_),
    .C1(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__a22o_1 _5888_ (.A1(_1393_),
    .A2(_0766_),
    .B1(_0198_),
    .B2(_1395_),
    .X(_1396_));
 sky130_fd_sc_hd__inv_2 _5889_ (.A(_1396_),
    .Y(_1397_));
 sky130_fd_sc_hd__a22o_1 _5890_ (.A1(_1333_),
    .A2(_0766_),
    .B1(_0769_),
    .B2(_1361_),
    .X(_1398_));
 sky130_fd_sc_hd__nand2_1 _5891_ (.A(_1398_),
    .B(_1280_),
    .Y(_1399_));
 sky130_fd_sc_hd__o21ai_1 _5892_ (.A1(_1280_),
    .A2(_1397_),
    .B1(_1399_),
    .Y(_1400_));
 sky130_fd_sc_hd__and2_1 _5893_ (.A(_1400_),
    .B(_0487_),
    .X(_1401_));
 sky130_fd_sc_hd__a221o_1 _5894_ (.A1(_0645_),
    .A2(_1361_),
    .B1(_1391_),
    .B2(_0670_),
    .C1(_1401_),
    .X(net617));
 sky130_fd_sc_hd__a22o_1 _5895_ (.A1(_1361_),
    .A2(_0766_),
    .B1(_0769_),
    .B2(_1393_),
    .X(_1402_));
 sky130_fd_sc_hd__o22a_1 _5896_ (.A1(net119),
    .A2(_0474_),
    .B1(net55),
    .B2(_0477_),
    .X(_1403_));
 sky130_fd_sc_hd__o221a_4 _5897_ (.A1(net220),
    .A2(_0471_),
    .B1(net157),
    .B2(_0468_),
    .C1(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__inv_2 _5898_ (.A(_1404_),
    .Y(_1405_));
 sky130_fd_sc_hd__nand2_1 _5899_ (.A(_1395_),
    .B(_0767_),
    .Y(_1406_));
 sky130_fd_sc_hd__o21ai_1 _5900_ (.A1(_0855_),
    .A2(_1405_),
    .B1(_1406_),
    .Y(_1407_));
 sky130_fd_sc_hd__mux2_1 _5901_ (.A0(_1402_),
    .A1(_1407_),
    .S(_0886_),
    .X(_1408_));
 sky130_fd_sc_hd__o22a_1 _5902_ (.A1(net117),
    .A2(_0454_),
    .B1(net53),
    .B2(_0456_),
    .X(_1409_));
 sky130_fd_sc_hd__o221a_4 _5903_ (.A1(net155),
    .A2(_0450_),
    .B1(net218),
    .B2(_0452_),
    .C1(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__nand2_1 _5904_ (.A(_1318_),
    .B(_0800_),
    .Y(_1411_));
 sky130_fd_sc_hd__inv_2 _5905_ (.A(_1411_),
    .Y(_1412_));
 sky130_fd_sc_hd__a21oi_1 _5906_ (.A1(_0523_),
    .A2(_1383_),
    .B1(_1412_),
    .Y(_1413_));
 sky130_fd_sc_hd__or3_1 _5907_ (.A(_1007_),
    .B(_0704_),
    .C(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__inv_2 _5908_ (.A(_1382_),
    .Y(_1415_));
 sky130_fd_sc_hd__nand2_1 _5909_ (.A(_1415_),
    .B(_0677_),
    .Y(_1416_));
 sky130_fd_sc_hd__o22a_1 _5910_ (.A1(net119),
    .A2(_0625_),
    .B1(net55),
    .B2(_0626_),
    .X(_1417_));
 sky130_fd_sc_hd__o221a_4 _5911_ (.A1(net220),
    .A2(_0409_),
    .B1(net157),
    .B2(_0408_),
    .C1(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__nand2_1 _5912_ (.A(_1418_),
    .B(_0785_),
    .Y(_1419_));
 sky130_fd_sc_hd__mux2_1 _5913_ (.A0(_1419_),
    .A1(_1368_),
    .S(_0555_),
    .X(_1420_));
 sky130_fd_sc_hd__nand2_1 _5914_ (.A(_1420_),
    .B(_0833_),
    .Y(_1421_));
 sky130_fd_sc_hd__o21ai_1 _5915_ (.A1(_0833_),
    .A2(_1348_),
    .B1(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__a22o_1 _5916_ (.A1(_0417_),
    .A2(_1365_),
    .B1(_1422_),
    .B2(_0419_),
    .X(_1423_));
 sky130_fd_sc_hd__a31o_2 _5917_ (.A1(_0592_),
    .A2(_1414_),
    .A3(_1416_),
    .B1(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__nand2_1 _5918_ (.A(_1424_),
    .B(_0682_),
    .Y(_1425_));
 sky130_fd_sc_hd__o211a_1 _5919_ (.A1(_0682_),
    .A2(_1410_),
    .B1(_0670_),
    .C1(_1425_),
    .X(_1426_));
 sky130_fd_sc_hd__a221o_1 _5920_ (.A1(_0645_),
    .A2(_1393_),
    .B1(_0660_),
    .B2(_1408_),
    .C1(_1426_),
    .X(net618));
 sky130_fd_sc_hd__o22a_1 _5921_ (.A1(net120),
    .A2(_0474_),
    .B1(net57),
    .B2(_0478_),
    .X(_1427_));
 sky130_fd_sc_hd__o221a_4 _5922_ (.A1(net158),
    .A2(_0468_),
    .B1(net221),
    .B2(_0471_),
    .C1(_1427_),
    .X(_1428_));
 sky130_fd_sc_hd__nand2_1 _5923_ (.A(_1428_),
    .B(_0888_),
    .Y(_1429_));
 sky130_fd_sc_hd__nand2_1 _5924_ (.A(_1404_),
    .B(_0888_),
    .Y(_1430_));
 sky130_fd_sc_hd__mux2_1 _5925_ (.A0(_1429_),
    .A1(_1430_),
    .S(_0855_),
    .X(_1431_));
 sky130_fd_sc_hd__nor2_1 _5926_ (.A(_0887_),
    .B(_1396_),
    .Y(_1432_));
 sky130_fd_sc_hd__a21oi_2 _5927_ (.A1(_0887_),
    .A2(_1431_),
    .B1(_1432_),
    .Y(_1433_));
 sky130_fd_sc_hd__o22a_1 _5928_ (.A1(net118),
    .A2(_0724_),
    .B1(net54),
    .B2(_0725_),
    .X(_1434_));
 sky130_fd_sc_hd__o221a_4 _5929_ (.A1(net156),
    .A2(_0637_),
    .B1(net219),
    .B2(_0723_),
    .C1(_1434_),
    .X(_1435_));
 sky130_fd_sc_hd__inv_2 _5930_ (.A(_1377_),
    .Y(_1436_));
 sky130_fd_sc_hd__inv_2 _5931_ (.A(net158),
    .Y(_1437_));
 sky130_fd_sc_hd__inv_2 _5932_ (.A(net221),
    .Y(_1438_));
 sky130_fd_sc_hd__a22oi_1 _5933_ (.A1(_0263_),
    .A2(net120),
    .B1(_0434_),
    .B2(net57),
    .Y(_1439_));
 sky130_fd_sc_hd__o221a_2 _5934_ (.A1(_1437_),
    .A2(_0424_),
    .B1(_1438_),
    .B2(_0429_),
    .C1(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__nor2_1 _5935_ (.A(_4204_),
    .B(_1440_),
    .Y(_1441_));
 sky130_fd_sc_hd__inv_2 _5936_ (.A(net220),
    .Y(_1442_));
 sky130_fd_sc_hd__inv_2 _5937_ (.A(net157),
    .Y(_1443_));
 sky130_fd_sc_hd__a22oi_1 _5938_ (.A1(_0263_),
    .A2(net119),
    .B1(_0434_),
    .B2(net55),
    .Y(_1444_));
 sky130_fd_sc_hd__o221a_2 _5939_ (.A1(_1442_),
    .A2(_0429_),
    .B1(_1443_),
    .B2(_0424_),
    .C1(_1444_),
    .X(_1445_));
 sky130_fd_sc_hd__or3_1 _5940_ (.A(_4127_),
    .B(_4119_),
    .C(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__inv_2 _5941_ (.A(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__a21o_1 _5942_ (.A1(_0522_),
    .A2(_1441_),
    .B1(_1447_),
    .X(_1448_));
 sky130_fd_sc_hd__mux2_1 _5943_ (.A0(_1448_),
    .A1(_1384_),
    .S(_0813_),
    .X(_1449_));
 sky130_fd_sc_hd__a22o_1 _5944_ (.A1(_0677_),
    .A2(_1436_),
    .B1(_1449_),
    .B2(_0443_),
    .X(_1450_));
 sky130_fd_sc_hd__o22a_1 _5945_ (.A1(net120),
    .A2(_0411_),
    .B1(net57),
    .B2(_0413_),
    .X(_1451_));
 sky130_fd_sc_hd__o221a_2 _5946_ (.A1(net158),
    .A2(_0407_),
    .B1(net221),
    .B2(_0409_),
    .C1(_1451_),
    .X(_1452_));
 sky130_fd_sc_hd__nand2_1 _5947_ (.A(_1452_),
    .B(_4272_),
    .Y(_1453_));
 sky130_fd_sc_hd__or2_1 _5948_ (.A(_0557_),
    .B(_1419_),
    .X(_1454_));
 sky130_fd_sc_hd__o21ai_1 _5949_ (.A1(_0555_),
    .A2(_1453_),
    .B1(_1454_),
    .Y(_1455_));
 sky130_fd_sc_hd__nand2_1 _5950_ (.A(_1455_),
    .B(_0833_),
    .Y(_1456_));
 sky130_fd_sc_hd__o21ai_2 _5951_ (.A1(_0833_),
    .A2(_1369_),
    .B1(_1456_),
    .Y(_1457_));
 sky130_fd_sc_hd__a22o_1 _5952_ (.A1(_0417_),
    .A2(_1367_),
    .B1(_1457_),
    .B2(_0419_),
    .X(_1458_));
 sky130_fd_sc_hd__a211o_1 _5953_ (.A1(_1450_),
    .A2(_0592_),
    .B1(_0465_),
    .C1(_1458_),
    .X(_1459_));
 sky130_fd_sc_hd__o211a_1 _5954_ (.A1(_0682_),
    .A2(_1435_),
    .B1(_0601_),
    .C1(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__a221o_1 _5955_ (.A1(_0645_),
    .A2(_1395_),
    .B1(_0660_),
    .B2(_1433_),
    .C1(_1460_),
    .X(net619));
 sky130_fd_sc_hd__o22a_1 _5956_ (.A1(net121),
    .A2(_0475_),
    .B1(net58),
    .B2(_0478_),
    .X(_1461_));
 sky130_fd_sc_hd__o221a_4 _5957_ (.A1(net159),
    .A2(_0468_),
    .B1(net222),
    .B2(_0472_),
    .C1(_1461_),
    .X(_1462_));
 sky130_fd_sc_hd__nand2_1 _5958_ (.A(_1462_),
    .B(_0888_),
    .Y(_1463_));
 sky130_fd_sc_hd__mux2_1 _5959_ (.A0(_1463_),
    .A1(_1429_),
    .S(_0855_),
    .X(_1464_));
 sky130_fd_sc_hd__nor2_1 _5960_ (.A(_0887_),
    .B(_1407_),
    .Y(_1465_));
 sky130_fd_sc_hd__a21oi_2 _5961_ (.A1(_1464_),
    .A2(_0887_),
    .B1(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__o22a_1 _5962_ (.A1(net119),
    .A2(_0724_),
    .B1(net55),
    .B2(_0725_),
    .X(_1467_));
 sky130_fd_sc_hd__o221a_4 _5963_ (.A1(net220),
    .A2(_0723_),
    .B1(net157),
    .B2(_0637_),
    .C1(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__inv_2 _5964_ (.A(_1445_),
    .Y(_1469_));
 sky130_fd_sc_hd__inv_2 _5965_ (.A(net159),
    .Y(_1470_));
 sky130_fd_sc_hd__inv_2 _5966_ (.A(net222),
    .Y(_1471_));
 sky130_fd_sc_hd__a22oi_1 _5967_ (.A1(_0263_),
    .A2(net121),
    .B1(_0434_),
    .B2(net58),
    .Y(_1472_));
 sky130_fd_sc_hd__o221a_2 _5968_ (.A1(_1470_),
    .A2(_0424_),
    .B1(_1471_),
    .B2(_0429_),
    .C1(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__inv_2 _5969_ (.A(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__nand2_1 _5970_ (.A(_1441_),
    .B(_4114_),
    .Y(_1475_));
 sky130_fd_sc_hd__inv_2 _5971_ (.A(_1475_),
    .Y(_1476_));
 sky130_fd_sc_hd__a31o_1 _5972_ (.A1(_1474_),
    .A2(_4127_),
    .A3(_0520_),
    .B1(_1476_),
    .X(_1477_));
 sky130_fd_sc_hd__o21ai_1 _5973_ (.A1(_0538_),
    .A2(_1445_),
    .B1(_0522_),
    .Y(_1478_));
 sky130_fd_sc_hd__o21a_2 _5974_ (.A1(_0522_),
    .A2(_1378_),
    .B1(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__mux2_1 _5975_ (.A0(_1477_),
    .A1(_1479_),
    .S(_0813_),
    .X(_1480_));
 sky130_fd_sc_hd__a22o_1 _5976_ (.A1(_0677_),
    .A2(_1469_),
    .B1(_1480_),
    .B2(_0443_),
    .X(_1481_));
 sky130_fd_sc_hd__o22a_1 _5977_ (.A1(net121),
    .A2(_0625_),
    .B1(net58),
    .B2(_0626_),
    .X(_1482_));
 sky130_fd_sc_hd__o221a_2 _5978_ (.A1(net159),
    .A2(_0408_),
    .B1(net222),
    .B2(_0624_),
    .C1(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__nand2_1 _5979_ (.A(_1483_),
    .B(_0785_),
    .Y(_1484_));
 sky130_fd_sc_hd__or2_1 _5980_ (.A(_0510_),
    .B(_1453_),
    .X(_1485_));
 sky130_fd_sc_hd__o21ai_1 _5981_ (.A1(_0555_),
    .A2(_1484_),
    .B1(_1485_),
    .Y(_1486_));
 sky130_fd_sc_hd__nand2_1 _5982_ (.A(_1486_),
    .B(_0833_),
    .Y(_1487_));
 sky130_fd_sc_hd__o21ai_2 _5983_ (.A1(_0833_),
    .A2(_1420_),
    .B1(_1487_),
    .Y(_1488_));
 sky130_fd_sc_hd__a22o_1 _5984_ (.A1(_0417_),
    .A2(_1418_),
    .B1(_1488_),
    .B2(_0419_),
    .X(_1489_));
 sky130_fd_sc_hd__a211o_1 _5985_ (.A1(_1481_),
    .A2(_0592_),
    .B1(_0465_),
    .C1(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__o211a_1 _5986_ (.A1(_0682_),
    .A2(_1468_),
    .B1(_0601_),
    .C1(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__a221o_1 _5987_ (.A1(_0645_),
    .A2(_1404_),
    .B1(_0660_),
    .B2(_1466_),
    .C1(_1491_),
    .X(net620));
 sky130_fd_sc_hd__inv_2 _5988_ (.A(net160),
    .Y(_1492_));
 sky130_fd_sc_hd__inv_2 _5989_ (.A(net223),
    .Y(_1493_));
 sky130_fd_sc_hd__a22oi_1 _5990_ (.A1(_0803_),
    .A2(net122),
    .B1(_0804_),
    .B2(net59),
    .Y(_1494_));
 sky130_fd_sc_hd__o221a_1 _5991_ (.A1(_1492_),
    .A2(_0425_),
    .B1(_1493_),
    .B2(_0430_),
    .C1(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__nor2_1 _5992_ (.A(_0910_),
    .B(_1495_),
    .Y(_1496_));
 sky130_fd_sc_hd__or3_1 _5993_ (.A(_4127_),
    .B(_4119_),
    .C(_1473_),
    .X(_1497_));
 sky130_fd_sc_hd__inv_2 _5994_ (.A(_1497_),
    .Y(_1498_));
 sky130_fd_sc_hd__a21o_1 _5995_ (.A1(_0522_),
    .A2(_1496_),
    .B1(_1498_),
    .X(_1499_));
 sky130_fd_sc_hd__mux2_1 _5996_ (.A0(_1499_),
    .A1(_1448_),
    .S(_0813_),
    .X(_1500_));
 sky130_fd_sc_hd__nand2_1 _5997_ (.A(_1500_),
    .B(_0706_),
    .Y(_1501_));
 sky130_fd_sc_hd__inv_2 _5998_ (.A(_1440_),
    .Y(_1502_));
 sky130_fd_sc_hd__nand2_1 _5999_ (.A(_1502_),
    .B(_0441_),
    .Y(_1503_));
 sky130_fd_sc_hd__a21o_1 _6000_ (.A1(_1501_),
    .A2(_1503_),
    .B1(_4268_),
    .X(_1504_));
 sky130_fd_sc_hd__nand2_1 _6001_ (.A(_1455_),
    .B(_0719_),
    .Y(_1505_));
 sky130_fd_sc_hd__inv_2 _6002_ (.A(_1452_),
    .Y(_1506_));
 sky130_fd_sc_hd__a21bo_1 _6003_ (.A1(_1503_),
    .A2(_0287_),
    .B1_N(_0550_),
    .X(_1507_));
 sky130_fd_sc_hd__a22o_1 _6004_ (.A1(_0632_),
    .A2(_1506_),
    .B1(_1501_),
    .B2(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__a31o_2 _6005_ (.A1(_1504_),
    .A2(_4233_),
    .A3(_1505_),
    .B1(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__nand2_1 _6006_ (.A(_1509_),
    .B(_0668_),
    .Y(_1510_));
 sky130_fd_sc_hd__o22a_1 _6007_ (.A1(net120),
    .A2(_0454_),
    .B1(net57),
    .B2(_0456_),
    .X(_1511_));
 sky130_fd_sc_hd__o221a_4 _6008_ (.A1(net158),
    .A2(_0450_),
    .B1(net221),
    .B2(_0452_),
    .C1(_1511_),
    .X(_1512_));
 sky130_fd_sc_hd__o21a_1 _6009_ (.A1(_0682_),
    .A2(_1512_),
    .B1(_0670_),
    .X(_1513_));
 sky130_fd_sc_hd__a22o_1 _6010_ (.A1(_0567_),
    .A2(_1428_),
    .B1(_1510_),
    .B2(_1513_),
    .X(net621));
 sky130_fd_sc_hd__o22a_1 _6011_ (.A1(net124),
    .A2(_0625_),
    .B1(net60),
    .B2(_0626_),
    .X(_1514_));
 sky130_fd_sc_hd__o221a_2 _6012_ (.A1(net161),
    .A2(_0408_),
    .B1(net224),
    .B2(_0624_),
    .C1(_1514_),
    .X(_1515_));
 sky130_fd_sc_hd__nand2_1 _6013_ (.A(_1515_),
    .B(_0785_),
    .Y(_1516_));
 sky130_fd_sc_hd__o22a_1 _6014_ (.A1(net122),
    .A2(_0411_),
    .B1(net59),
    .B2(_0413_),
    .X(_1517_));
 sky130_fd_sc_hd__o221a_2 _6015_ (.A1(net160),
    .A2(_0407_),
    .B1(net223),
    .B2(_0409_),
    .C1(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__nand2_1 _6016_ (.A(_1518_),
    .B(_4272_),
    .Y(_1519_));
 sky130_fd_sc_hd__or2_1 _6017_ (.A(_0510_),
    .B(_1519_),
    .X(_1520_));
 sky130_fd_sc_hd__o21ai_1 _6018_ (.A1(_0555_),
    .A2(_1516_),
    .B1(_1520_),
    .Y(_1521_));
 sky130_fd_sc_hd__mux2_1 _6019_ (.A0(_1521_),
    .A1(_1486_),
    .S(_0718_),
    .X(_1522_));
 sky130_fd_sc_hd__inv_2 _6020_ (.A(net161),
    .Y(_1523_));
 sky130_fd_sc_hd__inv_2 _6021_ (.A(net224),
    .Y(_1524_));
 sky130_fd_sc_hd__a22oi_1 _6022_ (.A1(_0263_),
    .A2(net124),
    .B1(_0804_),
    .B2(net60),
    .Y(_1525_));
 sky130_fd_sc_hd__o221a_2 _6023_ (.A1(_1523_),
    .A2(_0424_),
    .B1(_1524_),
    .B2(_0429_),
    .C1(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__nor2_1 _6024_ (.A(_4204_),
    .B(_1526_),
    .Y(_1527_));
 sky130_fd_sc_hd__mux2_1 _6025_ (.A0(_1496_),
    .A1(_1527_),
    .S(_4127_),
    .X(_1528_));
 sky130_fd_sc_hd__mux2_1 _6026_ (.A0(_1477_),
    .A1(_1528_),
    .S(_0703_),
    .X(_1529_));
 sky130_fd_sc_hd__a22o_1 _6027_ (.A1(_0441_),
    .A2(_1474_),
    .B1(_1529_),
    .B2(_0443_),
    .X(_1530_));
 sky130_fd_sc_hd__inv_2 _6028_ (.A(_1483_),
    .Y(_1531_));
 sky130_fd_sc_hd__nor2_1 _6029_ (.A(_0418_),
    .B(_1531_),
    .Y(_1532_));
 sky130_fd_sc_hd__a221o_2 _6030_ (.A1(_0419_),
    .A2(_1522_),
    .B1(_1530_),
    .B2(_0592_),
    .C1(_1532_),
    .X(_1533_));
 sky130_fd_sc_hd__o22a_1 _6031_ (.A1(net121),
    .A2(_0454_),
    .B1(net58),
    .B2(_0456_),
    .X(_1534_));
 sky130_fd_sc_hd__o221a_4 _6032_ (.A1(net159),
    .A2(_0450_),
    .B1(net222),
    .B2(_0452_),
    .C1(_1534_),
    .X(_1535_));
 sky130_fd_sc_hd__mux2_1 _6033_ (.A0(_1533_),
    .A1(_1535_),
    .S(_0465_),
    .X(_1536_));
 sky130_fd_sc_hd__mux2_1 _6034_ (.A0(_1536_),
    .A1(_1462_),
    .S(_0490_),
    .X(_1537_));
 sky130_fd_sc_hd__buf_1 _6035_ (.A(_1537_),
    .X(net622));
 sky130_fd_sc_hd__o22a_1 _6036_ (.A1(net122),
    .A2(_0475_),
    .B1(net59),
    .B2(_0479_),
    .X(_1538_));
 sky130_fd_sc_hd__o221a_4 _6037_ (.A1(net160),
    .A2(_0646_),
    .B1(net223),
    .B2(_0472_),
    .C1(_1538_),
    .X(_1539_));
 sky130_fd_sc_hd__o22a_1 _6038_ (.A1(net125),
    .A2(_0625_),
    .B1(net61),
    .B2(_0626_),
    .X(_1540_));
 sky130_fd_sc_hd__o221a_4 _6039_ (.A1(net163),
    .A2(_0408_),
    .B1(net225),
    .B2(_0624_),
    .C1(_1540_),
    .X(_1541_));
 sky130_fd_sc_hd__nand2_1 _6040_ (.A(_1541_),
    .B(_0785_),
    .Y(_1542_));
 sky130_fd_sc_hd__mux2_2 _6041_ (.A0(_1516_),
    .A1(_1542_),
    .S(_0558_),
    .X(_1543_));
 sky130_fd_sc_hd__or2_1 _6042_ (.A(_0557_),
    .B(_1484_),
    .X(_1544_));
 sky130_fd_sc_hd__o21ai_1 _6043_ (.A1(_0555_),
    .A2(_1519_),
    .B1(_1544_),
    .Y(_1545_));
 sky130_fd_sc_hd__nand2_1 _6044_ (.A(_1545_),
    .B(_0719_),
    .Y(_1546_));
 sky130_fd_sc_hd__o21ai_2 _6045_ (.A1(_0719_),
    .A2(_1543_),
    .B1(_1546_),
    .Y(_1547_));
 sky130_fd_sc_hd__inv_2 _6046_ (.A(_1495_),
    .Y(_1548_));
 sky130_fd_sc_hd__inv_2 _6047_ (.A(net163),
    .Y(_1549_));
 sky130_fd_sc_hd__inv_2 _6048_ (.A(net225),
    .Y(_1550_));
 sky130_fd_sc_hd__a22oi_1 _6049_ (.A1(_0803_),
    .A2(net125),
    .B1(_0804_),
    .B2(net61),
    .Y(_1551_));
 sky130_fd_sc_hd__o221a_2 _6050_ (.A1(_1549_),
    .A2(_0425_),
    .B1(_1550_),
    .B2(_0430_),
    .C1(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__nand2_1 _6051_ (.A(_1527_),
    .B(_0799_),
    .Y(_1553_));
 sky130_fd_sc_hd__o31a_1 _6052_ (.A1(_0799_),
    .A2(_0538_),
    .A3(_1552_),
    .B1(_1553_),
    .X(_1554_));
 sky130_fd_sc_hd__inv_2 _6053_ (.A(_1554_),
    .Y(_1555_));
 sky130_fd_sc_hd__mux2_1 _6054_ (.A0(_1499_),
    .A1(_1555_),
    .S(_0704_),
    .X(_1556_));
 sky130_fd_sc_hd__a22o_1 _6055_ (.A1(_0677_),
    .A2(_1548_),
    .B1(_1556_),
    .B2(_0706_),
    .X(_1557_));
 sky130_fd_sc_hd__a21o_1 _6056_ (.A1(_1518_),
    .A2(_0632_),
    .B1(_0633_),
    .X(_1558_));
 sky130_fd_sc_hd__a221o_2 _6057_ (.A1(_0631_),
    .A2(_1547_),
    .B1(_1557_),
    .B2(_0604_),
    .C1(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__inv_2 _6058_ (.A(_1539_),
    .Y(_1560_));
 sky130_fd_sc_hd__nand2_1 _6059_ (.A(_1462_),
    .B(_0767_),
    .Y(_1561_));
 sky130_fd_sc_hd__o21ai_2 _6060_ (.A1(_0855_),
    .A2(_1560_),
    .B1(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hd__o22a_1 _6061_ (.A1(net122),
    .A2(_0454_),
    .B1(net59),
    .B2(_0456_),
    .X(_1563_));
 sky130_fd_sc_hd__o221a_4 _6062_ (.A1(net160),
    .A2(_0637_),
    .B1(net223),
    .B2(_0452_),
    .C1(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__nand2_1 _6063_ (.A(_1564_),
    .B(_0844_),
    .Y(_1565_));
 sky130_fd_sc_hd__nand2_1 _6064_ (.A(_1565_),
    .B(_0462_),
    .Y(_1566_));
 sky130_fd_sc_hd__o21a_1 _6065_ (.A1(_0461_),
    .A2(_1564_),
    .B1(_0485_),
    .X(_1567_));
 sky130_fd_sc_hd__o211a_1 _6066_ (.A1(_0488_),
    .A2(_1562_),
    .B1(_1566_),
    .C1(_1567_),
    .X(_1568_));
 sky130_fd_sc_hd__a22o_1 _6067_ (.A1(_0490_),
    .A2(_1539_),
    .B1(_1559_),
    .B2(_1568_),
    .X(net623));
 sky130_fd_sc_hd__o22a_1 _6068_ (.A1(net126),
    .A2(_0411_),
    .B1(net62),
    .B2(_0413_),
    .X(_1569_));
 sky130_fd_sc_hd__o221a_2 _6069_ (.A1(net164),
    .A2(_0492_),
    .B1(net226),
    .B2(_0409_),
    .C1(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__nand2_1 _6070_ (.A(_1570_),
    .B(_4272_),
    .Y(_1571_));
 sky130_fd_sc_hd__mux2_1 _6071_ (.A0(_1571_),
    .A1(_1542_),
    .S(_0555_),
    .X(_1572_));
 sky130_fd_sc_hd__nand2_1 _6072_ (.A(_1521_),
    .B(_0718_),
    .Y(_1573_));
 sky130_fd_sc_hd__o21ai_2 _6073_ (.A1(_0719_),
    .A2(_1572_),
    .B1(_1573_),
    .Y(_1574_));
 sky130_fd_sc_hd__inv_2 _6074_ (.A(_1526_),
    .Y(_1575_));
 sky130_fd_sc_hd__inv_2 _6075_ (.A(net164),
    .Y(_1576_));
 sky130_fd_sc_hd__inv_2 _6076_ (.A(net226),
    .Y(_1577_));
 sky130_fd_sc_hd__a22oi_1 _6077_ (.A1(_0803_),
    .A2(net126),
    .B1(_0804_),
    .B2(net62),
    .Y(_1578_));
 sky130_fd_sc_hd__o221a_2 _6078_ (.A1(_1576_),
    .A2(_0425_),
    .B1(_1577_),
    .B2(_0430_),
    .C1(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__nor2_1 _6079_ (.A(_0910_),
    .B(_1579_),
    .Y(_1580_));
 sky130_fd_sc_hd__nor2_1 _6080_ (.A(_0538_),
    .B(_1552_),
    .Y(_1581_));
 sky130_fd_sc_hd__mux2_1 _6081_ (.A0(_1580_),
    .A1(_1581_),
    .S(_0799_),
    .X(_1582_));
 sky130_fd_sc_hd__mux2_1 _6082_ (.A0(_1582_),
    .A1(_1528_),
    .S(_0813_),
    .X(_1583_));
 sky130_fd_sc_hd__a22o_1 _6083_ (.A1(_0441_),
    .A2(_1575_),
    .B1(_1583_),
    .B2(_0443_),
    .X(_1584_));
 sky130_fd_sc_hd__and2_1 _6084_ (.A(_1515_),
    .B(_0417_),
    .X(_1585_));
 sky130_fd_sc_hd__a221o_1 _6085_ (.A1(_0419_),
    .A2(_1574_),
    .B1(_1584_),
    .B2(_0592_),
    .C1(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__o22a_1 _6086_ (.A1(net124),
    .A2(_0724_),
    .B1(net60),
    .B2(_0725_),
    .X(_1587_));
 sky130_fd_sc_hd__o221a_4 _6087_ (.A1(net161),
    .A2(_0637_),
    .B1(net224),
    .B2(_0723_),
    .C1(_1587_),
    .X(_1588_));
 sky130_fd_sc_hd__mux2_2 _6088_ (.A0(_1586_),
    .A1(_1588_),
    .S(_0465_),
    .X(_1589_));
 sky130_fd_sc_hd__o22a_1 _6089_ (.A1(net124),
    .A2(_0186_),
    .B1(net60),
    .B2(_0477_),
    .X(_1590_));
 sky130_fd_sc_hd__o221a_4 _6090_ (.A1(net161),
    .A2(_0467_),
    .B1(net224),
    .B2(_0185_),
    .C1(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__mux2_1 _6091_ (.A0(_1589_),
    .A1(_1591_),
    .S(_0490_),
    .X(_1592_));
 sky130_fd_sc_hd__buf_1 _6092_ (.A(_1592_),
    .X(net625));
 sky130_fd_sc_hd__o22a_1 _6093_ (.A1(net125),
    .A2(_0186_),
    .B1(net61),
    .B2(_0477_),
    .X(_1593_));
 sky130_fd_sc_hd__o221a_4 _6094_ (.A1(net163),
    .A2(_0467_),
    .B1(net225),
    .B2(_0185_),
    .C1(_1593_),
    .X(_1594_));
 sky130_fd_sc_hd__and2_1 _6095_ (.A(_1591_),
    .B(_0766_),
    .X(_1595_));
 sky130_fd_sc_hd__a21o_1 _6096_ (.A1(_0198_),
    .A2(_1594_),
    .B1(_1595_),
    .X(_1596_));
 sky130_fd_sc_hd__o22a_1 _6097_ (.A1(net127),
    .A2(_0123_),
    .B1(net63),
    .B2(_0122_),
    .X(_1597_));
 sky130_fd_sc_hd__o221a_4 _6098_ (.A1(net165),
    .A2(_0449_),
    .B1(net227),
    .B2(_0365_),
    .C1(_1597_),
    .X(_1598_));
 sky130_fd_sc_hd__nand2_1 _6099_ (.A(_1598_),
    .B(_0844_),
    .Y(_1599_));
 sky130_fd_sc_hd__o22a_1 _6100_ (.A1(net126),
    .A2(_0123_),
    .B1(net62),
    .B2(_0122_),
    .X(_1600_));
 sky130_fd_sc_hd__o221a_4 _6101_ (.A1(net164),
    .A2(_0128_),
    .B1(net226),
    .B2(_0365_),
    .C1(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__nand2_1 _6102_ (.A(_1601_),
    .B(_0152_),
    .Y(_1602_));
 sky130_fd_sc_hd__mux2_1 _6103_ (.A0(_1599_),
    .A1(_1602_),
    .S(_0090_),
    .X(_1603_));
 sky130_fd_sc_hd__o22a_1 _6104_ (.A1(net125),
    .A2(_0454_),
    .B1(net61),
    .B2(_0456_),
    .X(_1604_));
 sky130_fd_sc_hd__o221a_4 _6105_ (.A1(net163),
    .A2(_0450_),
    .B1(net225),
    .B2(_0452_),
    .C1(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__nand2_1 _6106_ (.A(_1605_),
    .B(_0844_),
    .Y(_1606_));
 sky130_fd_sc_hd__nand2_1 _6107_ (.A(_1588_),
    .B(_0844_),
    .Y(_1607_));
 sky130_fd_sc_hd__or2_1 _6108_ (.A(_0730_),
    .B(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__o21ai_4 _6109_ (.A1(_0090_),
    .A2(_1606_),
    .B1(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__nand2_1 _6110_ (.A(_1609_),
    .B(_0761_),
    .Y(_1610_));
 sky130_fd_sc_hd__o21ai_2 _6111_ (.A1(_0761_),
    .A2(_1603_),
    .B1(_1610_),
    .Y(_1611_));
 sky130_fd_sc_hd__or2_1 _6112_ (.A(_0461_),
    .B(_1605_),
    .X(_1612_));
 sky130_fd_sc_hd__o22a_1 _6113_ (.A1(net127),
    .A2(_0625_),
    .B1(net63),
    .B2(_0626_),
    .X(_1613_));
 sky130_fd_sc_hd__o221a_4 _6114_ (.A1(net165),
    .A2(_0492_),
    .B1(net227),
    .B2(_0624_),
    .C1(_1613_),
    .X(_1614_));
 sky130_fd_sc_hd__nand2_1 _6115_ (.A(_1614_),
    .B(_0785_),
    .Y(_1615_));
 sky130_fd_sc_hd__or2_1 _6116_ (.A(_0557_),
    .B(_1571_),
    .X(_1616_));
 sky130_fd_sc_hd__o21ai_1 _6117_ (.A1(_0555_),
    .A2(_1615_),
    .B1(_1616_),
    .Y(_1617_));
 sky130_fd_sc_hd__nand2_1 _6118_ (.A(_1617_),
    .B(_0833_),
    .Y(_1618_));
 sky130_fd_sc_hd__o21ai_4 _6119_ (.A1(_0833_),
    .A2(_1543_),
    .B1(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__a22o_1 _6120_ (.A1(_0663_),
    .A2(net165),
    .B1(_0664_),
    .B2(net227),
    .X(_1620_));
 sky130_fd_sc_hd__a221oi_4 _6121_ (.A1(net63),
    .A2(_0435_),
    .B1(net127),
    .B2(_0432_),
    .C1(_1620_),
    .Y(_1621_));
 sky130_fd_sc_hd__nand2_1 _6122_ (.A(_1580_),
    .B(_0800_),
    .Y(_1622_));
 sky130_fd_sc_hd__o21ai_1 _6123_ (.A1(_0800_),
    .A2(_1621_),
    .B1(_1622_),
    .Y(_1623_));
 sky130_fd_sc_hd__mux2_1 _6124_ (.A0(_1555_),
    .A1(_1623_),
    .S(_0703_),
    .X(_1624_));
 sky130_fd_sc_hd__nor2_1 _6125_ (.A(_0591_),
    .B(_1552_),
    .Y(_1625_));
 sky130_fd_sc_hd__a211o_1 _6126_ (.A1(_1624_),
    .A2(_0706_),
    .B1(_0422_),
    .C1(_1625_),
    .X(_1626_));
 sky130_fd_sc_hd__o221ai_4 _6127_ (.A1(_0418_),
    .A2(_1541_),
    .B1(_0420_),
    .B2(_1619_),
    .C1(_1626_),
    .Y(_1627_));
 sky130_fd_sc_hd__nand2_1 _6128_ (.A(_1627_),
    .B(_0682_),
    .Y(_1628_));
 sky130_fd_sc_hd__o2111a_1 _6129_ (.A1(_0463_),
    .A2(_1611_),
    .B1(_0601_),
    .C1(_1612_),
    .D1(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__a221o_1 _6130_ (.A1(_0645_),
    .A2(_1594_),
    .B1(_0660_),
    .B2(_1596_),
    .C1(_1629_),
    .X(net626));
 sky130_fd_sc_hd__o21ai_1 _6131_ (.A1(_0591_),
    .A2(_1579_),
    .B1(_0525_),
    .Y(_1630_));
 sky130_fd_sc_hd__a22o_1 _6132_ (.A1(_0550_),
    .A2(_1630_),
    .B1(_1582_),
    .B2(_0706_),
    .X(_1631_));
 sky130_fd_sc_hd__nand2_1 _6133_ (.A(_1572_),
    .B(_0631_),
    .Y(_1632_));
 sky130_fd_sc_hd__o21a_1 _6134_ (.A1(_0418_),
    .A2(_1570_),
    .B1(_0667_),
    .X(_1633_));
 sky130_fd_sc_hd__a32o_2 _6135_ (.A1(_1631_),
    .A2(_1632_),
    .A3(_1633_),
    .B1(_0535_),
    .B2(_1601_),
    .X(_1634_));
 sky130_fd_sc_hd__o22a_1 _6136_ (.A1(net126),
    .A2(_0474_),
    .B1(net62),
    .B2(_0478_),
    .X(_1635_));
 sky130_fd_sc_hd__o221a_4 _6137_ (.A1(net164),
    .A2(_0468_),
    .B1(net226),
    .B2(_0471_),
    .C1(_1635_),
    .X(_1636_));
 sky130_fd_sc_hd__o22a_1 _6138_ (.A1(net128),
    .A2(_0474_),
    .B1(net64),
    .B2(_0478_),
    .X(_1637_));
 sky130_fd_sc_hd__o221a_4 _6139_ (.A1(net2),
    .A2(_0471_),
    .B1(net166),
    .B2(_0468_),
    .C1(_1637_),
    .X(_1638_));
 sky130_fd_sc_hd__o22a_1 _6140_ (.A1(net127),
    .A2(_0474_),
    .B1(net63),
    .B2(_0478_),
    .X(_1639_));
 sky130_fd_sc_hd__o221a_4 _6141_ (.A1(net165),
    .A2(_0468_),
    .B1(net227),
    .B2(_0471_),
    .C1(_1639_),
    .X(_1640_));
 sky130_fd_sc_hd__a22o_1 _6142_ (.A1(_1638_),
    .A2(_0769_),
    .B1(_0767_),
    .B2(_1640_),
    .X(_1641_));
 sky130_fd_sc_hd__a22o_1 _6143_ (.A1(_1594_),
    .A2(_0767_),
    .B1(_0769_),
    .B2(_1636_),
    .X(_1642_));
 sky130_fd_sc_hd__mux2_1 _6144_ (.A0(_1641_),
    .A1(_1642_),
    .S(_1280_),
    .X(_1643_));
 sky130_fd_sc_hd__a22o_1 _6145_ (.A1(_0645_),
    .A2(_1636_),
    .B1(_1643_),
    .B2(_0660_),
    .X(_1644_));
 sky130_fd_sc_hd__a21o_1 _6146_ (.A1(_1634_),
    .A2(_0636_),
    .B1(_1644_),
    .X(net627));
 sky130_fd_sc_hd__o22a_1 _6147_ (.A1(net129),
    .A2(_0411_),
    .B1(net65),
    .B2(_0413_),
    .X(_1645_));
 sky130_fd_sc_hd__o221a_4 _6148_ (.A1(net167),
    .A2(_0492_),
    .B1(net3),
    .B2(_0409_),
    .C1(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__nand2_1 _6149_ (.A(_1646_),
    .B(_0785_),
    .Y(_1647_));
 sky130_fd_sc_hd__o22a_1 _6150_ (.A1(net128),
    .A2(_0411_),
    .B1(net64),
    .B2(_0413_),
    .X(_1648_));
 sky130_fd_sc_hd__o221a_2 _6151_ (.A1(net2),
    .A2(_0409_),
    .B1(net166),
    .B2(_0492_),
    .C1(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__nand2_1 _6152_ (.A(_1649_),
    .B(_0785_),
    .Y(_1650_));
 sky130_fd_sc_hd__mux2_1 _6153_ (.A0(_1647_),
    .A1(_1650_),
    .S(_4253_),
    .X(_1651_));
 sky130_fd_sc_hd__nand2_1 _6154_ (.A(_1651_),
    .B(_0781_),
    .Y(_1652_));
 sky130_fd_sc_hd__o21ai_1 _6155_ (.A1(_0781_),
    .A2(_1617_),
    .B1(_1652_),
    .Y(_1653_));
 sky130_fd_sc_hd__inv_2 _6156_ (.A(_1653_),
    .Y(_1654_));
 sky130_fd_sc_hd__inv_2 _6157_ (.A(net2),
    .Y(_1655_));
 sky130_fd_sc_hd__inv_2 _6158_ (.A(net166),
    .Y(_1656_));
 sky130_fd_sc_hd__a22oi_1 _6159_ (.A1(_0432_),
    .A2(net128),
    .B1(_0435_),
    .B2(net64),
    .Y(_1657_));
 sky130_fd_sc_hd__o221a_2 _6160_ (.A1(_1655_),
    .A2(_0431_),
    .B1(_1656_),
    .B2(_0426_),
    .C1(_1657_),
    .X(_1658_));
 sky130_fd_sc_hd__nor2_1 _6161_ (.A(_0539_),
    .B(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__a22o_1 _6162_ (.A1(_0663_),
    .A2(net167),
    .B1(_0664_),
    .B2(net3),
    .X(_1660_));
 sky130_fd_sc_hd__a221oi_4 _6163_ (.A1(net65),
    .A2(_0436_),
    .B1(net129),
    .B2(_0432_),
    .C1(_1660_),
    .Y(_1661_));
 sky130_fd_sc_hd__o21ai_1 _6164_ (.A1(_0539_),
    .A2(_1661_),
    .B1(_0522_),
    .Y(_1662_));
 sky130_fd_sc_hd__o21ai_1 _6165_ (.A1(_0522_),
    .A2(_1659_),
    .B1(_1662_),
    .Y(_1663_));
 sky130_fd_sc_hd__nand2_1 _6166_ (.A(_1663_),
    .B(_0703_),
    .Y(_1664_));
 sky130_fd_sc_hd__o21ai_1 _6167_ (.A1(_0703_),
    .A2(_1623_),
    .B1(_1664_),
    .Y(_1665_));
 sky130_fd_sc_hd__o221ai_1 _6168_ (.A1(_0591_),
    .A2(_1621_),
    .B1(_0444_),
    .B2(_1665_),
    .C1(_0592_),
    .Y(_1666_));
 sky130_fd_sc_hd__o221a_1 _6169_ (.A1(_0418_),
    .A2(_1614_),
    .B1(_0420_),
    .B2(_1654_),
    .C1(_1666_),
    .X(_1667_));
 sky130_fd_sc_hd__or2_1 _6170_ (.A(_0535_),
    .B(_1667_),
    .X(_1668_));
 sky130_fd_sc_hd__o22a_1 _6171_ (.A1(net129),
    .A2(_0123_),
    .B1(net65),
    .B2(_0122_),
    .X(_1669_));
 sky130_fd_sc_hd__o221a_4 _6172_ (.A1(net167),
    .A2(_0449_),
    .B1(net3),
    .B2(_0365_),
    .C1(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__nand2_1 _6173_ (.A(_1670_),
    .B(_0844_),
    .Y(_1671_));
 sky130_fd_sc_hd__o22a_1 _6174_ (.A1(net128),
    .A2(_0123_),
    .B1(net64),
    .B2(_0122_),
    .X(_1672_));
 sky130_fd_sc_hd__o221a_4 _6175_ (.A1(net2),
    .A2(_0365_),
    .B1(net166),
    .B2(_0449_),
    .C1(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__nand2_1 _6176_ (.A(_1673_),
    .B(_0844_),
    .Y(_1674_));
 sky130_fd_sc_hd__mux2_1 _6177_ (.A0(_1671_),
    .A1(_1674_),
    .S(_0090_),
    .X(_1675_));
 sky130_fd_sc_hd__mux2_1 _6178_ (.A0(_1603_),
    .A1(_1675_),
    .S(_0841_),
    .X(_1676_));
 sky130_fd_sc_hd__nand2_1 _6179_ (.A(_1676_),
    .B(_0462_),
    .Y(_1677_));
 sky130_fd_sc_hd__inv_2 _6180_ (.A(_1598_),
    .Y(_1678_));
 sky130_fd_sc_hd__nand2_1 _6181_ (.A(_1678_),
    .B(_0460_),
    .Y(_1679_));
 sky130_fd_sc_hd__o22a_1 _6182_ (.A1(net129),
    .A2(_0474_),
    .B1(net65),
    .B2(_0478_),
    .X(_1680_));
 sky130_fd_sc_hd__o221a_4 _6183_ (.A1(net167),
    .A2(_0468_),
    .B1(net3),
    .B2(_0471_),
    .C1(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__nand2_1 _6184_ (.A(_1681_),
    .B(_0888_),
    .Y(_1682_));
 sky130_fd_sc_hd__nand2_1 _6185_ (.A(_1638_),
    .B(_0888_),
    .Y(_1683_));
 sky130_fd_sc_hd__mux2_1 _6186_ (.A0(_1682_),
    .A1(_1683_),
    .S(_0855_),
    .X(_1684_));
 sky130_fd_sc_hd__a22o_1 _6187_ (.A1(_1636_),
    .A2(_0766_),
    .B1(_0769_),
    .B2(_1640_),
    .X(_1685_));
 sky130_fd_sc_hd__nor2_1 _6188_ (.A(_0887_),
    .B(_1685_),
    .Y(_1686_));
 sky130_fd_sc_hd__a21oi_1 _6189_ (.A1(_0887_),
    .A2(_1684_),
    .B1(_1686_),
    .Y(_1687_));
 sky130_fd_sc_hd__a22o_1 _6190_ (.A1(_0484_),
    .A2(_1640_),
    .B1(_1687_),
    .B2(_0660_),
    .X(_1688_));
 sky130_fd_sc_hd__a41o_2 _6191_ (.A1(_1668_),
    .A2(_0636_),
    .A3(_1677_),
    .A4(_1679_),
    .B1(_1688_),
    .X(net628));
 sky130_fd_sc_hd__inv_2 _6192_ (.A(_1649_),
    .Y(_1689_));
 sky130_fd_sc_hd__mux2_1 _6193_ (.A0(_1615_),
    .A1(_1650_),
    .S(_0557_),
    .X(_1690_));
 sky130_fd_sc_hd__o22a_1 _6194_ (.A1(net130),
    .A2(_0625_),
    .B1(net66),
    .B2(_0626_),
    .X(_1691_));
 sky130_fd_sc_hd__o221a_4 _6195_ (.A1(net168),
    .A2(_0408_),
    .B1(net4),
    .B2(_0624_),
    .C1(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__nand2_1 _6196_ (.A(_1692_),
    .B(_0785_),
    .Y(_1693_));
 sky130_fd_sc_hd__mux2_1 _6197_ (.A0(_1647_),
    .A1(_1693_),
    .S(_0557_),
    .X(_1694_));
 sky130_fd_sc_hd__mux2_1 _6198_ (.A0(_1690_),
    .A1(_1694_),
    .S(_0781_),
    .X(_1695_));
 sky130_fd_sc_hd__or4_1 _6199_ (.A(_1007_),
    .B(_0800_),
    .C(_4119_),
    .D(_1658_),
    .X(_1696_));
 sky130_fd_sc_hd__o211a_1 _6200_ (.A1(_0591_),
    .A2(_1658_),
    .B1(_0592_),
    .C1(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__a221o_1 _6201_ (.A1(_0632_),
    .A2(_1689_),
    .B1(_0631_),
    .B2(_1695_),
    .C1(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__nand2_1 _6202_ (.A(_1698_),
    .B(_0668_),
    .Y(_1699_));
 sky130_fd_sc_hd__nand2_1 _6203_ (.A(_1673_),
    .B(_0771_),
    .Y(_1700_));
 sky130_fd_sc_hd__o21ai_1 _6204_ (.A1(_0771_),
    .A2(_1599_),
    .B1(_1700_),
    .Y(_1701_));
 sky130_fd_sc_hd__o22a_1 _6205_ (.A1(net130),
    .A2(_0454_),
    .B1(net66),
    .B2(_0456_),
    .X(_1702_));
 sky130_fd_sc_hd__o221a_4 _6206_ (.A1(net168),
    .A2(_0450_),
    .B1(net4),
    .B2(_0452_),
    .C1(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__nand2_1 _6207_ (.A(_1703_),
    .B(_0844_),
    .Y(_1704_));
 sky130_fd_sc_hd__mux2_1 _6208_ (.A0(_1704_),
    .A1(_1671_),
    .S(_0090_),
    .X(_1705_));
 sky130_fd_sc_hd__nand2_1 _6209_ (.A(_1705_),
    .B(_0841_),
    .Y(_1706_));
 sky130_fd_sc_hd__o21ai_1 _6210_ (.A1(_0841_),
    .A2(_1701_),
    .B1(_1706_),
    .Y(_1707_));
 sky130_fd_sc_hd__nand2_1 _6211_ (.A(_1707_),
    .B(_0462_),
    .Y(_1708_));
 sky130_fd_sc_hd__or2_1 _6212_ (.A(_0461_),
    .B(_1673_),
    .X(_1709_));
 sky130_fd_sc_hd__o22a_1 _6213_ (.A1(net130),
    .A2(_0475_),
    .B1(net66),
    .B2(_0478_),
    .X(_1710_));
 sky130_fd_sc_hd__o221a_4 _6214_ (.A1(net168),
    .A2(_0646_),
    .B1(net4),
    .B2(_0472_),
    .C1(_1710_),
    .X(_1711_));
 sky130_fd_sc_hd__nand2_1 _6215_ (.A(_1711_),
    .B(_0888_),
    .Y(_1712_));
 sky130_fd_sc_hd__mux2_1 _6216_ (.A0(_1712_),
    .A1(_1682_),
    .S(_0855_),
    .X(_1713_));
 sky130_fd_sc_hd__nor2_1 _6217_ (.A(_0887_),
    .B(_1641_),
    .Y(_1714_));
 sky130_fd_sc_hd__a21oi_1 _6218_ (.A1(_0887_),
    .A2(_1713_),
    .B1(_1714_),
    .Y(_1715_));
 sky130_fd_sc_hd__a22o_1 _6219_ (.A1(_0484_),
    .A2(_1638_),
    .B1(_1715_),
    .B2(_0660_),
    .X(_1716_));
 sky130_fd_sc_hd__a41o_2 _6220_ (.A1(_1699_),
    .A2(_0636_),
    .A3(_1708_),
    .A4(_1709_),
    .B1(_1716_),
    .X(net629));
 sky130_fd_sc_hd__inv_2 _6221_ (.A(_1661_),
    .Y(_1717_));
 sky130_fd_sc_hd__a22o_1 _6222_ (.A1(_1646_),
    .A2(_0422_),
    .B1(_1717_),
    .B2(_0447_),
    .X(_1718_));
 sky130_fd_sc_hd__mux2_1 _6223_ (.A0(_1718_),
    .A1(_1670_),
    .S(_0465_),
    .X(_1719_));
 sky130_fd_sc_hd__mux2_1 _6224_ (.A0(_1719_),
    .A1(_1681_),
    .S(_0490_),
    .X(_1720_));
 sky130_fd_sc_hd__buf_1 _6225_ (.A(_1720_),
    .X(net630));
 sky130_fd_sc_hd__inv_2 _6226_ (.A(_1711_),
    .Y(_1721_));
 sky130_fd_sc_hd__inv_2 _6227_ (.A(net168),
    .Y(_1722_));
 sky130_fd_sc_hd__inv_2 _6228_ (.A(net4),
    .Y(_1723_));
 sky130_fd_sc_hd__a22oi_1 _6229_ (.A1(_0433_),
    .A2(net130),
    .B1(_0436_),
    .B2(net66),
    .Y(_1724_));
 sky130_fd_sc_hd__o221a_2 _6230_ (.A1(_1722_),
    .A2(_0426_),
    .B1(_1723_),
    .B2(_0431_),
    .C1(_1724_),
    .X(_1725_));
 sky130_fd_sc_hd__or4_1 _6231_ (.A(_1007_),
    .B(_0800_),
    .C(_4119_),
    .D(_1725_),
    .X(_1726_));
 sky130_fd_sc_hd__o21ai_1 _6232_ (.A1(_0591_),
    .A2(_1725_),
    .B1(_1726_),
    .Y(_1727_));
 sky130_fd_sc_hd__nand2_1 _6233_ (.A(_1727_),
    .B(_0604_),
    .Y(_1728_));
 sky130_fd_sc_hd__nand2_1 _6234_ (.A(_1692_),
    .B(_0422_),
    .Y(_1729_));
 sky130_fd_sc_hd__o21ai_1 _6235_ (.A1(_0682_),
    .A2(_1703_),
    .B1(_0670_),
    .Y(_1730_));
 sky130_fd_sc_hd__a31o_1 _6236_ (.A1(_1728_),
    .A2(_0668_),
    .A3(_1729_),
    .B1(_1730_),
    .X(_1731_));
 sky130_fd_sc_hd__o21ai_2 _6237_ (.A1(_0636_),
    .A2(_1721_),
    .B1(_1731_),
    .Y(net631));
 sky130_fd_sc_hd__o22a_1 _6238_ (.A1(net131),
    .A2(_0454_),
    .B1(net68),
    .B2(_0456_),
    .X(_1732_));
 sky130_fd_sc_hd__o221a_4 _6239_ (.A1(net169),
    .A2(_0450_),
    .B1(net5),
    .B2(_0452_),
    .C1(_1732_),
    .X(_1733_));
 sky130_fd_sc_hd__o22a_1 _6240_ (.A1(net131),
    .A2(_0412_),
    .B1(net68),
    .B2(_0414_),
    .X(_1734_));
 sky130_fd_sc_hd__o221a_2 _6241_ (.A1(net169),
    .A2(_0615_),
    .B1(net5),
    .B2(_0410_),
    .C1(_1734_),
    .X(_1735_));
 sky130_fd_sc_hd__a22o_1 _6242_ (.A1(_0663_),
    .A2(net169),
    .B1(_0664_),
    .B2(net5),
    .X(_1736_));
 sky130_fd_sc_hd__a221oi_1 _6243_ (.A1(net68),
    .A2(_0436_),
    .B1(net131),
    .B2(_0433_),
    .C1(_1736_),
    .Y(_1737_));
 sky130_fd_sc_hd__inv_2 _6244_ (.A(_1737_),
    .Y(_1738_));
 sky130_fd_sc_hd__a221o_1 _6245_ (.A1(_1735_),
    .A2(_0422_),
    .B1(_1738_),
    .B2(_0447_),
    .C1(_0465_),
    .X(_1739_));
 sky130_fd_sc_hd__o21a_1 _6246_ (.A1(_0682_),
    .A2(_1733_),
    .B1(_1739_),
    .X(_1740_));
 sky130_fd_sc_hd__o22a_1 _6247_ (.A1(net131),
    .A2(_0476_),
    .B1(net68),
    .B2(_0480_),
    .X(_1741_));
 sky130_fd_sc_hd__o221a_2 _6248_ (.A1(net169),
    .A2(_0470_),
    .B1(net5),
    .B2(_0473_),
    .C1(_1741_),
    .X(_1742_));
 sky130_fd_sc_hd__mux2_1 _6249_ (.A0(_1740_),
    .A1(_1742_),
    .S(_0489_),
    .X(_1743_));
 sky130_fd_sc_hd__buf_1 _6250_ (.A(_1743_),
    .X(net632));
 sky130_fd_sc_hd__o22a_1 _6251_ (.A1(net132),
    .A2(_0412_),
    .B1(net69),
    .B2(_0414_),
    .X(_1744_));
 sky130_fd_sc_hd__o221a_2 _6252_ (.A1(net170),
    .A2(_0615_),
    .B1(net6),
    .B2(_0410_),
    .C1(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__inv_2 _6253_ (.A(net170),
    .Y(_1746_));
 sky130_fd_sc_hd__inv_2 _6254_ (.A(net6),
    .Y(_1747_));
 sky130_fd_sc_hd__a22oi_1 _6255_ (.A1(_0432_),
    .A2(net132),
    .B1(_0436_),
    .B2(net69),
    .Y(_1748_));
 sky130_fd_sc_hd__o221a_2 _6256_ (.A1(_1746_),
    .A2(_0426_),
    .B1(_1747_),
    .B2(_0431_),
    .C1(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__inv_2 _6257_ (.A(_1749_),
    .Y(_1750_));
 sky130_fd_sc_hd__a221o_1 _6258_ (.A1(_1745_),
    .A2(_0422_),
    .B1(_1750_),
    .B2(_0447_),
    .C1(_0633_),
    .X(_1751_));
 sky130_fd_sc_hd__o22a_1 _6259_ (.A1(net132),
    .A2(_0455_),
    .B1(net69),
    .B2(_0457_),
    .X(_1752_));
 sky130_fd_sc_hd__o221a_2 _6260_ (.A1(net170),
    .A2(_0451_),
    .B1(net6),
    .B2(_0453_),
    .C1(_1752_),
    .X(_1753_));
 sky130_fd_sc_hd__or2_1 _6261_ (.A(_0667_),
    .B(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__o22a_1 _6262_ (.A1(net132),
    .A2(_0475_),
    .B1(net69),
    .B2(_0479_),
    .X(_1755_));
 sky130_fd_sc_hd__o221a_2 _6263_ (.A1(net170),
    .A2(_0469_),
    .B1(net6),
    .B2(_0472_),
    .C1(_1755_),
    .X(_1756_));
 sky130_fd_sc_hd__buf_6 _6264_ (.A(_0168_),
    .X(_1757_));
 sky130_fd_sc_hd__o21ai_1 _6265_ (.A1(_4105_),
    .A2(_1756_),
    .B1(_1757_),
    .Y(_1758_));
 sky130_fd_sc_hd__nand2_4 _6266_ (.A(_0488_),
    .B(_0483_),
    .Y(_1759_));
 sky130_fd_sc_hd__nand2_1 _6267_ (.A(_1758_),
    .B(_1759_),
    .Y(_1760_));
 sky130_fd_sc_hd__a32o_1 _6268_ (.A1(_1751_),
    .A2(_1754_),
    .A3(_1760_),
    .B1(_0490_),
    .B2(_1756_),
    .X(net633));
 sky130_fd_sc_hd__o22a_1 _6269_ (.A1(net133),
    .A2(_0476_),
    .B1(net70),
    .B2(_0479_),
    .X(_1761_));
 sky130_fd_sc_hd__o221a_2 _6270_ (.A1(net171),
    .A2(_0470_),
    .B1(net7),
    .B2(_0472_),
    .C1(_1761_),
    .X(_1762_));
 sky130_fd_sc_hd__a22o_1 _6271_ (.A1(_0663_),
    .A2(net171),
    .B1(_0664_),
    .B2(net7),
    .X(_1763_));
 sky130_fd_sc_hd__a221o_2 _6272_ (.A1(net70),
    .A2(_0436_),
    .B1(net133),
    .B2(_0433_),
    .C1(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__o22a_1 _6273_ (.A1(net133),
    .A2(_0412_),
    .B1(net70),
    .B2(_0414_),
    .X(_1765_));
 sky130_fd_sc_hd__o221a_2 _6274_ (.A1(net171),
    .A2(_0408_),
    .B1(net7),
    .B2(_0410_),
    .C1(_1765_),
    .X(_1766_));
 sky130_fd_sc_hd__o22a_1 _6275_ (.A1(net135),
    .A2(_0036_),
    .B1(net71),
    .B2(_4289_),
    .X(_1767_));
 sky130_fd_sc_hd__o221a_2 _6276_ (.A1(net172),
    .A2(_0407_),
    .B1(net8),
    .B2(_0038_),
    .C1(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__inv_2 _6277_ (.A(_1768_),
    .Y(_1769_));
 sky130_fd_sc_hd__nor2_1 _6278_ (.A(_4278_),
    .B(_1769_),
    .Y(_1770_));
 sky130_fd_sc_hd__o22a_1 _6279_ (.A1(net136),
    .A2(_0412_),
    .B1(net72),
    .B2(_0626_),
    .X(_1771_));
 sky130_fd_sc_hd__o221a_2 _6280_ (.A1(net174),
    .A2(_0408_),
    .B1(net9),
    .B2(_0624_),
    .C1(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__mux2_1 _6281_ (.A0(_1770_),
    .A1(_1772_),
    .S(_0557_),
    .X(_1773_));
 sky130_fd_sc_hd__a22o_1 _6282_ (.A1(_4268_),
    .A2(_1766_),
    .B1(_1773_),
    .B2(_0833_),
    .X(_1774_));
 sky130_fd_sc_hd__inv_2 _6283_ (.A(_1766_),
    .Y(_1775_));
 sky130_fd_sc_hd__nor2_1 _6284_ (.A(_0418_),
    .B(_1775_),
    .Y(_1776_));
 sky130_fd_sc_hd__a221o_1 _6285_ (.A1(_0447_),
    .A2(_1764_),
    .B1(_1774_),
    .B2(_0631_),
    .C1(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__o22a_1 _6286_ (.A1(net133),
    .A2(_0455_),
    .B1(net70),
    .B2(_0457_),
    .X(_1778_));
 sky130_fd_sc_hd__o221a_2 _6287_ (.A1(net171),
    .A2(_0451_),
    .B1(net7),
    .B2(_0453_),
    .C1(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__mux2_1 _6288_ (.A0(_1777_),
    .A1(_1779_),
    .S(_0633_),
    .X(_1780_));
 sky130_fd_sc_hd__o21ai_1 _6289_ (.A1(_4105_),
    .A2(_1762_),
    .B1(_1757_),
    .Y(_1781_));
 sky130_fd_sc_hd__nand2_1 _6290_ (.A(_1781_),
    .B(_1759_),
    .Y(_1782_));
 sky130_fd_sc_hd__a22o_1 _6291_ (.A1(_0490_),
    .A2(_1762_),
    .B1(_1780_),
    .B2(_1782_),
    .X(net634));
 sky130_fd_sc_hd__o22a_1 _6292_ (.A1(net136),
    .A2(_0475_),
    .B1(net72),
    .B2(_0479_),
    .X(_1783_));
 sky130_fd_sc_hd__o221a_4 _6293_ (.A1(net174),
    .A2(_0469_),
    .B1(net9),
    .B2(_0472_),
    .C1(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__o22a_1 _6294_ (.A1(net137),
    .A2(_0475_),
    .B1(net73),
    .B2(_0479_),
    .X(_1785_));
 sky130_fd_sc_hd__o221a_2 _6295_ (.A1(net10),
    .A2(_0472_),
    .B1(net175),
    .B2(_0469_),
    .C1(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__o22a_1 _6296_ (.A1(net135),
    .A2(_0475_),
    .B1(net71),
    .B2(_0479_),
    .X(_1787_));
 sky130_fd_sc_hd__o221a_4 _6297_ (.A1(net172),
    .A2(_0646_),
    .B1(net8),
    .B2(_0472_),
    .C1(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__a221o_1 _6298_ (.A1(_1784_),
    .A2(_0767_),
    .B1(_1786_),
    .B2(_0652_),
    .C1(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__inv_2 _6299_ (.A(net172),
    .Y(_1790_));
 sky130_fd_sc_hd__inv_2 _6300_ (.A(net8),
    .Y(_1791_));
 sky130_fd_sc_hd__a22oi_1 _6301_ (.A1(_0433_),
    .A2(net135),
    .B1(_0436_),
    .B2(net71),
    .Y(_1792_));
 sky130_fd_sc_hd__o221a_2 _6302_ (.A1(_1790_),
    .A2(_0426_),
    .B1(_1791_),
    .B2(_0431_),
    .C1(_1792_),
    .X(_1793_));
 sky130_fd_sc_hd__inv_2 _6303_ (.A(_1793_),
    .Y(_1794_));
 sky130_fd_sc_hd__nor2_1 _6304_ (.A(_0591_),
    .B(_1793_),
    .Y(_1795_));
 sky130_fd_sc_hd__a31o_1 _6305_ (.A1(_1794_),
    .A2(_0589_),
    .A3(_0590_),
    .B1(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__a22o_1 _6306_ (.A1(_0632_),
    .A2(_1768_),
    .B1(_1770_),
    .B2(_0419_),
    .X(_1797_));
 sky130_fd_sc_hd__a211o_1 _6307_ (.A1(_1796_),
    .A2(_0604_),
    .B1(_0633_),
    .C1(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__o21ai_1 _6308_ (.A1(_4105_),
    .A2(_1788_),
    .B1(_0168_),
    .Y(_1799_));
 sky130_fd_sc_hd__o22a_1 _6309_ (.A1(net135),
    .A2(_0455_),
    .B1(net71),
    .B2(_0457_),
    .X(_1800_));
 sky130_fd_sc_hd__o221a_4 _6310_ (.A1(net172),
    .A2(_0451_),
    .B1(net8),
    .B2(_0453_),
    .C1(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__o2bb2a_1 _6311_ (.A1_N(_1759_),
    .A2_N(_1799_),
    .B1(_0667_),
    .B2(_1801_),
    .X(_1802_));
 sky130_fd_sc_hd__nor2_1 _6312_ (.A(_4105_),
    .B(_1799_),
    .Y(_1803_));
 sky130_fd_sc_hd__a221o_1 _6313_ (.A1(_0660_),
    .A2(_1789_),
    .B1(_1798_),
    .B2(_1802_),
    .C1(_1803_),
    .X(net636));
 sky130_fd_sc_hd__nand2_1 _6314_ (.A(_4153_),
    .B(net72),
    .Y(_1804_));
 sky130_fd_sc_hd__nand2_1 _6315_ (.A(\arbiter.master_sel[0][0] ),
    .B(net136),
    .Y(_1805_));
 sky130_fd_sc_hd__a21oi_2 _6316_ (.A1(_1804_),
    .A2(_1805_),
    .B1(_4156_),
    .Y(_1806_));
 sky130_fd_sc_hd__a221o_2 _6317_ (.A1(net174),
    .A2(_0663_),
    .B1(net9),
    .B2(_0664_),
    .C1(_1806_),
    .X(_1807_));
 sky130_fd_sc_hd__o22a_1 _6318_ (.A1(net137),
    .A2(_0412_),
    .B1(net73),
    .B2(_0414_),
    .X(_1808_));
 sky130_fd_sc_hd__o221a_2 _6319_ (.A1(net10),
    .A2(_0410_),
    .B1(net175),
    .B2(_0615_),
    .C1(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__nand2_1 _6320_ (.A(_1809_),
    .B(_0785_),
    .Y(_1810_));
 sky130_fd_sc_hd__nand2_1 _6321_ (.A(_1810_),
    .B(_0555_),
    .Y(_1811_));
 sky130_fd_sc_hd__or2_1 _6322_ (.A(_0781_),
    .B(_1773_),
    .X(_1812_));
 sky130_fd_sc_hd__o2111a_1 _6323_ (.A1(_4271_),
    .A2(_0041_),
    .B1(_1811_),
    .C1(_0419_),
    .D1(_1812_),
    .X(_1813_));
 sky130_fd_sc_hd__a221o_1 _6324_ (.A1(_0632_),
    .A2(_1772_),
    .B1(_0447_),
    .B2(_1807_),
    .C1(_1813_),
    .X(_1814_));
 sky130_fd_sc_hd__o22a_1 _6325_ (.A1(net136),
    .A2(_0455_),
    .B1(net72),
    .B2(_0457_),
    .X(_1815_));
 sky130_fd_sc_hd__o221a_2 _6326_ (.A1(net174),
    .A2(_0451_),
    .B1(net9),
    .B2(_0453_),
    .C1(_1815_),
    .X(_1816_));
 sky130_fd_sc_hd__mux2_1 _6327_ (.A0(_1814_),
    .A1(_1816_),
    .S(_0633_),
    .X(_1817_));
 sky130_fd_sc_hd__o21ai_1 _6328_ (.A1(_4105_),
    .A2(_1784_),
    .B1(_1757_),
    .Y(_1818_));
 sky130_fd_sc_hd__nand2_1 _6329_ (.A(_1818_),
    .B(_1759_),
    .Y(_1819_));
 sky130_fd_sc_hd__a22o_1 _6330_ (.A1(_0490_),
    .A2(_1784_),
    .B1(_1817_),
    .B2(_1819_),
    .X(net637));
 sky130_fd_sc_hd__a22o_1 _6331_ (.A1(_0663_),
    .A2(net175),
    .B1(_0664_),
    .B2(net10),
    .X(_1820_));
 sky130_fd_sc_hd__a221oi_2 _6332_ (.A1(net73),
    .A2(_0436_),
    .B1(net137),
    .B2(_0433_),
    .C1(_1820_),
    .Y(_1821_));
 sky130_fd_sc_hd__inv_2 _6333_ (.A(_1821_),
    .Y(_1822_));
 sky130_fd_sc_hd__a21oi_1 _6334_ (.A1(_1810_),
    .A2(_0719_),
    .B1(_0420_),
    .Y(_1823_));
 sky130_fd_sc_hd__a221o_1 _6335_ (.A1(_1809_),
    .A2(_0417_),
    .B1(_0447_),
    .B2(_1822_),
    .C1(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__o22a_1 _6336_ (.A1(net137),
    .A2(_0455_),
    .B1(net73),
    .B2(_0457_),
    .X(_1825_));
 sky130_fd_sc_hd__o221a_1 _6337_ (.A1(net10),
    .A2(_0453_),
    .B1(net175),
    .B2(_0451_),
    .C1(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__mux2_1 _6338_ (.A0(_1824_),
    .A1(_1826_),
    .S(_0633_),
    .X(_1827_));
 sky130_fd_sc_hd__o21ai_1 _6339_ (.A1(_4105_),
    .A2(_1786_),
    .B1(_1757_),
    .Y(_1828_));
 sky130_fd_sc_hd__nand2_1 _6340_ (.A(_1828_),
    .B(_1759_),
    .Y(_1829_));
 sky130_fd_sc_hd__a22o_1 _6341_ (.A1(_0490_),
    .A2(_1786_),
    .B1(_1827_),
    .B2(_1829_),
    .X(net638));
 sky130_fd_sc_hd__and4_1 _6342_ (.A(_0041_),
    .B(_4233_),
    .C(_0558_),
    .D(\arbiter.slave_sel[1][1] ),
    .X(_1830_));
 sky130_fd_sc_hd__a221o_1 _6343_ (.A1(_0229_),
    .A2(_0447_),
    .B1(_0041_),
    .B2(_0632_),
    .C1(_0633_),
    .X(_1831_));
 sky130_fd_sc_hd__o21ai_1 _6344_ (.A1(_4105_),
    .A2(_0191_),
    .B1(_1757_),
    .Y(_1832_));
 sky130_fd_sc_hd__nand2_1 _6345_ (.A(_1832_),
    .B(_1759_),
    .Y(_1833_));
 sky130_fd_sc_hd__o221a_1 _6346_ (.A1(_0131_),
    .A2(_0682_),
    .B1(_1830_),
    .B2(_1831_),
    .C1(_1833_),
    .X(_1834_));
 sky130_fd_sc_hd__a21o_1 _6347_ (.A1(_0191_),
    .A2(_0567_),
    .B1(_1834_),
    .X(net639));
 sky130_fd_sc_hd__o22a_1 _6348_ (.A1(net139),
    .A2(_0412_),
    .B1(net75),
    .B2(_0414_),
    .X(_1835_));
 sky130_fd_sc_hd__o221a_2 _6349_ (.A1(net177),
    .A2(_0615_),
    .B1(net13),
    .B2(_0410_),
    .C1(_1835_),
    .X(_1836_));
 sky130_fd_sc_hd__a22o_1 _6350_ (.A1(_0663_),
    .A2(net177),
    .B1(_0664_),
    .B2(net13),
    .X(_1837_));
 sky130_fd_sc_hd__a221oi_1 _6351_ (.A1(net75),
    .A2(_0436_),
    .B1(net139),
    .B2(_0433_),
    .C1(_1837_),
    .Y(_1838_));
 sky130_fd_sc_hd__inv_2 _6352_ (.A(_1838_),
    .Y(_1839_));
 sky130_fd_sc_hd__a22o_1 _6353_ (.A1(_1836_),
    .A2(_0422_),
    .B1(_1839_),
    .B2(_0447_),
    .X(_1840_));
 sky130_fd_sc_hd__o22a_1 _6354_ (.A1(net139),
    .A2(_0455_),
    .B1(net75),
    .B2(_0457_),
    .X(_1841_));
 sky130_fd_sc_hd__o221a_2 _6355_ (.A1(net177),
    .A2(_0451_),
    .B1(net13),
    .B2(_0453_),
    .C1(_1841_),
    .X(_1842_));
 sky130_fd_sc_hd__mux2_1 _6356_ (.A0(_1840_),
    .A1(_1842_),
    .S(_0465_),
    .X(_1843_));
 sky130_fd_sc_hd__o22a_1 _6357_ (.A1(net139),
    .A2(_0476_),
    .B1(net75),
    .B2(_0480_),
    .X(_1844_));
 sky130_fd_sc_hd__o221a_2 _6358_ (.A1(net177),
    .A2(_0470_),
    .B1(net13),
    .B2(_0473_),
    .C1(_1844_),
    .X(_1845_));
 sky130_fd_sc_hd__mux2_1 _6359_ (.A0(_1843_),
    .A1(_1845_),
    .S(_0489_),
    .X(_1846_));
 sky130_fd_sc_hd__buf_1 _6360_ (.A(_1846_),
    .X(net640));
 sky130_fd_sc_hd__o22a_1 _6361_ (.A1(net140),
    .A2(_0475_),
    .B1(net76),
    .B2(_0479_),
    .X(_1847_));
 sky130_fd_sc_hd__o221a_2 _6362_ (.A1(net178),
    .A2(_0469_),
    .B1(net14),
    .B2(_0472_),
    .C1(_1847_),
    .X(_1848_));
 sky130_fd_sc_hd__o22a_1 _6363_ (.A1(net140),
    .A2(_0455_),
    .B1(net76),
    .B2(_0457_),
    .X(_1849_));
 sky130_fd_sc_hd__o221a_1 _6364_ (.A1(net178),
    .A2(_0451_),
    .B1(net14),
    .B2(_0453_),
    .C1(_1849_),
    .X(_1850_));
 sky130_fd_sc_hd__a22o_1 _6365_ (.A1(_0663_),
    .A2(net178),
    .B1(_0664_),
    .B2(net14),
    .X(_1851_));
 sky130_fd_sc_hd__a221oi_4 _6366_ (.A1(net76),
    .A2(_0436_),
    .B1(net140),
    .B2(_0433_),
    .C1(_1851_),
    .Y(_1852_));
 sky130_fd_sc_hd__nor2_1 _6367_ (.A(_0446_),
    .B(_1852_),
    .Y(_1853_));
 sky130_fd_sc_hd__o22a_1 _6368_ (.A1(net140),
    .A2(_0412_),
    .B1(net76),
    .B2(_0414_),
    .X(_1854_));
 sky130_fd_sc_hd__o221a_2 _6369_ (.A1(net178),
    .A2(_0615_),
    .B1(net14),
    .B2(_0410_),
    .C1(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__a22o_1 _6370_ (.A1(_1836_),
    .A2(_0613_),
    .B1(_0558_),
    .B2(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__o21a_1 _6371_ (.A1(_0418_),
    .A2(_1855_),
    .B1(_0667_),
    .X(_1857_));
 sky130_fd_sc_hd__o221a_1 _6372_ (.A1(_0422_),
    .A2(_1853_),
    .B1(_0420_),
    .B2(_1856_),
    .C1(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__a21o_1 _6373_ (.A1(_0535_),
    .A2(_1850_),
    .B1(_1858_),
    .X(_1859_));
 sky130_fd_sc_hd__o21ai_1 _6374_ (.A1(_4105_),
    .A2(_1848_),
    .B1(_1757_),
    .Y(_1860_));
 sky130_fd_sc_hd__nand2_1 _6375_ (.A(_1860_),
    .B(_1759_),
    .Y(_1861_));
 sky130_fd_sc_hd__a22o_1 _6376_ (.A1(_0490_),
    .A2(_1848_),
    .B1(_1859_),
    .B2(_1861_),
    .X(net641));
 sky130_fd_sc_hd__o22a_1 _6377_ (.A1(net141),
    .A2(_0412_),
    .B1(net77),
    .B2(_0414_),
    .X(_1862_));
 sky130_fd_sc_hd__o221a_1 _6378_ (.A1(net179),
    .A2(_0615_),
    .B1(net15),
    .B2(_0410_),
    .C1(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__inv_2 _6379_ (.A(_1863_),
    .Y(_1864_));
 sky130_fd_sc_hd__a22o_1 _6380_ (.A1(_0433_),
    .A2(net141),
    .B1(_0436_),
    .B2(net77),
    .X(_1865_));
 sky130_fd_sc_hd__a221oi_4 _6381_ (.A1(net179),
    .A2(_0663_),
    .B1(net15),
    .B2(_0664_),
    .C1(_1865_),
    .Y(_1866_));
 sky130_fd_sc_hd__o22a_1 _6382_ (.A1(_0592_),
    .A2(_1864_),
    .B1(_0662_),
    .B2(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__o22a_1 _6383_ (.A1(net141),
    .A2(_0455_),
    .B1(net77),
    .B2(_0457_),
    .X(_1868_));
 sky130_fd_sc_hd__o221a_2 _6384_ (.A1(net179),
    .A2(_0451_),
    .B1(net15),
    .B2(_0453_),
    .C1(_1868_),
    .X(_1869_));
 sky130_fd_sc_hd__inv_2 _6385_ (.A(_1869_),
    .Y(_1870_));
 sky130_fd_sc_hd__mux2_1 _6386_ (.A0(_1867_),
    .A1(_1870_),
    .S(_0633_),
    .X(_1871_));
 sky130_fd_sc_hd__o22a_1 _6387_ (.A1(net141),
    .A2(_0476_),
    .B1(net77),
    .B2(_0480_),
    .X(_1872_));
 sky130_fd_sc_hd__o221a_2 _6388_ (.A1(net179),
    .A2(_0470_),
    .B1(net15),
    .B2(_0473_),
    .C1(_1872_),
    .X(_1873_));
 sky130_fd_sc_hd__nor2_1 _6389_ (.A(_0636_),
    .B(_1873_),
    .Y(_1874_));
 sky130_fd_sc_hd__a21oi_2 _6390_ (.A1(_1871_),
    .A2(_0636_),
    .B1(_1874_),
    .Y(net642));
 sky130_fd_sc_hd__o22a_1 _6391_ (.A1(net142),
    .A2(_0455_),
    .B1(net79),
    .B2(_0457_),
    .X(_1875_));
 sky130_fd_sc_hd__o221a_2 _6392_ (.A1(net180),
    .A2(_0451_),
    .B1(net16),
    .B2(_0453_),
    .C1(_1875_),
    .X(_1876_));
 sky130_fd_sc_hd__o22a_1 _6393_ (.A1(net142),
    .A2(_0412_),
    .B1(net79),
    .B2(_0414_),
    .X(_1877_));
 sky130_fd_sc_hd__o221a_2 _6394_ (.A1(net180),
    .A2(_0615_),
    .B1(net16),
    .B2(_0410_),
    .C1(_1877_),
    .X(_1878_));
 sky130_fd_sc_hd__and2_1 _6395_ (.A(_1878_),
    .B(_0288_),
    .X(_1879_));
 sky130_fd_sc_hd__a22o_1 _6396_ (.A1(_0663_),
    .A2(net180),
    .B1(_0664_),
    .B2(net16),
    .X(_1880_));
 sky130_fd_sc_hd__a221o_2 _6397_ (.A1(net79),
    .A2(_0436_),
    .B1(net142),
    .B2(_0433_),
    .C1(_1880_),
    .X(_1881_));
 sky130_fd_sc_hd__a221o_1 _6398_ (.A1(_1879_),
    .A2(_0422_),
    .B1(_1881_),
    .B2(_0447_),
    .C1(_0633_),
    .X(_1882_));
 sky130_fd_sc_hd__o21ai_1 _6399_ (.A1(_0668_),
    .A2(_1876_),
    .B1(_1882_),
    .Y(_1883_));
 sky130_fd_sc_hd__o22a_1 _6400_ (.A1(net142),
    .A2(_0476_),
    .B1(net79),
    .B2(_0480_),
    .X(_1884_));
 sky130_fd_sc_hd__o221a_2 _6401_ (.A1(net180),
    .A2(_0470_),
    .B1(net16),
    .B2(_0473_),
    .C1(_1884_),
    .X(_1885_));
 sky130_fd_sc_hd__nor2_1 _6402_ (.A(_0636_),
    .B(_1885_),
    .Y(_1886_));
 sky130_fd_sc_hd__a21oi_2 _6403_ (.A1(_1883_),
    .A2(_0636_),
    .B1(_1886_),
    .Y(net643));
 sky130_fd_sc_hd__nor2_4 _6404_ (.A(_4100_),
    .B(_0056_),
    .Y(_1887_));
 sky130_fd_sc_hd__inv_2 _6405_ (.A(_1887_),
    .Y(_1888_));
 sky130_fd_sc_hd__nand2_8 _6406_ (.A(_4280_),
    .B(_4233_),
    .Y(_1889_));
 sky130_fd_sc_hd__nand2_2 _6407_ (.A(_1888_),
    .B(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__buf_8 _6408_ (.A(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__nor2_8 _6409_ (.A(_4100_),
    .B(_0440_),
    .Y(_1892_));
 sky130_fd_sc_hd__inv_2 _6410_ (.A(_1892_),
    .Y(_1893_));
 sky130_fd_sc_hd__buf_12 _6411_ (.A(_4213_),
    .X(_1894_));
 sky130_fd_sc_hd__nand2_8 _6412_ (.A(_1894_),
    .B(_0588_),
    .Y(_1895_));
 sky130_fd_sc_hd__nand2_2 _6413_ (.A(_1893_),
    .B(_1895_),
    .Y(_1896_));
 sky130_fd_sc_hd__inv_2 _6414_ (.A(_1896_),
    .Y(_1897_));
 sky130_fd_sc_hd__nor2_4 _6415_ (.A(_1890_),
    .B(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__a22o_1 _6416_ (.A1(_0416_),
    .A2(_1891_),
    .B1(_0439_),
    .B2(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__nor2_8 _6417_ (.A(_4100_),
    .B(_0134_),
    .Y(_1900_));
 sky130_fd_sc_hd__inv_2 _6418_ (.A(_1900_),
    .Y(_1901_));
 sky130_fd_sc_hd__nand2_4 _6419_ (.A(_0143_),
    .B(_4239_),
    .Y(_1902_));
 sky130_fd_sc_hd__nand2_2 _6420_ (.A(_1901_),
    .B(_1902_),
    .Y(_1903_));
 sky130_fd_sc_hd__buf_6 _6421_ (.A(_1903_),
    .X(_1904_));
 sky130_fd_sc_hd__mux2_1 _6422_ (.A0(_1899_),
    .A1(_0459_),
    .S(_1904_),
    .X(_1905_));
 sky130_fd_sc_hd__nor2_8 _6423_ (.A(_4100_),
    .B(_0483_),
    .Y(_1906_));
 sky130_fd_sc_hd__inv_2 _6424_ (.A(_1906_),
    .Y(_1907_));
 sky130_fd_sc_hd__nand2_8 _6425_ (.A(_0652_),
    .B(_0209_),
    .Y(_1908_));
 sky130_fd_sc_hd__nand2_1 _6426_ (.A(_1907_),
    .B(_1908_),
    .Y(_1909_));
 sky130_fd_sc_hd__buf_8 _6427_ (.A(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__buf_6 _6428_ (.A(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__mux2_2 _6429_ (.A0(_1905_),
    .A1(_0482_),
    .S(_1911_),
    .X(_1912_));
 sky130_fd_sc_hd__buf_1 _6430_ (.A(_1912_),
    .X(net682));
 sky130_fd_sc_hd__nand2_1 _6431_ (.A(_1889_),
    .B(_0056_),
    .Y(_1913_));
 sky130_fd_sc_hd__buf_6 _6432_ (.A(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__a21o_1 _6433_ (.A1(_0499_),
    .A2(_1896_),
    .B1(_1914_),
    .X(_1915_));
 sky130_fd_sc_hd__nand2_1 _6434_ (.A(_4235_),
    .B(_4100_),
    .Y(_1916_));
 sky130_fd_sc_hd__buf_6 _6435_ (.A(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__inv_2 _6436_ (.A(_1917_),
    .Y(_1918_));
 sky130_fd_sc_hd__o21ai_1 _6437_ (.A1(_1895_),
    .A2(_0498_),
    .B1(_1918_),
    .Y(_1919_));
 sky130_fd_sc_hd__buf_8 _6438_ (.A(_1888_),
    .X(_1920_));
 sky130_fd_sc_hd__or2_1 _6439_ (.A(_1920_),
    .B(_0494_),
    .X(_1921_));
 sky130_fd_sc_hd__nand2_1 _6440_ (.A(_0494_),
    .B(_4272_),
    .Y(_1922_));
 sky130_fd_sc_hd__inv_6 _6441_ (.A(_1889_),
    .Y(_1923_));
 sky130_fd_sc_hd__buf_6 _6442_ (.A(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__nand2_1 _6443_ (.A(_1922_),
    .B(_1924_),
    .Y(_1925_));
 sky130_fd_sc_hd__buf_6 _6444_ (.A(_1903_),
    .X(_1926_));
 sky130_fd_sc_hd__a41o_1 _6445_ (.A1(_1915_),
    .A2(_1919_),
    .A3(_1921_),
    .A4(_1925_),
    .B1(_1926_),
    .X(_1927_));
 sky130_fd_sc_hd__inv_2 _6446_ (.A(_1903_),
    .Y(_1928_));
 sky130_fd_sc_hd__clkbuf_8 _6447_ (.A(_1928_),
    .X(_1929_));
 sky130_fd_sc_hd__inv_2 _6448_ (.A(_1909_),
    .Y(_1930_));
 sky130_fd_sc_hd__buf_8 _6449_ (.A(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__clkbuf_8 _6450_ (.A(_1931_),
    .X(_1932_));
 sky130_fd_sc_hd__o21a_1 _6451_ (.A1(_1929_),
    .A2(_0502_),
    .B1(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__a22o_2 _6452_ (.A1(_0505_),
    .A2(_1911_),
    .B1(_1927_),
    .B2(_1933_),
    .X(net683));
 sky130_fd_sc_hd__a21bo_1 _6453_ (.A1(_0555_),
    .A2(_1922_),
    .B1_N(_0511_),
    .X(_1934_));
 sky130_fd_sc_hd__a31o_1 _6454_ (.A1(_0416_),
    .A2(_0558_),
    .A3(_0785_),
    .B1(_0781_),
    .X(_1935_));
 sky130_fd_sc_hd__a21boi_1 _6455_ (.A1(_1934_),
    .A2(_0833_),
    .B1_N(_1935_),
    .Y(_1936_));
 sky130_fd_sc_hd__nand2_1 _6456_ (.A(_0499_),
    .B(_0520_),
    .Y(_1937_));
 sky130_fd_sc_hd__nand2_1 _6457_ (.A(_1937_),
    .B(_0800_),
    .Y(_1938_));
 sky130_fd_sc_hd__inv_2 _6458_ (.A(_1895_),
    .Y(_1939_));
 sky130_fd_sc_hd__a32o_1 _6459_ (.A1(_1938_),
    .A2(_0524_),
    .A3(_1939_),
    .B1(_0519_),
    .B2(_1892_),
    .X(_1940_));
 sky130_fd_sc_hd__inv_6 _6460_ (.A(_1891_),
    .Y(_1941_));
 sky130_fd_sc_hd__inv_2 _6461_ (.A(_0508_),
    .Y(_1942_));
 sky130_fd_sc_hd__nor2_1 _6462_ (.A(_1888_),
    .B(_1942_),
    .Y(_1943_));
 sky130_fd_sc_hd__a221o_1 _6463_ (.A1(_1936_),
    .A2(_1923_),
    .B1(_1940_),
    .B2(_1941_),
    .C1(_1943_),
    .X(_1944_));
 sky130_fd_sc_hd__mux2_1 _6464_ (.A0(_1944_),
    .A1(_0530_),
    .S(_1904_),
    .X(_1945_));
 sky130_fd_sc_hd__mux2_2 _6465_ (.A0(_1945_),
    .A1(_0533_),
    .S(_1910_),
    .X(_1946_));
 sky130_fd_sc_hd__buf_1 _6466_ (.A(_1946_),
    .X(net684));
 sky130_fd_sc_hd__buf_8 _6467_ (.A(_1928_),
    .X(_1947_));
 sky130_fd_sc_hd__a221o_1 _6468_ (.A1(_0553_),
    .A2(_1887_),
    .B1(_0560_),
    .B2(_1923_),
    .C1(_1926_),
    .X(_1948_));
 sky130_fd_sc_hd__or2_1 _6469_ (.A(_0862_),
    .B(_0546_),
    .X(_1949_));
 sky130_fd_sc_hd__nand2_1 _6470_ (.A(_1937_),
    .B(_0523_),
    .Y(_1950_));
 sky130_fd_sc_hd__o21ai_1 _6471_ (.A1(_4119_),
    .A2(_0438_),
    .B1(_0800_),
    .Y(_1951_));
 sky130_fd_sc_hd__a21o_1 _6472_ (.A1(_1950_),
    .A2(_1951_),
    .B1(_0704_),
    .X(_1952_));
 sky130_fd_sc_hd__clkbuf_8 _6473_ (.A(_1939_),
    .X(_1953_));
 sky130_fd_sc_hd__inv_2 _6474_ (.A(_0543_),
    .Y(_1954_));
 sky130_fd_sc_hd__buf_6 _6475_ (.A(_1892_),
    .X(_1955_));
 sky130_fd_sc_hd__a32o_1 _6476_ (.A1(_1949_),
    .A2(_1952_),
    .A3(_1953_),
    .B1(_1954_),
    .B2(_1955_),
    .X(_1956_));
 sky130_fd_sc_hd__and2_1 _6477_ (.A(_1956_),
    .B(_1941_),
    .X(_1957_));
 sky130_fd_sc_hd__o221a_1 _6478_ (.A1(_0537_),
    .A2(_1947_),
    .B1(_1948_),
    .B2(_1957_),
    .C1(_1932_),
    .X(_1958_));
 sky130_fd_sc_hd__a21o_2 _6479_ (.A1(_0565_),
    .A2(_1911_),
    .B1(_1958_),
    .X(net686));
 sky130_fd_sc_hd__a22o_1 _6480_ (.A1(_0586_),
    .A2(_1892_),
    .B1(_0587_),
    .B2(_1953_),
    .X(_1959_));
 sky130_fd_sc_hd__nand2_1 _6481_ (.A(_1934_),
    .B(_0718_),
    .Y(_1960_));
 sky130_fd_sc_hd__o21ai_1 _6482_ (.A1(_0718_),
    .A2(_0597_),
    .B1(_1960_),
    .Y(_1961_));
 sky130_fd_sc_hd__a2bb2o_1 _6483_ (.A1_N(_1889_),
    .A2_N(_1961_),
    .B1(_0581_),
    .B2(_1887_),
    .X(_1962_));
 sky130_fd_sc_hd__a21o_1 _6484_ (.A1(_1941_),
    .A2(_1959_),
    .B1(_1962_),
    .X(_1963_));
 sky130_fd_sc_hd__mux2_1 _6485_ (.A0(_1963_),
    .A1(_0571_),
    .S(_1904_),
    .X(_1964_));
 sky130_fd_sc_hd__mux2_4 _6486_ (.A0(_1964_),
    .A1(_0569_),
    .S(_1910_),
    .X(_1965_));
 sky130_fd_sc_hd__buf_1 _6487_ (.A(_1965_),
    .X(net687));
 sky130_fd_sc_hd__nand2_1 _6488_ (.A(_0609_),
    .B(_1896_),
    .Y(_1966_));
 sky130_fd_sc_hd__inv_2 _6489_ (.A(_0621_),
    .Y(_1967_));
 sky130_fd_sc_hd__mux2_1 _6490_ (.A0(_1966_),
    .A1(_1967_),
    .S(_1891_),
    .X(_1968_));
 sky130_fd_sc_hd__nand2_1 _6491_ (.A(_1968_),
    .B(_1929_),
    .Y(_1969_));
 sky130_fd_sc_hd__o21a_1 _6492_ (.A1(_1929_),
    .A2(_0574_),
    .B1(_1931_),
    .X(_1970_));
 sky130_fd_sc_hd__a22o_2 _6493_ (.A1(_0648_),
    .A2(_1911_),
    .B1(_1969_),
    .B2(_1970_),
    .X(net688));
 sky130_fd_sc_hd__inv_2 _6494_ (.A(_1894_),
    .Y(_1971_));
 sky130_fd_sc_hd__or3_1 _6495_ (.A(_1007_),
    .B(_1971_),
    .C(net730),
    .X(_1972_));
 sky130_fd_sc_hd__buf_6 _6496_ (.A(_1893_),
    .X(_1973_));
 sky130_fd_sc_hd__nor2_1 _6497_ (.A(_1973_),
    .B(net730),
    .Y(_1974_));
 sky130_fd_sc_hd__o21ai_1 _6498_ (.A1(_1914_),
    .A2(_1974_),
    .B1(_1917_),
    .Y(_1975_));
 sky130_fd_sc_hd__inv_2 _6499_ (.A(_0617_),
    .Y(_1976_));
 sky130_fd_sc_hd__buf_12 _6500_ (.A(_4280_),
    .X(_1977_));
 sky130_fd_sc_hd__a221o_1 _6501_ (.A1(_1977_),
    .A2(_1976_),
    .B1(_0597_),
    .B2(_4268_),
    .C1(_1889_),
    .X(_1978_));
 sky130_fd_sc_hd__o21ai_1 _6502_ (.A1(_1976_),
    .A2(_1920_),
    .B1(_1978_),
    .Y(_1979_));
 sky130_fd_sc_hd__a21o_1 _6503_ (.A1(_1972_),
    .A2(_1975_),
    .B1(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__buf_6 _6504_ (.A(_1902_),
    .X(_1981_));
 sky130_fd_sc_hd__nor2_1 _6505_ (.A(_1981_),
    .B(_0579_),
    .Y(_1982_));
 sky130_fd_sc_hd__buf_8 _6506_ (.A(_1901_),
    .X(_1983_));
 sky130_fd_sc_hd__nor2_1 _6507_ (.A(_1983_),
    .B(_0576_),
    .Y(_1984_));
 sky130_fd_sc_hd__a2111o_1 _6508_ (.A1(_1980_),
    .A2(_1947_),
    .B1(_1910_),
    .C1(_1982_),
    .D1(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__o21ai_2 _6509_ (.A1(_0657_),
    .A2(_1932_),
    .B1(_1985_),
    .Y(net689));
 sky130_fd_sc_hd__clkbuf_8 _6510_ (.A(_1906_),
    .X(_1986_));
 sky130_fd_sc_hd__inv_2 _6511_ (.A(_1908_),
    .Y(_1987_));
 sky130_fd_sc_hd__clkbuf_8 _6512_ (.A(_1987_),
    .X(_1988_));
 sky130_fd_sc_hd__buf_12 _6513_ (.A(_1894_),
    .X(_1989_));
 sky130_fd_sc_hd__nor2_1 _6514_ (.A(_1973_),
    .B(_0675_),
    .Y(_1990_));
 sky130_fd_sc_hd__a31o_1 _6515_ (.A1(_0676_),
    .A2(_0588_),
    .A3(_1989_),
    .B1(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__nand2_1 _6516_ (.A(_1991_),
    .B(_1941_),
    .Y(_1992_));
 sky130_fd_sc_hd__nand2_1 _6517_ (.A(_1992_),
    .B(_1928_),
    .Y(_1993_));
 sky130_fd_sc_hd__a2bb2o_1 _6518_ (.A1_N(_1889_),
    .A2_N(_0623_),
    .B1(_0683_),
    .B2(_1887_),
    .X(_1994_));
 sky130_fd_sc_hd__o21a_1 _6519_ (.A1(_1901_),
    .A2(_0639_),
    .B1(_1930_),
    .X(_1995_));
 sky130_fd_sc_hd__o221a_1 _6520_ (.A1(_0642_),
    .A2(_1981_),
    .B1(_1993_),
    .B2(_1994_),
    .C1(_1995_),
    .X(_1996_));
 sky130_fd_sc_hd__a221o_1 _6521_ (.A1(_0650_),
    .A2(_1986_),
    .B1(_0659_),
    .B2(_1988_),
    .C1(_1996_),
    .X(net690));
 sky130_fd_sc_hd__buf_6 _6522_ (.A(_1953_),
    .X(_1997_));
 sky130_fd_sc_hd__a22o_1 _6523_ (.A1(_0693_),
    .A2(_1955_),
    .B1(_0695_),
    .B2(_1997_),
    .X(_1998_));
 sky130_fd_sc_hd__buf_6 _6524_ (.A(_1941_),
    .X(_1999_));
 sky130_fd_sc_hd__nand2_1 _6525_ (.A(_1998_),
    .B(_1999_),
    .Y(_2000_));
 sky130_fd_sc_hd__inv_2 _6526_ (.A(_0715_),
    .Y(_2001_));
 sky130_fd_sc_hd__o2bb2a_1 _6527_ (.A1_N(_1924_),
    .A2_N(_0716_),
    .B1(_2001_),
    .B2(_1920_),
    .X(_2002_));
 sky130_fd_sc_hd__inv_2 _6528_ (.A(_1902_),
    .Y(_2003_));
 sky130_fd_sc_hd__clkbuf_8 _6529_ (.A(_2003_),
    .X(_2004_));
 sky130_fd_sc_hd__a221o_1 _6530_ (.A1(_0728_),
    .A2(_1900_),
    .B1(_0732_),
    .B2(_2004_),
    .C1(_1910_),
    .X(_2005_));
 sky130_fd_sc_hd__a31o_1 _6531_ (.A1(_2000_),
    .A2(_1929_),
    .A3(_2002_),
    .B1(_2005_),
    .X(_2006_));
 sky130_fd_sc_hd__a22o_1 _6532_ (.A1(_0650_),
    .A2(_0767_),
    .B1(_0769_),
    .B2(_0688_),
    .X(_2007_));
 sky130_fd_sc_hd__a22oi_1 _6533_ (.A1(_0688_),
    .A2(_1986_),
    .B1(_2007_),
    .B2(_1988_),
    .Y(_2008_));
 sky130_fd_sc_hd__nand2_1 _6534_ (.A(_2006_),
    .B(_2008_),
    .Y(net691));
 sky130_fd_sc_hd__inv_2 _6535_ (.A(_0743_),
    .Y(_2009_));
 sky130_fd_sc_hd__or2_1 _6536_ (.A(_0198_),
    .B(_0690_),
    .X(_2010_));
 sky130_fd_sc_hd__o21ai_1 _6537_ (.A1(_0855_),
    .A2(_2009_),
    .B1(_2010_),
    .Y(_2011_));
 sky130_fd_sc_hd__inv_2 _6538_ (.A(_2011_),
    .Y(_2012_));
 sky130_fd_sc_hd__a22o_1 _6539_ (.A1(_0698_),
    .A2(_0522_),
    .B1(_0693_),
    .B2(_0694_),
    .X(_2013_));
 sky130_fd_sc_hd__mux2_1 _6540_ (.A0(_2013_),
    .A1(_0679_),
    .S(_0862_),
    .X(_2014_));
 sky130_fd_sc_hd__a22o_1 _6541_ (.A1(_0698_),
    .A2(_1955_),
    .B1(_2014_),
    .B2(_1997_),
    .X(_2015_));
 sky130_fd_sc_hd__nand2_1 _6542_ (.A(_2015_),
    .B(_1999_),
    .Y(_2016_));
 sky130_fd_sc_hd__nand2_1 _6543_ (.A(_1976_),
    .B(_0785_),
    .Y(_2017_));
 sky130_fd_sc_hd__nand2_1 _6544_ (.A(_0683_),
    .B(_0785_),
    .Y(_2018_));
 sky130_fd_sc_hd__mux2_1 _6545_ (.A0(_2017_),
    .A1(_2018_),
    .S(_0558_),
    .X(_2019_));
 sky130_fd_sc_hd__a22o_1 _6546_ (.A1(_0710_),
    .A2(_0510_),
    .B1(_0612_),
    .B2(_0715_),
    .X(_2020_));
 sky130_fd_sc_hd__nor2_1 _6547_ (.A(_0719_),
    .B(_2020_),
    .Y(_2021_));
 sky130_fd_sc_hd__a211o_1 _6548_ (.A1(_0719_),
    .A2(_2019_),
    .B1(_1889_),
    .C1(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__buf_6 _6549_ (.A(_1887_),
    .X(_2023_));
 sky130_fd_sc_hd__nand2_1 _6550_ (.A(_0710_),
    .B(_2023_),
    .Y(_2024_));
 sky130_fd_sc_hd__inv_2 _6551_ (.A(_0739_),
    .Y(_2025_));
 sky130_fd_sc_hd__a22o_1 _6552_ (.A1(_0739_),
    .A2(_0730_),
    .B1(_0729_),
    .B2(_0727_),
    .X(_2026_));
 sky130_fd_sc_hd__inv_2 _6553_ (.A(_2026_),
    .Y(_2027_));
 sky130_fd_sc_hd__a221o_1 _6554_ (.A1(_2025_),
    .A2(_1900_),
    .B1(_2027_),
    .B2(_2003_),
    .C1(_1910_),
    .X(_2028_));
 sky130_fd_sc_hd__a41o_1 _6555_ (.A1(_2016_),
    .A2(_1947_),
    .A3(_2022_),
    .A4(_2024_),
    .B1(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__o221ai_4 _6556_ (.A1(_0742_),
    .A2(_1907_),
    .B1(_2012_),
    .B2(_1908_),
    .C1(_2029_),
    .Y(net692));
 sky130_fd_sc_hd__nand2_1 _6557_ (.A(_0705_),
    .B(_1997_),
    .Y(_2030_));
 sky130_fd_sc_hd__nor2_1 _6558_ (.A(_1973_),
    .B(_0700_),
    .Y(_2031_));
 sky130_fd_sc_hd__o21ai_1 _6559_ (.A1(_1914_),
    .A2(_2031_),
    .B1(_1917_),
    .Y(_2032_));
 sky130_fd_sc_hd__nor2_1 _6560_ (.A(_1889_),
    .B(_0720_),
    .Y(_2033_));
 sky130_fd_sc_hd__a221o_1 _6561_ (.A1(_0748_),
    .A2(_2023_),
    .B1(_2030_),
    .B2(_2032_),
    .C1(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__nand2_1 _6562_ (.A(_2034_),
    .B(_1929_),
    .Y(_2035_));
 sky130_fd_sc_hd__nand2_1 _6563_ (.A(_0732_),
    .B(_0761_),
    .Y(_2036_));
 sky130_fd_sc_hd__o21ai_1 _6564_ (.A1(_0761_),
    .A2(_0758_),
    .B1(_2036_),
    .Y(_2037_));
 sky130_fd_sc_hd__nand2_1 _6565_ (.A(_2037_),
    .B(_2004_),
    .Y(_2038_));
 sky130_fd_sc_hd__or2_1 _6566_ (.A(_1983_),
    .B(_0752_),
    .X(_2039_));
 sky130_fd_sc_hd__nand2_1 _6567_ (.A(_0746_),
    .B(_0888_),
    .Y(_2040_));
 sky130_fd_sc_hd__mux2_1 _6568_ (.A0(_2009_),
    .A1(_2040_),
    .S(_0769_),
    .X(_2041_));
 sky130_fd_sc_hd__nor2_1 _6569_ (.A(_0887_),
    .B(_2007_),
    .Y(_2042_));
 sky130_fd_sc_hd__a21oi_1 _6570_ (.A1(_2041_),
    .A2(_0887_),
    .B1(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__a22o_1 _6571_ (.A1(_0746_),
    .A2(_1906_),
    .B1(_2043_),
    .B2(_1988_),
    .X(_2044_));
 sky130_fd_sc_hd__a41o_1 _6572_ (.A1(_2035_),
    .A2(_1932_),
    .A3(_2038_),
    .A4(_2039_),
    .B1(_2044_),
    .X(net693));
 sky130_fd_sc_hd__or2_1 _6573_ (.A(_0781_),
    .B(_2020_),
    .X(_2045_));
 sky130_fd_sc_hd__o21ai_1 _6574_ (.A1(_0719_),
    .A2(_0782_),
    .B1(_2045_),
    .Y(_2046_));
 sky130_fd_sc_hd__or4b_1 _6575_ (.A(_1007_),
    .B(_0800_),
    .C(_4118_),
    .D_N(_0812_),
    .X(_2047_));
 sky130_fd_sc_hd__nor2_1 _6576_ (.A(_1973_),
    .B(_0797_),
    .Y(_2048_));
 sky130_fd_sc_hd__o21ai_1 _6577_ (.A1(_1914_),
    .A2(_2048_),
    .B1(_1917_),
    .Y(_2049_));
 sky130_fd_sc_hd__nor2_1 _6578_ (.A(_1920_),
    .B(_0780_),
    .Y(_2050_));
 sky130_fd_sc_hd__a221o_1 _6579_ (.A1(_2046_),
    .A2(_1924_),
    .B1(_2047_),
    .B2(_2049_),
    .C1(_2050_),
    .X(_2051_));
 sky130_fd_sc_hd__nand2_1 _6580_ (.A(_2051_),
    .B(_1929_),
    .Y(_2052_));
 sky130_fd_sc_hd__nand2_1 _6581_ (.A(_2027_),
    .B(_0761_),
    .Y(_2053_));
 sky130_fd_sc_hd__o21ai_1 _6582_ (.A1(_0761_),
    .A2(_0775_),
    .B1(_2053_),
    .Y(_2054_));
 sky130_fd_sc_hd__nand2_1 _6583_ (.A(_2054_),
    .B(_2004_),
    .Y(_2055_));
 sky130_fd_sc_hd__nand2_1 _6584_ (.A(_0777_),
    .B(_1900_),
    .Y(_2056_));
 sky130_fd_sc_hd__nand2_1 _6585_ (.A(_2012_),
    .B(_1280_),
    .Y(_2057_));
 sky130_fd_sc_hd__o21ai_1 _6586_ (.A1(_1280_),
    .A2(_0770_),
    .B1(_2057_),
    .Y(_2058_));
 sky130_fd_sc_hd__inv_2 _6587_ (.A(_2058_),
    .Y(_2059_));
 sky130_fd_sc_hd__a22o_1 _6588_ (.A1(_0765_),
    .A2(_1906_),
    .B1(_2059_),
    .B2(_1988_),
    .X(_2060_));
 sky130_fd_sc_hd__a41o_1 _6589_ (.A1(_2052_),
    .A2(_1932_),
    .A3(_2055_),
    .A4(_2056_),
    .B1(_2060_),
    .X(net694));
 sky130_fd_sc_hd__or2_1 _6590_ (.A(_0704_),
    .B(_0702_),
    .X(_2061_));
 sky130_fd_sc_hd__or2_1 _6591_ (.A(_0862_),
    .B(_0821_),
    .X(_2062_));
 sky130_fd_sc_hd__a32o_1 _6592_ (.A1(_2061_),
    .A2(_2062_),
    .A3(_1953_),
    .B1(_0808_),
    .B2(_1955_),
    .X(_2063_));
 sky130_fd_sc_hd__or2_1 _6593_ (.A(_0781_),
    .B(_0713_),
    .X(_2064_));
 sky130_fd_sc_hd__o21ai_1 _6594_ (.A1(_0719_),
    .A2(_0834_),
    .B1(_2064_),
    .Y(_2065_));
 sky130_fd_sc_hd__a2bb2o_1 _6595_ (.A1_N(_1889_),
    .A2_N(_2065_),
    .B1(_0788_),
    .B2(_2023_),
    .X(_2066_));
 sky130_fd_sc_hd__a211o_1 _6596_ (.A1(_2063_),
    .A2(_1999_),
    .B1(_1926_),
    .C1(_2066_),
    .X(_2067_));
 sky130_fd_sc_hd__or2_1 _6597_ (.A(_1981_),
    .B(_0762_),
    .X(_2068_));
 sky130_fd_sc_hd__nand2_1 _6598_ (.A(_0851_),
    .B(_1900_),
    .Y(_2069_));
 sky130_fd_sc_hd__a22o_1 _6599_ (.A1(_0854_),
    .A2(_1906_),
    .B1(_0858_),
    .B2(_1988_),
    .X(_2070_));
 sky130_fd_sc_hd__a41o_1 _6600_ (.A1(_2067_),
    .A2(_1932_),
    .A3(_2068_),
    .A4(_2069_),
    .B1(_2070_),
    .X(net695));
 sky130_fd_sc_hd__a22o_1 _6601_ (.A1(_0826_),
    .A2(_1955_),
    .B1(_0814_),
    .B2(_1997_),
    .X(_2071_));
 sky130_fd_sc_hd__a22o_1 _6602_ (.A1(_0784_),
    .A2(_2023_),
    .B1(_0793_),
    .B2(_1924_),
    .X(_2072_));
 sky130_fd_sc_hd__a211o_1 _6603_ (.A1(_2071_),
    .A2(_1999_),
    .B1(_1926_),
    .C1(_2072_),
    .X(_2073_));
 sky130_fd_sc_hd__o221a_1 _6604_ (.A1(_0773_),
    .A2(_1983_),
    .B1(_1981_),
    .B2(_0776_),
    .C1(_1931_),
    .X(_2074_));
 sky130_fd_sc_hd__a22o_1 _6605_ (.A1(_0885_),
    .A2(_1911_),
    .B1(_2073_),
    .B2(_2074_),
    .X(net697));
 sky130_fd_sc_hd__a22o_1 _6606_ (.A1(_0863_),
    .A2(_1955_),
    .B1(_0831_),
    .B2(_1997_),
    .X(_2075_));
 sky130_fd_sc_hd__a22o_1 _6607_ (.A1(_0628_),
    .A2(_2023_),
    .B1(_0838_),
    .B2(_1924_),
    .X(_2076_));
 sky130_fd_sc_hd__a211o_1 _6608_ (.A1(_2075_),
    .A2(_1999_),
    .B1(_1926_),
    .C1(_2076_),
    .X(_2077_));
 sky130_fd_sc_hd__nand2_1 _6609_ (.A(_0849_),
    .B(_2004_),
    .Y(_2078_));
 sky130_fd_sc_hd__o21a_1 _6610_ (.A1(_1983_),
    .A2(_0843_),
    .B1(_1931_),
    .X(_2079_));
 sky130_fd_sc_hd__nand2_1 _6611_ (.A(_0896_),
    .B(_0769_),
    .Y(_2080_));
 sky130_fd_sc_hd__o21ai_1 _6612_ (.A1(_0769_),
    .A2(_0889_),
    .B1(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__or2_1 _6613_ (.A(_1280_),
    .B(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__a22o_1 _6614_ (.A1(_0896_),
    .A2(_1986_),
    .B1(_2082_),
    .B2(_1988_),
    .X(_2083_));
 sky130_fd_sc_hd__a31o_1 _6615_ (.A1(_2077_),
    .A2(_2078_),
    .A3(_2079_),
    .B1(_2083_),
    .X(net698));
 sky130_fd_sc_hd__nand2_1 _6616_ (.A(_0872_),
    .B(_1997_),
    .Y(_2084_));
 sky130_fd_sc_hd__nor2_1 _6617_ (.A(_1973_),
    .B(_0867_),
    .Y(_2085_));
 sky130_fd_sc_hd__o21ai_1 _6618_ (.A1(_1914_),
    .A2(_2085_),
    .B1(_1917_),
    .Y(_2086_));
 sky130_fd_sc_hd__a22o_1 _6619_ (.A1(_0925_),
    .A2(_1891_),
    .B1(_2084_),
    .B2(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__nand2_1 _6620_ (.A(_2087_),
    .B(_1929_),
    .Y(_2088_));
 sky130_fd_sc_hd__nand2_1 _6621_ (.A(_0881_),
    .B(_2004_),
    .Y(_2089_));
 sky130_fd_sc_hd__inv_2 _6622_ (.A(_0877_),
    .Y(_2090_));
 sky130_fd_sc_hd__nand2_1 _6623_ (.A(_2090_),
    .B(_1900_),
    .Y(_2091_));
 sky130_fd_sc_hd__a22o_1 _6624_ (.A1(_0893_),
    .A2(_1906_),
    .B1(_0901_),
    .B2(_1988_),
    .X(_2092_));
 sky130_fd_sc_hd__a41o_1 _6625_ (.A1(_2088_),
    .A2(_1932_),
    .A3(_2089_),
    .A4(_2091_),
    .B1(_2092_),
    .X(net699));
 sky130_fd_sc_hd__nand2_1 _6626_ (.A(_0940_),
    .B(_0888_),
    .Y(_2093_));
 sky130_fd_sc_hd__mux2_1 _6627_ (.A0(_0894_),
    .A1(_2093_),
    .S(_0769_),
    .X(_2094_));
 sky130_fd_sc_hd__nand2_1 _6628_ (.A(_2094_),
    .B(_0887_),
    .Y(_2095_));
 sky130_fd_sc_hd__o21ai_1 _6629_ (.A1(_0887_),
    .A2(_2081_),
    .B1(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__nand2_1 _6630_ (.A(_0940_),
    .B(_1986_),
    .Y(_2097_));
 sky130_fd_sc_hd__a22o_1 _6631_ (.A1(_0948_),
    .A2(_1955_),
    .B1(_0920_),
    .B2(_1997_),
    .X(_2098_));
 sky130_fd_sc_hd__nand2_1 _6632_ (.A(_2098_),
    .B(_1999_),
    .Y(_2099_));
 sky130_fd_sc_hd__nand2_1 _6633_ (.A(_0909_),
    .B(_1924_),
    .Y(_2100_));
 sky130_fd_sc_hd__nand2_1 _6634_ (.A(_0904_),
    .B(_2023_),
    .Y(_2101_));
 sky130_fd_sc_hd__inv_2 _6635_ (.A(_0955_),
    .Y(_2102_));
 sky130_fd_sc_hd__a22o_1 _6636_ (.A1(_0877_),
    .A2(_0729_),
    .B1(_0730_),
    .B2(_0955_),
    .X(_2103_));
 sky130_fd_sc_hd__inv_2 _6637_ (.A(_2103_),
    .Y(_2104_));
 sky130_fd_sc_hd__a221o_1 _6638_ (.A1(_2102_),
    .A2(_1900_),
    .B1(_2104_),
    .B2(_2003_),
    .C1(_1910_),
    .X(_2105_));
 sky130_fd_sc_hd__a41o_1 _6639_ (.A1(_2099_),
    .A2(_1947_),
    .A3(_2100_),
    .A4(_2101_),
    .B1(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__o211ai_2 _6640_ (.A1(_2096_),
    .A2(_1908_),
    .B1(_2097_),
    .C1(_2106_),
    .Y(net700));
 sky130_fd_sc_hd__a22o_1 _6641_ (.A1(_0980_),
    .A2(_0730_),
    .B1(_0729_),
    .B2(_0955_),
    .X(_2107_));
 sky130_fd_sc_hd__inv_2 _6642_ (.A(_2107_),
    .Y(_2108_));
 sky130_fd_sc_hd__mux2_1 _6643_ (.A0(_0879_),
    .A1(_2108_),
    .S(_0841_),
    .X(_2109_));
 sky130_fd_sc_hd__inv_2 _6644_ (.A(_0971_),
    .Y(_2110_));
 sky130_fd_sc_hd__nand2_1 _6645_ (.A(_0932_),
    .B(_1953_),
    .Y(_2111_));
 sky130_fd_sc_hd__nor2_1 _6646_ (.A(_1973_),
    .B(_0929_),
    .Y(_2112_));
 sky130_fd_sc_hd__o21ai_1 _6647_ (.A1(_1914_),
    .A2(_2112_),
    .B1(_1917_),
    .Y(_2113_));
 sky130_fd_sc_hd__nor2_1 _6648_ (.A(_1920_),
    .B(_0944_),
    .Y(_2114_));
 sky130_fd_sc_hd__a221o_1 _6649_ (.A1(_2110_),
    .A2(_1923_),
    .B1(_2111_),
    .B2(_2113_),
    .C1(_2114_),
    .X(_2115_));
 sky130_fd_sc_hd__o21ai_1 _6650_ (.A1(_1983_),
    .A2(_0980_),
    .B1(_1930_),
    .Y(_2116_));
 sky130_fd_sc_hd__a221o_1 _6651_ (.A1(_2109_),
    .A2(_2004_),
    .B1(_2115_),
    .B2(_1947_),
    .C1(_2116_),
    .X(_2117_));
 sky130_fd_sc_hd__a21bo_1 _6652_ (.A1(_0983_),
    .A2(_1911_),
    .B1_N(_2117_),
    .X(net701));
 sky130_fd_sc_hd__inv_2 _6653_ (.A(_0966_),
    .Y(_2118_));
 sky130_fd_sc_hd__a21o_1 _6654_ (.A1(_1008_),
    .A2(_0704_),
    .B1(_0950_),
    .X(_2119_));
 sky130_fd_sc_hd__a22o_1 _6655_ (.A1(_2118_),
    .A2(_1955_),
    .B1(_2119_),
    .B2(_1997_),
    .X(_2120_));
 sky130_fd_sc_hd__a22o_1 _6656_ (.A1(_0942_),
    .A2(_2023_),
    .B1(_0947_),
    .B2(_1924_),
    .X(_2121_));
 sky130_fd_sc_hd__a211o_1 _6657_ (.A1(_2120_),
    .A2(_1999_),
    .B1(_1926_),
    .C1(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__nand2_1 _6658_ (.A(_1014_),
    .B(_0844_),
    .Y(_2123_));
 sky130_fd_sc_hd__nand2_1 _6659_ (.A(_0980_),
    .B(_0844_),
    .Y(_2124_));
 sky130_fd_sc_hd__mux2_1 _6660_ (.A0(_2123_),
    .A1(_2124_),
    .S(_0090_),
    .X(_2125_));
 sky130_fd_sc_hd__mux2_1 _6661_ (.A0(_2104_),
    .A1(_2125_),
    .S(_0841_),
    .X(_2126_));
 sky130_fd_sc_hd__nand2_1 _6662_ (.A(_2126_),
    .B(_2004_),
    .Y(_2127_));
 sky130_fd_sc_hd__o211a_1 _6663_ (.A1(_1014_),
    .A2(_1983_),
    .B1(_1931_),
    .C1(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__a22o_2 _6664_ (.A1(_0986_),
    .A2(_1911_),
    .B1(_2122_),
    .B2(_2128_),
    .X(net702));
 sky130_fd_sc_hd__a22o_1 _6665_ (.A1(_1014_),
    .A2(_0111_),
    .B1(_0730_),
    .B2(_1019_),
    .X(_2129_));
 sky130_fd_sc_hd__inv_2 _6666_ (.A(_2129_),
    .Y(_2130_));
 sky130_fd_sc_hd__mux2_1 _6667_ (.A0(_2108_),
    .A1(_2130_),
    .S(_0841_),
    .X(_2131_));
 sky130_fd_sc_hd__nand2_1 _6668_ (.A(_0969_),
    .B(_1953_),
    .Y(_2132_));
 sky130_fd_sc_hd__nor2_1 _6669_ (.A(_1973_),
    .B(_0961_),
    .Y(_2133_));
 sky130_fd_sc_hd__o21ai_1 _6670_ (.A1(_1914_),
    .A2(_2133_),
    .B1(_1917_),
    .Y(_2134_));
 sky130_fd_sc_hd__nor2_1 _6671_ (.A(_1920_),
    .B(_0973_),
    .Y(_2135_));
 sky130_fd_sc_hd__a221o_1 _6672_ (.A1(_0976_),
    .A2(_1923_),
    .B1(_2132_),
    .B2(_2134_),
    .C1(_2135_),
    .X(_2136_));
 sky130_fd_sc_hd__o21ai_1 _6673_ (.A1(_1901_),
    .A2(_1019_),
    .B1(_1930_),
    .Y(_2137_));
 sky130_fd_sc_hd__a221o_1 _6674_ (.A1(_2131_),
    .A2(_2004_),
    .B1(_2136_),
    .B2(_1947_),
    .C1(_2137_),
    .X(_2138_));
 sky130_fd_sc_hd__a21bo_1 _6675_ (.A1(_1017_),
    .A2(_1911_),
    .B1_N(_2138_),
    .X(net703));
 sky130_fd_sc_hd__or4b_1 _6676_ (.A(_1007_),
    .B(_0800_),
    .C(_4118_),
    .D_N(_1059_),
    .X(_2139_));
 sky130_fd_sc_hd__nor2_1 _6677_ (.A(_1973_),
    .B(_1034_),
    .Y(_2140_));
 sky130_fd_sc_hd__o21ai_1 _6678_ (.A1(_1914_),
    .A2(_2140_),
    .B1(_1917_),
    .Y(_2141_));
 sky130_fd_sc_hd__nor2_1 _6679_ (.A(_1920_),
    .B(_0990_),
    .Y(_2142_));
 sky130_fd_sc_hd__a221o_1 _6680_ (.A1(_0993_),
    .A2(_1923_),
    .B1(_2139_),
    .B2(_2141_),
    .C1(_2142_),
    .X(_2143_));
 sky130_fd_sc_hd__nand2_1 _6681_ (.A(_2143_),
    .B(_1929_),
    .Y(_2144_));
 sky130_fd_sc_hd__a22o_1 _6682_ (.A1(_1019_),
    .A2(_0572_),
    .B1(_0771_),
    .B2(_1064_),
    .X(_2145_));
 sky130_fd_sc_hd__or2_1 _6683_ (.A(_1981_),
    .B(_2145_),
    .X(_2146_));
 sky130_fd_sc_hd__o21a_1 _6684_ (.A1(_1983_),
    .A2(_1064_),
    .B1(_1931_),
    .X(_2147_));
 sky130_fd_sc_hd__a32o_2 _6685_ (.A1(_2144_),
    .A2(_2146_),
    .A3(_2147_),
    .B1(_1050_),
    .B2(_1911_),
    .X(net704));
 sky130_fd_sc_hd__a2bb2o_1 _6686_ (.A1_N(_1895_),
    .A2_N(_1038_),
    .B1(_1068_),
    .B2(_1955_),
    .X(_2148_));
 sky130_fd_sc_hd__a22o_1 _6687_ (.A1(_1021_),
    .A2(_2023_),
    .B1(_1023_),
    .B2(_1924_),
    .X(_2149_));
 sky130_fd_sc_hd__a211o_1 _6688_ (.A1(_2148_),
    .A2(_1999_),
    .B1(_1926_),
    .C1(_2149_),
    .X(_2150_));
 sky130_fd_sc_hd__mux2_1 _6689_ (.A0(_1079_),
    .A1(_2130_),
    .S(_0761_),
    .X(_2151_));
 sky130_fd_sc_hd__inv_2 _6690_ (.A(_2151_),
    .Y(_2152_));
 sky130_fd_sc_hd__o221a_1 _6691_ (.A1(_1077_),
    .A2(_1983_),
    .B1(_1981_),
    .B2(_2152_),
    .C1(_1931_),
    .X(_2153_));
 sky130_fd_sc_hd__a22o_2 _6692_ (.A1(_1067_),
    .A2(_1911_),
    .B1(_2150_),
    .B2(_2153_),
    .X(net705));
 sky130_fd_sc_hd__mux2_1 _6693_ (.A0(_1059_),
    .A1(_1098_),
    .S(_0704_),
    .X(_2154_));
 sky130_fd_sc_hd__nand2_1 _6694_ (.A(_2154_),
    .B(_1953_),
    .Y(_2155_));
 sky130_fd_sc_hd__nor2_1 _6695_ (.A(_1973_),
    .B(_1096_),
    .Y(_2156_));
 sky130_fd_sc_hd__o21ai_1 _6696_ (.A1(_1914_),
    .A2(_2156_),
    .B1(_1917_),
    .Y(_2157_));
 sky130_fd_sc_hd__nor2_1 _6697_ (.A(_1920_),
    .B(_1052_),
    .Y(_2158_));
 sky130_fd_sc_hd__a221o_1 _6698_ (.A1(_1055_),
    .A2(_1923_),
    .B1(_2155_),
    .B2(_2157_),
    .C1(_2158_),
    .X(_2159_));
 sky130_fd_sc_hd__nand2_1 _6699_ (.A(_2159_),
    .B(_1929_),
    .Y(_2160_));
 sky130_fd_sc_hd__a22o_1 _6700_ (.A1(_1077_),
    .A2(_0572_),
    .B1(_0771_),
    .B2(_1081_),
    .X(_2161_));
 sky130_fd_sc_hd__or2_1 _6701_ (.A(_1981_),
    .B(_2161_),
    .X(_2162_));
 sky130_fd_sc_hd__o21a_1 _6702_ (.A1(_1983_),
    .A2(_1081_),
    .B1(_1931_),
    .X(_2163_));
 sky130_fd_sc_hd__a32o_2 _6703_ (.A1(_2160_),
    .A2(_2162_),
    .A3(_2163_),
    .B1(_1106_),
    .B2(_1911_),
    .X(net706));
 sky130_fd_sc_hd__o21a_1 _6704_ (.A1(_1901_),
    .A2(_1083_),
    .B1(_1930_),
    .X(_2164_));
 sky130_fd_sc_hd__mux2_1 _6705_ (.A0(_1129_),
    .A1(_1036_),
    .S(_0862_),
    .X(_2165_));
 sky130_fd_sc_hd__a22o_1 _6706_ (.A1(_1112_),
    .A2(_1892_),
    .B1(_2165_),
    .B2(_1953_),
    .X(_2166_));
 sky130_fd_sc_hd__a22o_1 _6707_ (.A1(_1071_),
    .A2(_1887_),
    .B1(_1073_),
    .B2(_1923_),
    .X(_2167_));
 sky130_fd_sc_hd__a211o_1 _6708_ (.A1(_2166_),
    .A2(_1941_),
    .B1(_1904_),
    .C1(_2167_),
    .X(_2168_));
 sky130_fd_sc_hd__o211a_1 _6709_ (.A1(_1087_),
    .A2(_1981_),
    .B1(_2164_),
    .C1(_2168_),
    .X(_2169_));
 sky130_fd_sc_hd__a221o_1 _6710_ (.A1(_1153_),
    .A2(_1986_),
    .B1(_1163_),
    .B2(_1988_),
    .C1(_2169_),
    .X(net708));
 sky130_fd_sc_hd__mux2_1 _6711_ (.A0(_1185_),
    .A1(_1098_),
    .S(_0813_),
    .X(_2170_));
 sky130_fd_sc_hd__a22o_1 _6712_ (.A1(_1174_),
    .A2(_1892_),
    .B1(_2170_),
    .B2(_1953_),
    .X(_2171_));
 sky130_fd_sc_hd__and2_1 _6713_ (.A(_2171_),
    .B(_1941_),
    .X(_2172_));
 sky130_fd_sc_hd__a221o_1 _6714_ (.A1(_1090_),
    .A2(_1887_),
    .B1(_1092_),
    .B2(_1923_),
    .C1(_1904_),
    .X(_2173_));
 sky130_fd_sc_hd__o221a_2 _6715_ (.A1(_1144_),
    .A2(_1947_),
    .B1(_2172_),
    .B2(_2173_),
    .C1(_1931_),
    .X(_2174_));
 sky130_fd_sc_hd__a221o_2 _6716_ (.A1(_1158_),
    .A2(_1986_),
    .B1(_1167_),
    .B2(_1988_),
    .C1(_2174_),
    .X(net709));
 sky130_fd_sc_hd__a2bb2o_1 _6717_ (.A1_N(_1895_),
    .A2_N(_1131_),
    .B1(_1117_),
    .B2(_1955_),
    .X(_2175_));
 sky130_fd_sc_hd__a22o_1 _6718_ (.A1(_0995_),
    .A2(_1887_),
    .B1(_1137_),
    .B2(_1923_),
    .X(_2176_));
 sky130_fd_sc_hd__a211o_1 _6719_ (.A1(_2175_),
    .A2(_1999_),
    .B1(_1926_),
    .C1(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__nand2_1 _6720_ (.A(_1149_),
    .B(_2004_),
    .Y(_2178_));
 sky130_fd_sc_hd__nand2_1 _6721_ (.A(_1142_),
    .B(_1900_),
    .Y(_2179_));
 sky130_fd_sc_hd__a22o_1 _6722_ (.A1(_1155_),
    .A2(_1906_),
    .B1(_1165_),
    .B2(_1988_),
    .X(_2180_));
 sky130_fd_sc_hd__a41o_1 _6723_ (.A1(_2177_),
    .A2(_1932_),
    .A3(_2178_),
    .A4(_2179_),
    .B1(_2180_),
    .X(net710));
 sky130_fd_sc_hd__or2_1 _6724_ (.A(_1895_),
    .B(_1187_),
    .X(_2181_));
 sky130_fd_sc_hd__nor2_1 _6725_ (.A(_1973_),
    .B(_1180_),
    .Y(_2182_));
 sky130_fd_sc_hd__o21ai_1 _6726_ (.A1(_1914_),
    .A2(_2182_),
    .B1(_1917_),
    .Y(_2183_));
 sky130_fd_sc_hd__nor2_1 _6727_ (.A(_1920_),
    .B(_0997_),
    .Y(_2184_));
 sky130_fd_sc_hd__a221o_2 _6728_ (.A1(_1191_),
    .A2(_1924_),
    .B1(_2181_),
    .B2(_2183_),
    .C1(_2184_),
    .X(_2185_));
 sky130_fd_sc_hd__nand2_1 _6729_ (.A(_2185_),
    .B(_1929_),
    .Y(_2186_));
 sky130_fd_sc_hd__a22o_1 _6730_ (.A1(_1141_),
    .A2(_0572_),
    .B1(_0771_),
    .B2(_1213_),
    .X(_2187_));
 sky130_fd_sc_hd__or2_1 _6731_ (.A(_1981_),
    .B(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__inv_2 _6732_ (.A(_1213_),
    .Y(_2189_));
 sky130_fd_sc_hd__nand2_1 _6733_ (.A(_2189_),
    .B(_1900_),
    .Y(_2190_));
 sky130_fd_sc_hd__a22o_1 _6734_ (.A1(_1169_),
    .A2(_1906_),
    .B1(_1173_),
    .B2(_1988_),
    .X(_2191_));
 sky130_fd_sc_hd__a41o_2 _6735_ (.A1(_2186_),
    .A2(_1932_),
    .A3(_2188_),
    .A4(_2190_),
    .B1(_2191_),
    .X(net711));
 sky130_fd_sc_hd__o21a_1 _6736_ (.A1(_1901_),
    .A2(_1215_),
    .B1(_1930_),
    .X(_2192_));
 sky130_fd_sc_hd__inv_2 _6737_ (.A(_1203_),
    .Y(_2193_));
 sky130_fd_sc_hd__a22o_1 _6738_ (.A1(_2193_),
    .A2(_1892_),
    .B1(_1208_),
    .B2(_1953_),
    .X(_2194_));
 sky130_fd_sc_hd__a22o_1 _6739_ (.A1(_1000_),
    .A2(_1887_),
    .B1(_1199_),
    .B2(_1923_),
    .X(_2195_));
 sky130_fd_sc_hd__a211o_1 _6740_ (.A1(_2194_),
    .A2(_1941_),
    .B1(_1904_),
    .C1(_2195_),
    .X(_2196_));
 sky130_fd_sc_hd__o211a_1 _6741_ (.A1(_1219_),
    .A2(_1981_),
    .B1(_2192_),
    .C1(_2196_),
    .X(_2197_));
 sky130_fd_sc_hd__a221o_2 _6742_ (.A1(_1232_),
    .A2(_1986_),
    .B1(_1233_),
    .B2(_1988_),
    .C1(_2197_),
    .X(net712));
 sky130_fd_sc_hd__nand2_1 _6743_ (.A(_1169_),
    .B(_0769_),
    .Y(_2198_));
 sky130_fd_sc_hd__nor2_1 _6744_ (.A(_1279_),
    .B(_1287_),
    .Y(_2199_));
 sky130_fd_sc_hd__a31o_1 _6745_ (.A1(_1280_),
    .A2(_1171_),
    .A3(_2198_),
    .B1(_2199_),
    .X(_2200_));
 sky130_fd_sc_hd__inv_2 _6746_ (.A(_2200_),
    .Y(_2201_));
 sky130_fd_sc_hd__a22o_1 _6747_ (.A1(_1215_),
    .A2(_0572_),
    .B1(_0771_),
    .B2(_1277_),
    .X(_2202_));
 sky130_fd_sc_hd__o21a_1 _6748_ (.A1(_1901_),
    .A2(_1277_),
    .B1(_1930_),
    .X(_2203_));
 sky130_fd_sc_hd__nand2_1 _6749_ (.A(_1002_),
    .B(_2023_),
    .Y(_2204_));
 sky130_fd_sc_hd__a22o_1 _6750_ (.A1(_1257_),
    .A2(_1892_),
    .B1(_1227_),
    .B2(_1953_),
    .X(_2205_));
 sky130_fd_sc_hd__nand2_1 _6751_ (.A(_2205_),
    .B(_1941_),
    .Y(_2206_));
 sky130_fd_sc_hd__o2111ai_4 _6752_ (.A1(_1005_),
    .A2(_1889_),
    .B1(_1947_),
    .C1(_2204_),
    .D1(_2206_),
    .Y(_2207_));
 sky130_fd_sc_hd__o211a_1 _6753_ (.A1(_2202_),
    .A2(_1981_),
    .B1(_2203_),
    .C1(_2207_),
    .X(_2208_));
 sky130_fd_sc_hd__a221o_1 _6754_ (.A1(_1256_),
    .A2(_1986_),
    .B1(_2201_),
    .B2(_1988_),
    .C1(_2208_),
    .X(net713));
 sky130_fd_sc_hd__nand2_1 _6755_ (.A(_1242_),
    .B(_1997_),
    .Y(_2209_));
 sky130_fd_sc_hd__nor2_1 _6756_ (.A(_1973_),
    .B(_1238_),
    .Y(_2210_));
 sky130_fd_sc_hd__o21ai_1 _6757_ (.A1(_1914_),
    .A2(_2210_),
    .B1(_1917_),
    .Y(_2211_));
 sky130_fd_sc_hd__nor2_1 _6758_ (.A(_1920_),
    .B(_1246_),
    .Y(_2212_));
 sky130_fd_sc_hd__a221o_2 _6759_ (.A1(_1249_),
    .A2(_1924_),
    .B1(_2209_),
    .B2(_2211_),
    .C1(_2212_),
    .X(_2213_));
 sky130_fd_sc_hd__nand2_1 _6760_ (.A(_2213_),
    .B(_1929_),
    .Y(_2214_));
 sky130_fd_sc_hd__nand2_1 _6761_ (.A(_1306_),
    .B(_2004_),
    .Y(_2215_));
 sky130_fd_sc_hd__nand2_1 _6762_ (.A(_1310_),
    .B(_1900_),
    .Y(_2216_));
 sky130_fd_sc_hd__a22o_1 _6763_ (.A1(_1256_),
    .A2(_0766_),
    .B1(_0198_),
    .B2(_1282_),
    .X(_2217_));
 sky130_fd_sc_hd__inv_2 _6764_ (.A(_2217_),
    .Y(_2218_));
 sky130_fd_sc_hd__nand2_1 _6765_ (.A(_2218_),
    .B(_0886_),
    .Y(_2219_));
 sky130_fd_sc_hd__o21ai_1 _6766_ (.A1(_0886_),
    .A2(_1233_),
    .B1(_2219_),
    .Y(_2220_));
 sky130_fd_sc_hd__inv_2 _6767_ (.A(_2220_),
    .Y(_2221_));
 sky130_fd_sc_hd__a22o_1 _6768_ (.A1(_1282_),
    .A2(_1906_),
    .B1(_2221_),
    .B2(_1988_),
    .X(_2222_));
 sky130_fd_sc_hd__a41o_2 _6769_ (.A1(_2214_),
    .A2(_1932_),
    .A3(_2215_),
    .A4(_2216_),
    .B1(_2222_),
    .X(net714));
 sky130_fd_sc_hd__inv_2 _6770_ (.A(_1299_),
    .Y(_2223_));
 sky130_fd_sc_hd__nand2_1 _6771_ (.A(_1304_),
    .B(_0572_),
    .Y(_2224_));
 sky130_fd_sc_hd__o21ai_1 _6772_ (.A1(_0090_),
    .A2(_2223_),
    .B1(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__o21a_1 _6773_ (.A1(_1901_),
    .A2(_1299_),
    .B1(_1930_),
    .X(_2226_));
 sky130_fd_sc_hd__a22o_1 _6774_ (.A1(_1260_),
    .A2(_1892_),
    .B1(_1266_),
    .B2(_1953_),
    .X(_2227_));
 sky130_fd_sc_hd__a2bb2o_1 _6775_ (.A1_N(_1889_),
    .A2_N(_1273_),
    .B1(_1269_),
    .B2(_1887_),
    .X(_2228_));
 sky130_fd_sc_hd__a211o_1 _6776_ (.A1(_2227_),
    .A2(_1941_),
    .B1(_1904_),
    .C1(_2228_),
    .X(_2229_));
 sky130_fd_sc_hd__o211a_1 _6777_ (.A1(_2225_),
    .A2(_1981_),
    .B1(_2226_),
    .C1(_2229_),
    .X(_2230_));
 sky130_fd_sc_hd__a221o_1 _6778_ (.A1(_1284_),
    .A2(_1986_),
    .B1(_1289_),
    .B2(_1988_),
    .C1(_2230_),
    .X(net715));
 sky130_fd_sc_hd__o21ai_2 _6779_ (.A1(_0719_),
    .A2(_1350_),
    .B1(_1292_),
    .Y(_2231_));
 sky130_fd_sc_hd__nor2_1 _6780_ (.A(_0704_),
    .B(_1241_),
    .Y(_2232_));
 sky130_fd_sc_hd__a211o_1 _6781_ (.A1(_1340_),
    .A2(_0704_),
    .B1(_2232_),
    .C1(_1895_),
    .X(_2233_));
 sky130_fd_sc_hd__nor2_1 _6782_ (.A(_1973_),
    .B(_1322_),
    .Y(_2234_));
 sky130_fd_sc_hd__o21ai_1 _6783_ (.A1(_1914_),
    .A2(_2234_),
    .B1(_1917_),
    .Y(_2235_));
 sky130_fd_sc_hd__nand2_1 _6784_ (.A(_2233_),
    .B(_2235_),
    .Y(_2236_));
 sky130_fd_sc_hd__o221a_1 _6785_ (.A1(_1335_),
    .A2(_1920_),
    .B1(_2231_),
    .B2(_1889_),
    .C1(_2236_),
    .X(_2237_));
 sky130_fd_sc_hd__or2_2 _6786_ (.A(_1926_),
    .B(_2237_),
    .X(_2238_));
 sky130_fd_sc_hd__nand2_1 _6787_ (.A(_1308_),
    .B(_2004_),
    .Y(_2239_));
 sky130_fd_sc_hd__or2_1 _6788_ (.A(_1983_),
    .B(_1301_),
    .X(_2240_));
 sky130_fd_sc_hd__mux2_1 _6789_ (.A0(_1358_),
    .A1(_2218_),
    .S(_1280_),
    .X(_2241_));
 sky130_fd_sc_hd__a2bb2o_1 _6790_ (.A1_N(_1908_),
    .A2_N(_2241_),
    .B1(_1333_),
    .B2(_1986_),
    .X(_2242_));
 sky130_fd_sc_hd__a41o_1 _6791_ (.A1(_2238_),
    .A2(_1932_),
    .A3(_2239_),
    .A4(_2240_),
    .B1(_2242_),
    .X(net716));
 sky130_fd_sc_hd__a22o_1 _6792_ (.A1(_1373_),
    .A2(_1955_),
    .B1(_1325_),
    .B2(_1997_),
    .X(_2243_));
 sky130_fd_sc_hd__mux2_1 _6793_ (.A0(_1271_),
    .A1(_1363_),
    .S(_0717_),
    .X(_2244_));
 sky130_fd_sc_hd__a2bb2o_1 _6794_ (.A1_N(_1889_),
    .A2_N(_2244_),
    .B1(_1347_),
    .B2(_2023_),
    .X(_2245_));
 sky130_fd_sc_hd__a211o_1 _6795_ (.A1(_2243_),
    .A2(_1999_),
    .B1(_1926_),
    .C1(_2245_),
    .X(_2246_));
 sky130_fd_sc_hd__a22o_1 _6796_ (.A1(_1301_),
    .A2(_0729_),
    .B1(_0730_),
    .B2(_1390_),
    .X(_2247_));
 sky130_fd_sc_hd__inv_2 _6797_ (.A(_2247_),
    .Y(_2248_));
 sky130_fd_sc_hd__nand2_1 _6798_ (.A(_2248_),
    .B(_0841_),
    .Y(_2249_));
 sky130_fd_sc_hd__o21ai_1 _6799_ (.A1(_0841_),
    .A2(_2225_),
    .B1(_2249_),
    .Y(_2250_));
 sky130_fd_sc_hd__nand2_1 _6800_ (.A(_2250_),
    .B(_2004_),
    .Y(_2251_));
 sky130_fd_sc_hd__or2_1 _6801_ (.A(_1983_),
    .B(_1390_),
    .X(_2252_));
 sky130_fd_sc_hd__nand2_1 _6802_ (.A(_1286_),
    .B(_1280_),
    .Y(_2253_));
 sky130_fd_sc_hd__o21ai_1 _6803_ (.A1(_1280_),
    .A2(_1398_),
    .B1(_2253_),
    .Y(_2254_));
 sky130_fd_sc_hd__inv_2 _6804_ (.A(_2254_),
    .Y(_2255_));
 sky130_fd_sc_hd__a22o_1 _6805_ (.A1(_1361_),
    .A2(_1906_),
    .B1(_2255_),
    .B2(_1987_),
    .X(_2256_));
 sky130_fd_sc_hd__a41o_2 _6806_ (.A1(_2246_),
    .A2(_1932_),
    .A3(_2251_),
    .A4(_2252_),
    .B1(_2256_),
    .X(net717));
 sky130_fd_sc_hd__nor2_1 _6807_ (.A(_0862_),
    .B(_1413_),
    .Y(_2257_));
 sky130_fd_sc_hd__o21ai_1 _6808_ (.A1(_2257_),
    .A2(_1341_),
    .B1(_1997_),
    .Y(_2258_));
 sky130_fd_sc_hd__nor2_1 _6809_ (.A(_1973_),
    .B(_1382_),
    .Y(_2259_));
 sky130_fd_sc_hd__o21ai_1 _6810_ (.A1(_1914_),
    .A2(_2259_),
    .B1(_1917_),
    .Y(_2260_));
 sky130_fd_sc_hd__nor2_1 _6811_ (.A(_1920_),
    .B(_1345_),
    .Y(_2261_));
 sky130_fd_sc_hd__a221o_2 _6812_ (.A1(_1352_),
    .A2(_1924_),
    .B1(_2258_),
    .B2(_2260_),
    .C1(_2261_),
    .X(_2262_));
 sky130_fd_sc_hd__nand2_1 _6813_ (.A(_2262_),
    .B(_1929_),
    .Y(_2263_));
 sky130_fd_sc_hd__a22o_1 _6814_ (.A1(_1390_),
    .A2(_0572_),
    .B1(_0771_),
    .B2(_1410_),
    .X(_2264_));
 sky130_fd_sc_hd__or2_1 _6815_ (.A(_1981_),
    .B(_2264_),
    .X(_2265_));
 sky130_fd_sc_hd__inv_2 _6816_ (.A(_1410_),
    .Y(_2266_));
 sky130_fd_sc_hd__nand2_1 _6817_ (.A(_2266_),
    .B(_1900_),
    .Y(_2267_));
 sky130_fd_sc_hd__nand2_1 _6818_ (.A(_1358_),
    .B(_1280_),
    .Y(_2268_));
 sky130_fd_sc_hd__o21ai_1 _6819_ (.A1(_1280_),
    .A2(_1402_),
    .B1(_2268_),
    .Y(_2269_));
 sky130_fd_sc_hd__inv_2 _6820_ (.A(_2269_),
    .Y(_2270_));
 sky130_fd_sc_hd__a22o_1 _6821_ (.A1(_1393_),
    .A2(_1906_),
    .B1(_2270_),
    .B2(_1987_),
    .X(_2271_));
 sky130_fd_sc_hd__a41o_2 _6822_ (.A1(_2263_),
    .A2(_1932_),
    .A3(_2265_),
    .A4(_2267_),
    .B1(_2271_),
    .X(net719));
 sky130_fd_sc_hd__o21ai_1 _6823_ (.A1(_0197_),
    .A2(_1400_),
    .B1(_0209_),
    .Y(_2272_));
 sky130_fd_sc_hd__a22o_2 _6824_ (.A1(_1367_),
    .A2(_2023_),
    .B1(_1372_),
    .B2(_1924_),
    .X(_2273_));
 sky130_fd_sc_hd__a22o_1 _6825_ (.A1(_1436_),
    .A2(_1892_),
    .B1(_1385_),
    .B2(_1953_),
    .X(_2274_));
 sky130_fd_sc_hd__a21o_1 _6826_ (.A1(_2274_),
    .A2(_1941_),
    .B1(_1926_),
    .X(_2275_));
 sky130_fd_sc_hd__nand2_1 _6827_ (.A(_1435_),
    .B(_0844_),
    .Y(_2276_));
 sky130_fd_sc_hd__nand2_1 _6828_ (.A(_1410_),
    .B(_0844_),
    .Y(_2277_));
 sky130_fd_sc_hd__mux2_1 _6829_ (.A0(_2276_),
    .A1(_2277_),
    .S(_0090_),
    .X(_2278_));
 sky130_fd_sc_hd__mux2_1 _6830_ (.A0(_2248_),
    .A1(_2278_),
    .S(_0841_),
    .X(_2279_));
 sky130_fd_sc_hd__nand2_1 _6831_ (.A(_2279_),
    .B(_2004_),
    .Y(_2280_));
 sky130_fd_sc_hd__o221ai_4 _6832_ (.A1(_1435_),
    .A2(_1983_),
    .B1(_2273_),
    .B2(_2275_),
    .C1(_2280_),
    .Y(_2281_));
 sky130_fd_sc_hd__o21ai_1 _6833_ (.A1(_0197_),
    .A2(_2272_),
    .B1(_2281_),
    .Y(_2282_));
 sky130_fd_sc_hd__o21ai_4 _6834_ (.A1(_4100_),
    .A2(_0166_),
    .B1(_0138_),
    .Y(_2283_));
 sky130_fd_sc_hd__nand2_1 _6835_ (.A(_2272_),
    .B(_2283_),
    .Y(_2284_));
 sky130_fd_sc_hd__a22o_1 _6836_ (.A1(_1395_),
    .A2(_1986_),
    .B1(_2282_),
    .B2(_2284_),
    .X(net720));
 sky130_fd_sc_hd__nor2_1 _6837_ (.A(_0862_),
    .B(_1479_),
    .Y(_2285_));
 sky130_fd_sc_hd__a211o_1 _6838_ (.A1(_1413_),
    .A2(_0862_),
    .B1(_1895_),
    .C1(_2285_),
    .X(_2286_));
 sky130_fd_sc_hd__nor2_1 _6839_ (.A(_1973_),
    .B(_1445_),
    .Y(_2287_));
 sky130_fd_sc_hd__o21ai_1 _6840_ (.A1(_1914_),
    .A2(_2287_),
    .B1(_1917_),
    .Y(_2288_));
 sky130_fd_sc_hd__nor2_1 _6841_ (.A(_1920_),
    .B(_1418_),
    .Y(_2289_));
 sky130_fd_sc_hd__a221o_2 _6842_ (.A1(_1422_),
    .A2(_1924_),
    .B1(_2286_),
    .B2(_2288_),
    .C1(_2289_),
    .X(_2290_));
 sky130_fd_sc_hd__nand2_1 _6843_ (.A(_2290_),
    .B(_1929_),
    .Y(_2291_));
 sky130_fd_sc_hd__a22o_1 _6844_ (.A1(_1435_),
    .A2(_0729_),
    .B1(_0730_),
    .B2(_1468_),
    .X(_2292_));
 sky130_fd_sc_hd__inv_2 _6845_ (.A(_2292_),
    .Y(_2293_));
 sky130_fd_sc_hd__nand2_1 _6846_ (.A(_2293_),
    .B(_2004_),
    .Y(_2294_));
 sky130_fd_sc_hd__inv_2 _6847_ (.A(_1468_),
    .Y(_2295_));
 sky130_fd_sc_hd__nand2_1 _6848_ (.A(_2295_),
    .B(_1900_),
    .Y(_2296_));
 sky130_fd_sc_hd__a22o_1 _6849_ (.A1(_1404_),
    .A2(_1906_),
    .B1(_1408_),
    .B2(_1987_),
    .X(_2297_));
 sky130_fd_sc_hd__a41o_2 _6850_ (.A1(_2291_),
    .A2(_1932_),
    .A3(_2294_),
    .A4(_2296_),
    .B1(_2297_),
    .X(net721));
 sky130_fd_sc_hd__nand2_1 _6851_ (.A(_1449_),
    .B(_1997_),
    .Y(_2298_));
 sky130_fd_sc_hd__nor2_1 _6852_ (.A(_1973_),
    .B(_1440_),
    .Y(_2299_));
 sky130_fd_sc_hd__o21ai_1 _6853_ (.A1(_1914_),
    .A2(_2299_),
    .B1(_1917_),
    .Y(_2300_));
 sky130_fd_sc_hd__nor2_1 _6854_ (.A(_1889_),
    .B(_1457_),
    .Y(_2301_));
 sky130_fd_sc_hd__a221o_2 _6855_ (.A1(_1506_),
    .A2(_2023_),
    .B1(_2298_),
    .B2(_2300_),
    .C1(_2301_),
    .X(_2302_));
 sky130_fd_sc_hd__nand2_1 _6856_ (.A(_2302_),
    .B(_1929_),
    .Y(_2303_));
 sky130_fd_sc_hd__a22o_1 _6857_ (.A1(_1468_),
    .A2(_0572_),
    .B1(_0771_),
    .B2(_1512_),
    .X(_2304_));
 sky130_fd_sc_hd__inv_2 _6858_ (.A(_2304_),
    .Y(_2305_));
 sky130_fd_sc_hd__nand2_1 _6859_ (.A(_2305_),
    .B(_2004_),
    .Y(_2306_));
 sky130_fd_sc_hd__inv_2 _6860_ (.A(_1512_),
    .Y(_2307_));
 sky130_fd_sc_hd__nand2_1 _6861_ (.A(_2307_),
    .B(_1900_),
    .Y(_2308_));
 sky130_fd_sc_hd__a22o_1 _6862_ (.A1(_1428_),
    .A2(_1906_),
    .B1(_1433_),
    .B2(_1987_),
    .X(_2309_));
 sky130_fd_sc_hd__a41o_2 _6863_ (.A1(_2303_),
    .A2(_1932_),
    .A3(_2306_),
    .A4(_2308_),
    .B1(_2309_),
    .X(net722));
 sky130_fd_sc_hd__a22o_1 _6864_ (.A1(_1474_),
    .A2(_1955_),
    .B1(_1480_),
    .B2(_1997_),
    .X(_2310_));
 sky130_fd_sc_hd__a22o_1 _6865_ (.A1(_1483_),
    .A2(_2023_),
    .B1(_1488_),
    .B2(_1923_),
    .X(_2311_));
 sky130_fd_sc_hd__a211o_2 _6866_ (.A1(_2310_),
    .A2(_1999_),
    .B1(_1926_),
    .C1(_2311_),
    .X(_2312_));
 sky130_fd_sc_hd__nand2_1 _6867_ (.A(_1535_),
    .B(_0844_),
    .Y(_2313_));
 sky130_fd_sc_hd__nand2_1 _6868_ (.A(_1512_),
    .B(_0844_),
    .Y(_2314_));
 sky130_fd_sc_hd__mux2_1 _6869_ (.A0(_2313_),
    .A1(_2314_),
    .S(_0090_),
    .X(_2315_));
 sky130_fd_sc_hd__mux2_1 _6870_ (.A0(_2293_),
    .A1(_2315_),
    .S(_0841_),
    .X(_2316_));
 sky130_fd_sc_hd__nand2_1 _6871_ (.A(_2316_),
    .B(_2004_),
    .Y(_2317_));
 sky130_fd_sc_hd__o21a_1 _6872_ (.A1(_1983_),
    .A2(_1535_),
    .B1(_1931_),
    .X(_2318_));
 sky130_fd_sc_hd__a22o_1 _6873_ (.A1(_1462_),
    .A2(_1986_),
    .B1(_1466_),
    .B2(_1988_),
    .X(_2319_));
 sky130_fd_sc_hd__a31o_2 _6874_ (.A1(_2312_),
    .A2(_2317_),
    .A3(_2318_),
    .B1(_2319_),
    .X(net723));
 sky130_fd_sc_hd__nand2_1 _6875_ (.A(_1545_),
    .B(_0833_),
    .Y(_2320_));
 sky130_fd_sc_hd__nand3_1 _6876_ (.A(_1505_),
    .B(_2320_),
    .C(_1923_),
    .Y(_2321_));
 sky130_fd_sc_hd__a21o_1 _6877_ (.A1(_1548_),
    .A2(_1892_),
    .B1(_1913_),
    .X(_2322_));
 sky130_fd_sc_hd__a22o_1 _6878_ (.A1(_1916_),
    .A2(_2322_),
    .B1(_1500_),
    .B2(_1939_),
    .X(_2323_));
 sky130_fd_sc_hd__o211a_2 _6879_ (.A1(_1518_),
    .A2(_1920_),
    .B1(_2321_),
    .C1(_2323_),
    .X(_2324_));
 sky130_fd_sc_hd__a22o_1 _6880_ (.A1(_1535_),
    .A2(_0729_),
    .B1(_0771_),
    .B2(_1564_),
    .X(_2325_));
 sky130_fd_sc_hd__inv_2 _6881_ (.A(_2325_),
    .Y(_2326_));
 sky130_fd_sc_hd__nand2_1 _6882_ (.A(_2326_),
    .B(_2003_),
    .Y(_2327_));
 sky130_fd_sc_hd__o221a_1 _6883_ (.A1(_1564_),
    .A2(_1901_),
    .B1(_1926_),
    .B2(_2324_),
    .C1(_2327_),
    .X(_2328_));
 sky130_fd_sc_hd__a31o_1 _6884_ (.A1(_0209_),
    .A2(_0652_),
    .A3(_1562_),
    .B1(_2328_),
    .X(_2329_));
 sky130_fd_sc_hd__o21ai_1 _6885_ (.A1(_0197_),
    .A2(_1562_),
    .B1(_0209_),
    .Y(_2330_));
 sky130_fd_sc_hd__nand2_1 _6886_ (.A(_2330_),
    .B(_2283_),
    .Y(_2331_));
 sky130_fd_sc_hd__a22o_1 _6887_ (.A1(_1539_),
    .A2(_1986_),
    .B1(_2329_),
    .B2(_2331_),
    .X(net724));
 sky130_fd_sc_hd__a22o_1 _6888_ (.A1(_1575_),
    .A2(_1955_),
    .B1(_1529_),
    .B2(_1953_),
    .X(_2332_));
 sky130_fd_sc_hd__nand2_1 _6889_ (.A(_2332_),
    .B(_1999_),
    .Y(_2333_));
 sky130_fd_sc_hd__nand2_1 _6890_ (.A(_1522_),
    .B(_1924_),
    .Y(_2334_));
 sky130_fd_sc_hd__nand2_1 _6891_ (.A(_1515_),
    .B(_2023_),
    .Y(_2335_));
 sky130_fd_sc_hd__or2_1 _6892_ (.A(_0771_),
    .B(_1565_),
    .X(_2336_));
 sky130_fd_sc_hd__o21ai_2 _6893_ (.A1(_0090_),
    .A2(_1607_),
    .B1(_2336_),
    .Y(_2337_));
 sky130_fd_sc_hd__o221ai_4 _6894_ (.A1(_1588_),
    .A2(_1983_),
    .B1(_1981_),
    .B2(_2337_),
    .C1(_1931_),
    .Y(_2338_));
 sky130_fd_sc_hd__a41o_2 _6895_ (.A1(_2333_),
    .A2(_1947_),
    .A3(_2334_),
    .A4(_2335_),
    .B1(_2338_),
    .X(_2339_));
 sky130_fd_sc_hd__a21bo_1 _6896_ (.A1(_1591_),
    .A2(_1911_),
    .B1_N(_2339_),
    .X(net725));
 sky130_fd_sc_hd__inv_2 _6897_ (.A(_1552_),
    .Y(_2340_));
 sky130_fd_sc_hd__a22o_1 _6898_ (.A1(_2340_),
    .A2(_1955_),
    .B1(_1556_),
    .B2(_1953_),
    .X(_2341_));
 sky130_fd_sc_hd__nand2_1 _6899_ (.A(_2341_),
    .B(_1941_),
    .Y(_2342_));
 sky130_fd_sc_hd__nand2_1 _6900_ (.A(_1547_),
    .B(_1924_),
    .Y(_2343_));
 sky130_fd_sc_hd__nand2_1 _6901_ (.A(_1541_),
    .B(_2023_),
    .Y(_2344_));
 sky130_fd_sc_hd__o221ai_4 _6902_ (.A1(_1605_),
    .A2(_1983_),
    .B1(_1902_),
    .B2(_1609_),
    .C1(_1931_),
    .Y(_2345_));
 sky130_fd_sc_hd__a41o_2 _6903_ (.A1(_2342_),
    .A2(_1947_),
    .A3(_2343_),
    .A4(_2344_),
    .B1(_2345_),
    .X(_2346_));
 sky130_fd_sc_hd__a21bo_1 _6904_ (.A1(_1594_),
    .A2(_1911_),
    .B1_N(_2346_),
    .X(net726));
 sky130_fd_sc_hd__a22o_1 _6905_ (.A1(_1539_),
    .A2(_0767_),
    .B1(_0769_),
    .B2(_1591_),
    .X(_2347_));
 sky130_fd_sc_hd__or2_1 _6906_ (.A(_1280_),
    .B(_1642_),
    .X(_2348_));
 sky130_fd_sc_hd__o21ai_2 _6907_ (.A1(_0887_),
    .A2(_2347_),
    .B1(_2348_),
    .Y(_2349_));
 sky130_fd_sc_hd__nand2_1 _6908_ (.A(_1636_),
    .B(_1986_),
    .Y(_2350_));
 sky130_fd_sc_hd__inv_2 _6909_ (.A(_1579_),
    .Y(_2351_));
 sky130_fd_sc_hd__a22o_1 _6910_ (.A1(_2351_),
    .A2(_1955_),
    .B1(_1583_),
    .B2(_1997_),
    .X(_2352_));
 sky130_fd_sc_hd__nand2_1 _6911_ (.A(_2352_),
    .B(_1999_),
    .Y(_2353_));
 sky130_fd_sc_hd__nand2_1 _6912_ (.A(_1574_),
    .B(_1924_),
    .Y(_2354_));
 sky130_fd_sc_hd__nand2_1 _6913_ (.A(_1570_),
    .B(_2023_),
    .Y(_2355_));
 sky130_fd_sc_hd__or2_1 _6914_ (.A(_0771_),
    .B(_1606_),
    .X(_2356_));
 sky130_fd_sc_hd__o21ai_2 _6915_ (.A1(_0090_),
    .A2(_1602_),
    .B1(_2356_),
    .Y(_2357_));
 sky130_fd_sc_hd__o221ai_4 _6916_ (.A1(_1601_),
    .A2(_1983_),
    .B1(_1981_),
    .B2(_2357_),
    .C1(_1931_),
    .Y(_2358_));
 sky130_fd_sc_hd__a41o_2 _6917_ (.A1(_2353_),
    .A2(_1947_),
    .A3(_2354_),
    .A4(_2355_),
    .B1(_2358_),
    .X(_2359_));
 sky130_fd_sc_hd__o211ai_4 _6918_ (.A1(_2349_),
    .A2(_1908_),
    .B1(_2350_),
    .C1(_2359_),
    .Y(net727));
 sky130_fd_sc_hd__nor2_1 _6919_ (.A(_1893_),
    .B(_1621_),
    .Y(_2360_));
 sky130_fd_sc_hd__o21a_1 _6920_ (.A1(_1914_),
    .A2(_2360_),
    .B1(_1917_),
    .X(_2361_));
 sky130_fd_sc_hd__a31o_1 _6921_ (.A1(_1624_),
    .A2(_0589_),
    .A3(_1989_),
    .B1(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__o221a_1 _6922_ (.A1(_1614_),
    .A2(_1920_),
    .B1(_1619_),
    .B2(_1889_),
    .C1(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__or2_1 _6923_ (.A(_1926_),
    .B(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__or2_1 _6924_ (.A(_1981_),
    .B(_1611_),
    .X(_2365_));
 sky130_fd_sc_hd__nand2_1 _6925_ (.A(_1678_),
    .B(_1900_),
    .Y(_2366_));
 sky130_fd_sc_hd__or2_1 _6926_ (.A(_0886_),
    .B(_1596_),
    .X(_2367_));
 sky130_fd_sc_hd__o21ai_1 _6927_ (.A1(_1280_),
    .A2(_1685_),
    .B1(_2367_),
    .Y(_2368_));
 sky130_fd_sc_hd__inv_2 _6928_ (.A(_2368_),
    .Y(_2369_));
 sky130_fd_sc_hd__a22o_1 _6929_ (.A1(_1640_),
    .A2(_1906_),
    .B1(_2369_),
    .B2(_1987_),
    .X(_2370_));
 sky130_fd_sc_hd__a41o_2 _6930_ (.A1(_2364_),
    .A2(_1932_),
    .A3(_2365_),
    .A4(_2366_),
    .B1(_2370_),
    .X(net728));
 sky130_fd_sc_hd__inv_2 _6931_ (.A(_1658_),
    .Y(_2371_));
 sky130_fd_sc_hd__a22o_1 _6932_ (.A1(_2371_),
    .A2(_1955_),
    .B1(_1659_),
    .B2(_1997_),
    .X(_2372_));
 sky130_fd_sc_hd__nor2_1 _6933_ (.A(_1999_),
    .B(_1689_),
    .Y(_2373_));
 sky130_fd_sc_hd__a211o_1 _6934_ (.A1(_2372_),
    .A2(_1999_),
    .B1(_1926_),
    .C1(_2373_),
    .X(_2374_));
 sky130_fd_sc_hd__o21a_1 _6935_ (.A1(_1929_),
    .A2(_1673_),
    .B1(_1931_),
    .X(_2375_));
 sky130_fd_sc_hd__a22o_2 _6936_ (.A1(_1638_),
    .A2(_1911_),
    .B1(_2374_),
    .B2(_2375_),
    .X(net503));
 sky130_fd_sc_hd__and2_1 _6937_ (.A(_1646_),
    .B(_0288_),
    .X(_2376_));
 sky130_fd_sc_hd__a221o_1 _6938_ (.A1(_1717_),
    .A2(_1898_),
    .B1(_2376_),
    .B2(_1891_),
    .C1(_1903_),
    .X(_2377_));
 sky130_fd_sc_hd__o21a_1 _6939_ (.A1(_1670_),
    .A2(_1928_),
    .B1(_2377_),
    .X(_2378_));
 sky130_fd_sc_hd__inv_2 _6940_ (.A(_2283_),
    .Y(_2379_));
 sky130_fd_sc_hd__or2_1 _6941_ (.A(_0197_),
    .B(_1681_),
    .X(_2380_));
 sky130_fd_sc_hd__o211a_1 _6942_ (.A1(_0652_),
    .A2(_2378_),
    .B1(_0209_),
    .C1(_2380_),
    .X(_2381_));
 sky130_fd_sc_hd__a221o_1 _6943_ (.A1(_1681_),
    .A2(_1986_),
    .B1(_2378_),
    .B2(_2379_),
    .C1(_2381_),
    .X(net504));
 sky130_fd_sc_hd__inv_2 _6944_ (.A(_1725_),
    .Y(_2382_));
 sky130_fd_sc_hd__a22o_1 _6945_ (.A1(_1692_),
    .A2(_1891_),
    .B1(_2382_),
    .B2(_1898_),
    .X(_2383_));
 sky130_fd_sc_hd__mux2_1 _6946_ (.A0(_2383_),
    .A1(_1703_),
    .S(_1903_),
    .X(_2384_));
 sky130_fd_sc_hd__or2_1 _6947_ (.A(_0652_),
    .B(_2384_),
    .X(_2385_));
 sky130_fd_sc_hd__nand2_1 _6948_ (.A(_1721_),
    .B(_0652_),
    .Y(_2386_));
 sky130_fd_sc_hd__a22o_1 _6949_ (.A1(_1711_),
    .A2(_1986_),
    .B1(_2384_),
    .B2(_2379_),
    .X(_2387_));
 sky130_fd_sc_hd__a31o_1 _6950_ (.A1(_0209_),
    .A2(_2385_),
    .A3(_2386_),
    .B1(_2387_),
    .X(net505));
 sky130_fd_sc_hd__a22o_1 _6951_ (.A1(_1735_),
    .A2(_1891_),
    .B1(_1738_),
    .B2(_1898_),
    .X(_2388_));
 sky130_fd_sc_hd__mux2_1 _6952_ (.A0(_2388_),
    .A1(_1733_),
    .S(_1904_),
    .X(_2389_));
 sky130_fd_sc_hd__mux2_1 _6953_ (.A0(_2389_),
    .A1(_1742_),
    .S(_1910_),
    .X(_2390_));
 sky130_fd_sc_hd__clkbuf_2 _6954_ (.A(_2390_),
    .X(net506));
 sky130_fd_sc_hd__o21ai_1 _6955_ (.A1(_1973_),
    .A2(_1749_),
    .B1(_1941_),
    .Y(_2391_));
 sky130_fd_sc_hd__a31o_1 _6956_ (.A1(_0520_),
    .A2(_1750_),
    .A3(_1997_),
    .B1(_2391_),
    .X(_2392_));
 sky130_fd_sc_hd__o21ai_1 _6957_ (.A1(_1745_),
    .A2(_1999_),
    .B1(_2392_),
    .Y(_2393_));
 sky130_fd_sc_hd__nand2_1 _6958_ (.A(_2393_),
    .B(_1929_),
    .Y(_2394_));
 sky130_fd_sc_hd__o21a_1 _6959_ (.A1(_1947_),
    .A2(_1753_),
    .B1(_1931_),
    .X(_2395_));
 sky130_fd_sc_hd__a22o_2 _6960_ (.A1(_1756_),
    .A2(_1911_),
    .B1(_2394_),
    .B2(_2395_),
    .X(net507));
 sky130_fd_sc_hd__a22o_1 _6961_ (.A1(_1766_),
    .A2(_1891_),
    .B1(_1764_),
    .B2(_1898_),
    .X(_2396_));
 sky130_fd_sc_hd__mux2_1 _6962_ (.A0(_2396_),
    .A1(_1779_),
    .S(_1904_),
    .X(_2397_));
 sky130_fd_sc_hd__mux2_1 _6963_ (.A0(_2397_),
    .A1(_1762_),
    .S(_1910_),
    .X(_2398_));
 sky130_fd_sc_hd__clkbuf_2 _6964_ (.A(_2398_),
    .X(net508));
 sky130_fd_sc_hd__nor2_1 _6965_ (.A(_0539_),
    .B(_1793_),
    .Y(_2399_));
 sky130_fd_sc_hd__a221o_1 _6966_ (.A1(_1794_),
    .A2(_1892_),
    .B1(_2399_),
    .B2(_1953_),
    .C1(_1891_),
    .X(_2400_));
 sky130_fd_sc_hd__o221a_1 _6967_ (.A1(_1768_),
    .A2(_1920_),
    .B1(_1770_),
    .B2(_1889_),
    .C1(_2400_),
    .X(_2401_));
 sky130_fd_sc_hd__or2_1 _6968_ (.A(_1926_),
    .B(_2401_),
    .X(_2402_));
 sky130_fd_sc_hd__o21a_1 _6969_ (.A1(_1947_),
    .A2(_1801_),
    .B1(_1931_),
    .X(_2403_));
 sky130_fd_sc_hd__a22o_2 _6970_ (.A1(_1788_),
    .A2(_1911_),
    .B1(_2402_),
    .B2(_2403_),
    .X(net509));
 sky130_fd_sc_hd__and2_1 _6971_ (.A(_1772_),
    .B(_0288_),
    .X(_2404_));
 sky130_fd_sc_hd__a221o_1 _6972_ (.A1(_1807_),
    .A2(_1898_),
    .B1(_2404_),
    .B2(_1891_),
    .C1(_1904_),
    .X(_2405_));
 sky130_fd_sc_hd__o21a_1 _6973_ (.A1(_1816_),
    .A2(_1947_),
    .B1(_2405_),
    .X(_2406_));
 sky130_fd_sc_hd__mux2_1 _6974_ (.A0(_2406_),
    .A1(_1784_),
    .S(_1910_),
    .X(_2407_));
 sky130_fd_sc_hd__buf_2 _6975_ (.A(_2407_),
    .X(net510));
 sky130_fd_sc_hd__a22o_1 _6976_ (.A1(_1809_),
    .A2(_1891_),
    .B1(_1822_),
    .B2(_1898_),
    .X(_2408_));
 sky130_fd_sc_hd__mux2_1 _6977_ (.A0(_2408_),
    .A1(_1826_),
    .S(_1904_),
    .X(_2409_));
 sky130_fd_sc_hd__mux2_1 _6978_ (.A0(_2409_),
    .A1(_1786_),
    .S(_1910_),
    .X(_2410_));
 sky130_fd_sc_hd__clkbuf_2 _6979_ (.A(_2410_),
    .X(net511));
 sky130_fd_sc_hd__nor2_2 _6980_ (.A(_0287_),
    .B(_0284_),
    .Y(_2411_));
 sky130_fd_sc_hd__a221o_1 _6981_ (.A1(_0229_),
    .A2(_1898_),
    .B1(_2411_),
    .B2(_1891_),
    .C1(_1904_),
    .X(_2412_));
 sky130_fd_sc_hd__o21a_1 _6982_ (.A1(_0131_),
    .A2(_1947_),
    .B1(_2412_),
    .X(_2413_));
 sky130_fd_sc_hd__mux2_1 _6983_ (.A0(_2413_),
    .A1(_0191_),
    .S(_1910_),
    .X(_2414_));
 sky130_fd_sc_hd__buf_1 _6984_ (.A(_2414_),
    .X(net512));
 sky130_fd_sc_hd__a221o_1 _6985_ (.A1(_1836_),
    .A2(_1891_),
    .B1(_1839_),
    .B2(_1898_),
    .C1(_1904_),
    .X(_2415_));
 sky130_fd_sc_hd__o21a_1 _6986_ (.A1(_1842_),
    .A2(_1947_),
    .B1(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__mux2_1 _6987_ (.A0(_2416_),
    .A1(_1845_),
    .S(_1910_),
    .X(_2417_));
 sky130_fd_sc_hd__clkbuf_2 _6988_ (.A(_2417_),
    .X(net514));
 sky130_fd_sc_hd__and2b_1 _6989_ (.A_N(_1852_),
    .B(_1898_),
    .X(_2418_));
 sky130_fd_sc_hd__a21o_1 _6990_ (.A1(_1855_),
    .A2(_1891_),
    .B1(_2418_),
    .X(_2419_));
 sky130_fd_sc_hd__mux2_1 _6991_ (.A0(_2419_),
    .A1(_1850_),
    .S(_1904_),
    .X(_2420_));
 sky130_fd_sc_hd__mux2_1 _6992_ (.A0(_2420_),
    .A1(_1848_),
    .S(_1910_),
    .X(_2421_));
 sky130_fd_sc_hd__clkbuf_2 _6993_ (.A(_2421_),
    .X(net515));
 sky130_fd_sc_hd__or3_1 _6994_ (.A(_1897_),
    .B(_1891_),
    .C(_1866_),
    .X(_2422_));
 sky130_fd_sc_hd__o21ai_1 _6995_ (.A1(_1864_),
    .A2(_1941_),
    .B1(_2422_),
    .Y(_2423_));
 sky130_fd_sc_hd__mux2_1 _6996_ (.A0(_2423_),
    .A1(_1869_),
    .S(_1904_),
    .X(_2424_));
 sky130_fd_sc_hd__mux2_1 _6997_ (.A0(_2424_),
    .A1(_1873_),
    .S(_1910_),
    .X(_2425_));
 sky130_fd_sc_hd__clkbuf_2 _6998_ (.A(_2425_),
    .X(net516));
 sky130_fd_sc_hd__a22o_1 _6999_ (.A1(_1878_),
    .A2(_1891_),
    .B1(_1881_),
    .B2(_1898_),
    .X(_2426_));
 sky130_fd_sc_hd__mux2_1 _7000_ (.A0(_2426_),
    .A1(_1876_),
    .S(_1904_),
    .X(_2427_));
 sky130_fd_sc_hd__mux2_1 _7001_ (.A0(_2427_),
    .A1(_1885_),
    .S(_1910_),
    .X(_2428_));
 sky130_fd_sc_hd__clkbuf_2 _7002_ (.A(_2428_),
    .X(net517));
 sky130_fd_sc_hd__a22o_4 _7003_ (.A1(_4235_),
    .A2(_4098_),
    .B1(_4278_),
    .B2(_4233_),
    .X(_2429_));
 sky130_fd_sc_hd__buf_6 _7004_ (.A(_2429_),
    .X(_2430_));
 sky130_fd_sc_hd__inv_2 _7005_ (.A(_2429_),
    .Y(_2431_));
 sky130_fd_sc_hd__a22o_1 _7006_ (.A1(_0538_),
    .A2(_0588_),
    .B1(_4112_),
    .B2(_4098_),
    .X(_2432_));
 sky130_fd_sc_hd__and2_1 _7007_ (.A(_2431_),
    .B(_2432_),
    .X(_2433_));
 sky130_fd_sc_hd__buf_4 _7008_ (.A(_2433_),
    .X(_2434_));
 sky130_fd_sc_hd__a22o_1 _7009_ (.A1(_0416_),
    .A2(_2430_),
    .B1(_0439_),
    .B2(_2434_),
    .X(_2435_));
 sky130_fd_sc_hd__a22o_4 _7010_ (.A1(_0759_),
    .A2(_4239_),
    .B1(_4241_),
    .B2(_4098_),
    .X(_2436_));
 sky130_fd_sc_hd__buf_8 _7011_ (.A(_2436_),
    .X(_2437_));
 sky130_fd_sc_hd__mux2_1 _7012_ (.A0(_2435_),
    .A1(_0459_),
    .S(_2437_),
    .X(_2438_));
 sky130_fd_sc_hd__clkbuf_16 _7013_ (.A(_0741_),
    .X(_2439_));
 sky130_fd_sc_hd__a22o_1 _7014_ (.A1(_2439_),
    .A2(_0209_),
    .B1(_0168_),
    .B2(_4098_),
    .X(_2440_));
 sky130_fd_sc_hd__buf_6 _7015_ (.A(_2440_),
    .X(_2441_));
 sky130_fd_sc_hd__buf_8 _7016_ (.A(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__mux2_4 _7017_ (.A0(_2438_),
    .A1(_0482_),
    .S(_2442_),
    .X(_2443_));
 sky130_fd_sc_hd__buf_1 _7018_ (.A(_2443_),
    .X(net502));
 sky130_fd_sc_hd__buf_8 _7019_ (.A(_2429_),
    .X(_2444_));
 sky130_fd_sc_hd__clkbuf_8 _7020_ (.A(_2434_),
    .X(_2445_));
 sky130_fd_sc_hd__a221o_1 _7021_ (.A1(_0494_),
    .A2(_2444_),
    .B1(_0499_),
    .B2(_2445_),
    .C1(_2437_),
    .X(_2446_));
 sky130_fd_sc_hd__inv_6 _7022_ (.A(_2436_),
    .Y(_2447_));
 sky130_fd_sc_hd__clkbuf_8 _7023_ (.A(_2447_),
    .X(_2448_));
 sky130_fd_sc_hd__o21ba_1 _7024_ (.A1(_2448_),
    .A2(_0502_),
    .B1_N(_2441_),
    .X(_2449_));
 sky130_fd_sc_hd__a22o_2 _7025_ (.A1(_0505_),
    .A2(_2442_),
    .B1(_2446_),
    .B2(_2449_),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_8 _7026_ (.A(_2447_),
    .X(_2450_));
 sky130_fd_sc_hd__and2_1 _7027_ (.A(_0519_),
    .B(_2445_),
    .X(_2451_));
 sky130_fd_sc_hd__a21o_1 _7028_ (.A1(_0508_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2452_));
 sky130_fd_sc_hd__o22a_1 _7029_ (.A1(_0530_),
    .A2(_2450_),
    .B1(_2451_),
    .B2(_2452_),
    .X(_2453_));
 sky130_fd_sc_hd__mux2_4 _7030_ (.A0(_2453_),
    .A1(_0533_),
    .S(_2442_),
    .X(_2454_));
 sky130_fd_sc_hd__buf_1 _7031_ (.A(_2454_),
    .X(net652));
 sky130_fd_sc_hd__and2_1 _7032_ (.A(_1954_),
    .B(_2445_),
    .X(_2455_));
 sky130_fd_sc_hd__a21o_1 _7033_ (.A1(_0553_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2456_));
 sky130_fd_sc_hd__o22a_1 _7034_ (.A1(_0537_),
    .A2(_2450_),
    .B1(_2455_),
    .B2(_2456_),
    .X(_2457_));
 sky130_fd_sc_hd__mux2_4 _7035_ (.A0(_2457_),
    .A1(_0565_),
    .S(_2442_),
    .X(_2458_));
 sky130_fd_sc_hd__buf_1 _7036_ (.A(_2458_),
    .X(net663));
 sky130_fd_sc_hd__nor2_1 _7037_ (.A(_0287_),
    .B(_0595_),
    .Y(_2459_));
 sky130_fd_sc_hd__a221o_1 _7038_ (.A1(_0586_),
    .A2(_2434_),
    .B1(_2459_),
    .B2(_2429_),
    .C1(_2436_),
    .X(_2460_));
 sky130_fd_sc_hd__o21ai_1 _7039_ (.A1(_0571_),
    .A2(_2447_),
    .B1(_2460_),
    .Y(_2461_));
 sky130_fd_sc_hd__inv_2 _7040_ (.A(_2461_),
    .Y(_2462_));
 sky130_fd_sc_hd__mux2_4 _7041_ (.A0(_2462_),
    .A1(_0569_),
    .S(_2442_),
    .X(_2463_));
 sky130_fd_sc_hd__buf_1 _7042_ (.A(_2463_),
    .X(net674));
 sky130_fd_sc_hd__nor2_1 _7043_ (.A(_0287_),
    .B(_1967_),
    .Y(_2464_));
 sky130_fd_sc_hd__a221o_1 _7044_ (.A1(_0609_),
    .A2(_2434_),
    .B1(_2464_),
    .B2(_2429_),
    .C1(_2436_),
    .X(_2465_));
 sky130_fd_sc_hd__o21ai_2 _7045_ (.A1(_0574_),
    .A2(_2447_),
    .B1(_2465_),
    .Y(_2466_));
 sky130_fd_sc_hd__inv_2 _7046_ (.A(_2466_),
    .Y(_2467_));
 sky130_fd_sc_hd__mux2_1 _7047_ (.A0(_2467_),
    .A1(_0648_),
    .S(_2442_),
    .X(_2468_));
 sky130_fd_sc_hd__buf_1 _7048_ (.A(_2468_),
    .X(net685));
 sky130_fd_sc_hd__o21ai_1 _7049_ (.A1(_2431_),
    .A2(_0617_),
    .B1(_2447_),
    .Y(_2469_));
 sky130_fd_sc_hd__and2b_1 _7050_ (.A_N(net730),
    .B(_2445_),
    .X(_2470_));
 sky130_fd_sc_hd__o22a_1 _7051_ (.A1(_0576_),
    .A2(_2450_),
    .B1(_2469_),
    .B2(_2470_),
    .X(_2471_));
 sky130_fd_sc_hd__mux2_1 _7052_ (.A0(_2471_),
    .A1(_0656_),
    .S(_2442_),
    .X(_2472_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _7053_ (.A(_2472_),
    .X(net696));
 sky130_fd_sc_hd__o21ai_1 _7054_ (.A1(_2431_),
    .A2(_0619_),
    .B1(_2447_),
    .Y(_2473_));
 sky130_fd_sc_hd__and2_1 _7055_ (.A(_0676_),
    .B(_2445_),
    .X(_2474_));
 sky130_fd_sc_hd__o22a_1 _7056_ (.A1(_0639_),
    .A2(_2450_),
    .B1(_2473_),
    .B2(_2474_),
    .X(_2475_));
 sky130_fd_sc_hd__mux2_1 _7057_ (.A0(_2475_),
    .A1(_0650_),
    .S(_2442_),
    .X(_2476_));
 sky130_fd_sc_hd__buf_1 _7058_ (.A(_2476_),
    .X(net707));
 sky130_fd_sc_hd__buf_6 _7059_ (.A(_2429_),
    .X(_2477_));
 sky130_fd_sc_hd__buf_6 _7060_ (.A(_2434_),
    .X(_2478_));
 sky130_fd_sc_hd__buf_8 _7061_ (.A(_2436_),
    .X(_2479_));
 sky130_fd_sc_hd__a221o_1 _7062_ (.A1(_0715_),
    .A2(_2477_),
    .B1(_0693_),
    .B2(_2478_),
    .C1(_2479_),
    .X(_2480_));
 sky130_fd_sc_hd__o21a_1 _7063_ (.A1(_0727_),
    .A2(_2448_),
    .B1(_2480_),
    .X(_2481_));
 sky130_fd_sc_hd__mux2_1 _7064_ (.A0(_2481_),
    .A1(_0688_),
    .S(_2442_),
    .X(_2482_));
 sky130_fd_sc_hd__buf_1 _7065_ (.A(_2482_),
    .X(net718));
 sky130_fd_sc_hd__a221o_1 _7066_ (.A1(_0710_),
    .A2(_2477_),
    .B1(_0698_),
    .B2(_2478_),
    .C1(_2479_),
    .X(_2483_));
 sky130_fd_sc_hd__o21a_1 _7067_ (.A1(_0739_),
    .A2(_2448_),
    .B1(_2483_),
    .X(_2484_));
 sky130_fd_sc_hd__mux2_1 _7068_ (.A0(_2484_),
    .A1(_0736_),
    .S(_2442_),
    .X(_2485_));
 sky130_fd_sc_hd__buf_1 _7069_ (.A(_2485_),
    .X(net729));
 sky130_fd_sc_hd__a21o_1 _7070_ (.A1(_0712_),
    .A2(_2477_),
    .B1(_2479_),
    .X(_2486_));
 sky130_fd_sc_hd__and2_1 _7071_ (.A(_0701_),
    .B(_2445_),
    .X(_2487_));
 sky130_fd_sc_hd__o22a_1 _7072_ (.A1(_0752_),
    .A2(_2450_),
    .B1(_2486_),
    .B2(_2487_),
    .X(_2488_));
 sky130_fd_sc_hd__mux2_1 _7073_ (.A0(_2488_),
    .A1(_0746_),
    .S(_2442_),
    .X(_2489_));
 sky130_fd_sc_hd__buf_1 _7074_ (.A(_2489_),
    .X(net513));
 sky130_fd_sc_hd__a221o_1 _7075_ (.A1(_0780_),
    .A2(_2477_),
    .B1(_0819_),
    .B2(_2478_),
    .C1(_2479_),
    .X(_2490_));
 sky130_fd_sc_hd__o21a_1 _7076_ (.A1(_0754_),
    .A2(_2448_),
    .B1(_2490_),
    .X(_2491_));
 sky130_fd_sc_hd__mux2_1 _7077_ (.A0(_2491_),
    .A1(_0765_),
    .S(_2442_),
    .X(_2492_));
 sky130_fd_sc_hd__buf_1 _7078_ (.A(_2492_),
    .X(net524));
 sky130_fd_sc_hd__a221o_1 _7079_ (.A1(_0788_),
    .A2(_2477_),
    .B1(_0808_),
    .B2(_2478_),
    .C1(_2479_),
    .X(_2493_));
 sky130_fd_sc_hd__o21a_1 _7080_ (.A1(_0756_),
    .A2(_2448_),
    .B1(_2493_),
    .X(_2494_));
 sky130_fd_sc_hd__mux2_1 _7081_ (.A0(_2494_),
    .A1(_0854_),
    .S(_2442_),
    .X(_2495_));
 sky130_fd_sc_hd__buf_1 _7082_ (.A(_2495_),
    .X(net535));
 sky130_fd_sc_hd__and2_1 _7083_ (.A(_0826_),
    .B(_2445_),
    .X(_2496_));
 sky130_fd_sc_hd__a21o_1 _7084_ (.A1(_0784_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2497_));
 sky130_fd_sc_hd__o22a_1 _7085_ (.A1(_0773_),
    .A2(_2450_),
    .B1(_2496_),
    .B2(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__mux2_1 _7086_ (.A0(_2498_),
    .A1(_0885_),
    .S(_2442_),
    .X(_2499_));
 sky130_fd_sc_hd__buf_1 _7087_ (.A(_2499_),
    .X(net546));
 sky130_fd_sc_hd__buf_6 _7088_ (.A(_2434_),
    .X(_2500_));
 sky130_fd_sc_hd__clkbuf_8 _7089_ (.A(_2436_),
    .X(_2501_));
 sky130_fd_sc_hd__a221o_1 _7090_ (.A1(_0628_),
    .A2(_2477_),
    .B1(_0863_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2502_));
 sky130_fd_sc_hd__o21a_1 _7091_ (.A1(_0843_),
    .A2(_2448_),
    .B1(_2502_),
    .X(_2503_));
 sky130_fd_sc_hd__mux2_1 _7092_ (.A0(_2503_),
    .A1(_0896_),
    .S(_2442_),
    .X(_2504_));
 sky130_fd_sc_hd__buf_1 _7093_ (.A(_2504_),
    .X(net557));
 sky130_fd_sc_hd__inv_2 _7094_ (.A(_0867_),
    .Y(_2505_));
 sky130_fd_sc_hd__a221o_1 _7095_ (.A1(_0906_),
    .A2(_2430_),
    .B1(_2505_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2506_));
 sky130_fd_sc_hd__o21a_1 _7096_ (.A1(_0877_),
    .A2(_2448_),
    .B1(_2506_),
    .X(_2507_));
 sky130_fd_sc_hd__mux2_1 _7097_ (.A0(_2507_),
    .A1(_0893_),
    .S(_2442_),
    .X(_2508_));
 sky130_fd_sc_hd__buf_1 _7098_ (.A(_2508_),
    .X(net568));
 sky130_fd_sc_hd__and2_1 _7099_ (.A(_0948_),
    .B(_2445_),
    .X(_2509_));
 sky130_fd_sc_hd__a21o_1 _7100_ (.A1(_0904_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2510_));
 sky130_fd_sc_hd__o22a_1 _7101_ (.A1(_0955_),
    .A2(_2450_),
    .B1(_2509_),
    .B2(_2510_),
    .X(_2511_));
 sky130_fd_sc_hd__buf_6 _7102_ (.A(_2441_),
    .X(_2512_));
 sky130_fd_sc_hd__mux2_1 _7103_ (.A0(_2511_),
    .A1(_0940_),
    .S(_2512_),
    .X(_2513_));
 sky130_fd_sc_hd__buf_1 _7104_ (.A(_2513_),
    .X(net579));
 sky130_fd_sc_hd__and2_1 _7105_ (.A(_0957_),
    .B(_2445_),
    .X(_2514_));
 sky130_fd_sc_hd__a21o_1 _7106_ (.A1(_0944_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2515_));
 sky130_fd_sc_hd__o22a_2 _7107_ (.A1(_0980_),
    .A2(_2450_),
    .B1(_2514_),
    .B2(_2515_),
    .X(_2516_));
 sky130_fd_sc_hd__mux2_1 _7108_ (.A0(_2516_),
    .A1(_0983_),
    .S(_2512_),
    .X(_2517_));
 sky130_fd_sc_hd__buf_1 _7109_ (.A(_2517_),
    .X(net590));
 sky130_fd_sc_hd__and2_1 _7110_ (.A(_2118_),
    .B(_2445_),
    .X(_2518_));
 sky130_fd_sc_hd__a21o_1 _7111_ (.A1(_0942_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2519_));
 sky130_fd_sc_hd__o22a_2 _7112_ (.A1(_1014_),
    .A2(_2450_),
    .B1(_2518_),
    .B2(_2519_),
    .X(_2520_));
 sky130_fd_sc_hd__mux2_1 _7113_ (.A0(_2520_),
    .A1(_0986_),
    .S(_2512_),
    .X(_2521_));
 sky130_fd_sc_hd__buf_1 _7114_ (.A(_2521_),
    .X(net601));
 sky130_fd_sc_hd__and2_1 _7115_ (.A(_1025_),
    .B(_2478_),
    .X(_2522_));
 sky130_fd_sc_hd__a21o_1 _7116_ (.A1(_0973_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2523_));
 sky130_fd_sc_hd__o22a_1 _7117_ (.A1(_1019_),
    .A2(_2450_),
    .B1(_2522_),
    .B2(_2523_),
    .X(_2524_));
 sky130_fd_sc_hd__mux2_2 _7118_ (.A0(_2524_),
    .A1(_1017_),
    .S(_2512_),
    .X(_2525_));
 sky130_fd_sc_hd__buf_1 _7119_ (.A(_2525_),
    .X(net612));
 sky130_fd_sc_hd__inv_2 _7120_ (.A(_1034_),
    .Y(_2526_));
 sky130_fd_sc_hd__and2_1 _7121_ (.A(_2526_),
    .B(_2478_),
    .X(_2527_));
 sky130_fd_sc_hd__a21o_1 _7122_ (.A1(_0990_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2528_));
 sky130_fd_sc_hd__o22a_1 _7123_ (.A1(_1064_),
    .A2(_2450_),
    .B1(_2527_),
    .B2(_2528_),
    .X(_2529_));
 sky130_fd_sc_hd__mux2_2 _7124_ (.A0(_2529_),
    .A1(_1050_),
    .S(_2512_),
    .X(_2530_));
 sky130_fd_sc_hd__buf_1 _7125_ (.A(_2530_),
    .X(net624));
 sky130_fd_sc_hd__a221o_1 _7126_ (.A1(_1021_),
    .A2(_2430_),
    .B1(_1068_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2531_));
 sky130_fd_sc_hd__o21a_1 _7127_ (.A1(_1077_),
    .A2(_2448_),
    .B1(_2531_),
    .X(_2532_));
 sky130_fd_sc_hd__mux2_1 _7128_ (.A0(_2532_),
    .A1(_1067_),
    .S(_2512_),
    .X(_2533_));
 sky130_fd_sc_hd__buf_1 _7129_ (.A(_2533_),
    .X(net635));
 sky130_fd_sc_hd__a221o_2 _7130_ (.A1(_1052_),
    .A2(_2430_),
    .B1(_1099_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2534_));
 sky130_fd_sc_hd__o21a_1 _7131_ (.A1(_1081_),
    .A2(_2448_),
    .B1(_2534_),
    .X(_2535_));
 sky130_fd_sc_hd__mux2_1 _7132_ (.A0(_2535_),
    .A1(_1106_),
    .S(_2512_),
    .X(_2536_));
 sky130_fd_sc_hd__buf_1 _7133_ (.A(_2536_),
    .X(net644));
 sky130_fd_sc_hd__a221o_2 _7134_ (.A1(_1071_),
    .A2(_2430_),
    .B1(_1112_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2537_));
 sky130_fd_sc_hd__o21a_1 _7135_ (.A1(_1083_),
    .A2(_2448_),
    .B1(_2537_),
    .X(_2538_));
 sky130_fd_sc_hd__mux2_1 _7136_ (.A0(_2538_),
    .A1(_1153_),
    .S(_2512_),
    .X(_2539_));
 sky130_fd_sc_hd__buf_1 _7137_ (.A(_2539_),
    .X(net645));
 sky130_fd_sc_hd__buf_8 _7138_ (.A(_2447_),
    .X(_2540_));
 sky130_fd_sc_hd__and2_1 _7139_ (.A(_1174_),
    .B(_2478_),
    .X(_2541_));
 sky130_fd_sc_hd__a21o_1 _7140_ (.A1(_1090_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2542_));
 sky130_fd_sc_hd__o22a_2 _7141_ (.A1(_1144_),
    .A2(_2540_),
    .B1(_2541_),
    .B2(_2542_),
    .X(_2543_));
 sky130_fd_sc_hd__mux2_1 _7142_ (.A0(_2543_),
    .A1(_1158_),
    .S(_2512_),
    .X(_2544_));
 sky130_fd_sc_hd__buf_1 _7143_ (.A(_2544_),
    .X(net646));
 sky130_fd_sc_hd__a221o_1 _7144_ (.A1(_0995_),
    .A2(_2430_),
    .B1(_1117_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2545_));
 sky130_fd_sc_hd__o21a_1 _7145_ (.A1(_1141_),
    .A2(_2448_),
    .B1(_2545_),
    .X(_2546_));
 sky130_fd_sc_hd__mux2_1 _7146_ (.A0(_2546_),
    .A1(_1155_),
    .S(_2512_),
    .X(_2547_));
 sky130_fd_sc_hd__buf_1 _7147_ (.A(_2547_),
    .X(net647));
 sky130_fd_sc_hd__and2_1 _7148_ (.A(_1223_),
    .B(_2478_),
    .X(_2548_));
 sky130_fd_sc_hd__a21o_1 _7149_ (.A1(_0997_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2549_));
 sky130_fd_sc_hd__o22a_2 _7150_ (.A1(_1213_),
    .A2(_2540_),
    .B1(_2548_),
    .B2(_2549_),
    .X(_2550_));
 sky130_fd_sc_hd__mux2_1 _7151_ (.A0(_2550_),
    .A1(_1169_),
    .S(_2512_),
    .X(_2551_));
 sky130_fd_sc_hd__buf_1 _7152_ (.A(_2551_),
    .X(net648));
 sky130_fd_sc_hd__and2_1 _7153_ (.A(_2193_),
    .B(_2478_),
    .X(_2552_));
 sky130_fd_sc_hd__a21o_1 _7154_ (.A1(_1000_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2553_));
 sky130_fd_sc_hd__o22a_2 _7155_ (.A1(_1215_),
    .A2(_2540_),
    .B1(_2552_),
    .B2(_2553_),
    .X(_2554_));
 sky130_fd_sc_hd__mux2_1 _7156_ (.A0(_2554_),
    .A1(_1232_),
    .S(_2512_),
    .X(_2555_));
 sky130_fd_sc_hd__buf_1 _7157_ (.A(_2555_),
    .X(net649));
 sky130_fd_sc_hd__a221o_2 _7158_ (.A1(_1002_),
    .A2(_2430_),
    .B1(_1257_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2556_));
 sky130_fd_sc_hd__o21a_1 _7159_ (.A1(_1277_),
    .A2(_2448_),
    .B1(_2556_),
    .X(_2557_));
 sky130_fd_sc_hd__mux2_1 _7160_ (.A0(_2557_),
    .A1(_1256_),
    .S(_2512_),
    .X(_2558_));
 sky130_fd_sc_hd__buf_1 _7161_ (.A(_2558_),
    .X(net650));
 sky130_fd_sc_hd__a221o_2 _7162_ (.A1(_1246_),
    .A2(_2430_),
    .B1(_1294_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2559_));
 sky130_fd_sc_hd__o21a_1 _7163_ (.A1(_1304_),
    .A2(_2448_),
    .B1(_2559_),
    .X(_2560_));
 sky130_fd_sc_hd__mux2_1 _7164_ (.A0(_2560_),
    .A1(_1282_),
    .S(_2512_),
    .X(_2561_));
 sky130_fd_sc_hd__buf_1 _7165_ (.A(_2561_),
    .X(net651));
 sky130_fd_sc_hd__a21o_1 _7166_ (.A1(_1269_),
    .A2(_2477_),
    .B1(_2479_),
    .X(_2562_));
 sky130_fd_sc_hd__and2_1 _7167_ (.A(_1260_),
    .B(_2445_),
    .X(_2563_));
 sky130_fd_sc_hd__o22a_2 _7168_ (.A1(_1299_),
    .A2(_2540_),
    .B1(_2562_),
    .B2(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__mux2_2 _7169_ (.A0(_2564_),
    .A1(_1284_),
    .S(_2512_),
    .X(_2565_));
 sky130_fd_sc_hd__buf_1 _7170_ (.A(_2565_),
    .X(net653));
 sky130_fd_sc_hd__inv_2 _7171_ (.A(_1322_),
    .Y(_2566_));
 sky130_fd_sc_hd__and2_1 _7172_ (.A(_2566_),
    .B(_2478_),
    .X(_2567_));
 sky130_fd_sc_hd__a21o_1 _7173_ (.A1(_1335_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2568_));
 sky130_fd_sc_hd__o22a_2 _7174_ (.A1(_1301_),
    .A2(_2540_),
    .B1(_2567_),
    .B2(_2568_),
    .X(_2569_));
 sky130_fd_sc_hd__mux2_1 _7175_ (.A0(_2569_),
    .A1(_1333_),
    .S(_2512_),
    .X(_2570_));
 sky130_fd_sc_hd__buf_1 _7176_ (.A(_2570_),
    .X(net654));
 sky130_fd_sc_hd__and2_1 _7177_ (.A(_1373_),
    .B(_2478_),
    .X(_2571_));
 sky130_fd_sc_hd__a21o_1 _7178_ (.A1(_1347_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2572_));
 sky130_fd_sc_hd__o22a_2 _7179_ (.A1(_1390_),
    .A2(_2540_),
    .B1(_2571_),
    .B2(_2572_),
    .X(_2573_));
 sky130_fd_sc_hd__clkbuf_8 _7180_ (.A(_2441_),
    .X(_2574_));
 sky130_fd_sc_hd__mux2_1 _7181_ (.A0(_2573_),
    .A1(_1361_),
    .S(_2574_),
    .X(_2575_));
 sky130_fd_sc_hd__buf_1 _7182_ (.A(_2575_),
    .X(net655));
 sky130_fd_sc_hd__and2_1 _7183_ (.A(_1415_),
    .B(_2478_),
    .X(_2576_));
 sky130_fd_sc_hd__a21o_1 _7184_ (.A1(_1345_),
    .A2(_2444_),
    .B1(_2437_),
    .X(_2577_));
 sky130_fd_sc_hd__o22a_2 _7185_ (.A1(_1410_),
    .A2(_2540_),
    .B1(_2576_),
    .B2(_2577_),
    .X(_2578_));
 sky130_fd_sc_hd__mux2_4 _7186_ (.A0(_2578_),
    .A1(_1393_),
    .S(_2574_),
    .X(_2579_));
 sky130_fd_sc_hd__buf_1 _7187_ (.A(_2579_),
    .X(net656));
 sky130_fd_sc_hd__a221o_1 _7188_ (.A1(_1367_),
    .A2(_2430_),
    .B1(_1436_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2580_));
 sky130_fd_sc_hd__o21a_1 _7189_ (.A1(_1435_),
    .A2(_2448_),
    .B1(_2580_),
    .X(_2581_));
 sky130_fd_sc_hd__mux2_2 _7190_ (.A0(_2581_),
    .A1(_1395_),
    .S(_2574_),
    .X(_2582_));
 sky130_fd_sc_hd__buf_1 _7191_ (.A(_2582_),
    .X(net657));
 sky130_fd_sc_hd__and2_1 _7192_ (.A(_1469_),
    .B(_2478_),
    .X(_2583_));
 sky130_fd_sc_hd__a21o_1 _7193_ (.A1(_1418_),
    .A2(_2444_),
    .B1(_2479_),
    .X(_2584_));
 sky130_fd_sc_hd__o22a_2 _7194_ (.A1(_1468_),
    .A2(_2540_),
    .B1(_2583_),
    .B2(_2584_),
    .X(_2585_));
 sky130_fd_sc_hd__mux2_2 _7195_ (.A0(_2585_),
    .A1(_1404_),
    .S(_2574_),
    .X(_2586_));
 sky130_fd_sc_hd__buf_1 _7196_ (.A(_2586_),
    .X(net658));
 sky130_fd_sc_hd__a221o_2 _7197_ (.A1(_1452_),
    .A2(_2430_),
    .B1(_1502_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2587_));
 sky130_fd_sc_hd__o21a_1 _7198_ (.A1(_1512_),
    .A2(_2448_),
    .B1(_2587_),
    .X(_2588_));
 sky130_fd_sc_hd__mux2_2 _7199_ (.A0(_2588_),
    .A1(_1428_),
    .S(_2574_),
    .X(_2589_));
 sky130_fd_sc_hd__buf_1 _7200_ (.A(_2589_),
    .X(net659));
 sky130_fd_sc_hd__a221o_2 _7201_ (.A1(_1483_),
    .A2(_2430_),
    .B1(_1474_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2590_));
 sky130_fd_sc_hd__o21a_1 _7202_ (.A1(_1535_),
    .A2(_2448_),
    .B1(_2590_),
    .X(_2591_));
 sky130_fd_sc_hd__mux2_2 _7203_ (.A0(_2591_),
    .A1(_1462_),
    .S(_2574_),
    .X(_2592_));
 sky130_fd_sc_hd__buf_1 _7204_ (.A(_2592_),
    .X(net660));
 sky130_fd_sc_hd__a221o_1 _7205_ (.A1(_1518_),
    .A2(_2430_),
    .B1(_1548_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2593_));
 sky130_fd_sc_hd__o21a_1 _7206_ (.A1(_1564_),
    .A2(_2450_),
    .B1(_2593_),
    .X(_2594_));
 sky130_fd_sc_hd__mux2_2 _7207_ (.A0(_2594_),
    .A1(_1539_),
    .S(_2574_),
    .X(_2595_));
 sky130_fd_sc_hd__buf_1 _7208_ (.A(_2595_),
    .X(net661));
 sky130_fd_sc_hd__and2_1 _7209_ (.A(_1575_),
    .B(_2478_),
    .X(_2596_));
 sky130_fd_sc_hd__a21o_1 _7210_ (.A1(_1515_),
    .A2(_2477_),
    .B1(_2479_),
    .X(_2597_));
 sky130_fd_sc_hd__o22a_2 _7211_ (.A1(_1588_),
    .A2(_2540_),
    .B1(_2596_),
    .B2(_2597_),
    .X(_2598_));
 sky130_fd_sc_hd__mux2_2 _7212_ (.A0(_2598_),
    .A1(_1591_),
    .S(_2574_),
    .X(_2599_));
 sky130_fd_sc_hd__buf_1 _7213_ (.A(_2599_),
    .X(net662));
 sky130_fd_sc_hd__a221o_1 _7214_ (.A1(_1541_),
    .A2(_2430_),
    .B1(_2340_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2600_));
 sky130_fd_sc_hd__o21a_1 _7215_ (.A1(_1605_),
    .A2(_2450_),
    .B1(_2600_),
    .X(_2601_));
 sky130_fd_sc_hd__mux2_2 _7216_ (.A0(_2601_),
    .A1(_1594_),
    .S(_2574_),
    .X(_2602_));
 sky130_fd_sc_hd__buf_1 _7217_ (.A(_2602_),
    .X(net664));
 sky130_fd_sc_hd__and2_1 _7218_ (.A(_2351_),
    .B(_2478_),
    .X(_2603_));
 sky130_fd_sc_hd__a21o_1 _7219_ (.A1(_1570_),
    .A2(_2477_),
    .B1(_2479_),
    .X(_2604_));
 sky130_fd_sc_hd__o22a_2 _7220_ (.A1(_1601_),
    .A2(_2540_),
    .B1(_2603_),
    .B2(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__mux2_2 _7221_ (.A0(_2605_),
    .A1(_1636_),
    .S(_2574_),
    .X(_2606_));
 sky130_fd_sc_hd__buf_1 _7222_ (.A(_2606_),
    .X(net665));
 sky130_fd_sc_hd__a21o_1 _7223_ (.A1(_1614_),
    .A2(_2477_),
    .B1(_2479_),
    .X(_2607_));
 sky130_fd_sc_hd__and2b_1 _7224_ (.A_N(_1621_),
    .B(_2445_),
    .X(_2608_));
 sky130_fd_sc_hd__o22a_1 _7225_ (.A1(_1598_),
    .A2(_2540_),
    .B1(_2607_),
    .B2(_2608_),
    .X(_2609_));
 sky130_fd_sc_hd__mux2_2 _7226_ (.A0(_2609_),
    .A1(_1640_),
    .S(_2574_),
    .X(_2610_));
 sky130_fd_sc_hd__buf_1 _7227_ (.A(_2610_),
    .X(net666));
 sky130_fd_sc_hd__a221o_1 _7228_ (.A1(_1649_),
    .A2(_2430_),
    .B1(_2371_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2611_));
 sky130_fd_sc_hd__o21a_1 _7229_ (.A1(_1673_),
    .A2(_2450_),
    .B1(_2611_),
    .X(_2612_));
 sky130_fd_sc_hd__mux2_2 _7230_ (.A0(_2612_),
    .A1(_1638_),
    .S(_2574_),
    .X(_2613_));
 sky130_fd_sc_hd__buf_1 _7231_ (.A(_2613_),
    .X(net667));
 sky130_fd_sc_hd__a221o_1 _7232_ (.A1(_1717_),
    .A2(_2434_),
    .B1(_2376_),
    .B2(_2429_),
    .C1(_2436_),
    .X(_2614_));
 sky130_fd_sc_hd__o21ai_2 _7233_ (.A1(_1670_),
    .A2(_2447_),
    .B1(_2614_),
    .Y(_2615_));
 sky130_fd_sc_hd__inv_2 _7234_ (.A(_2615_),
    .Y(_2616_));
 sky130_fd_sc_hd__mux2_2 _7235_ (.A0(_2616_),
    .A1(_1681_),
    .S(_2574_),
    .X(_2617_));
 sky130_fd_sc_hd__buf_1 _7236_ (.A(_2617_),
    .X(net668));
 sky130_fd_sc_hd__a221o_1 _7237_ (.A1(_1692_),
    .A2(_2430_),
    .B1(_2382_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2618_));
 sky130_fd_sc_hd__o21a_1 _7238_ (.A1(_1703_),
    .A2(_2450_),
    .B1(_2618_),
    .X(_2619_));
 sky130_fd_sc_hd__mux2_2 _7239_ (.A0(_2619_),
    .A1(_1711_),
    .S(_2574_),
    .X(_2620_));
 sky130_fd_sc_hd__buf_1 _7240_ (.A(_2620_),
    .X(net669));
 sky130_fd_sc_hd__a21o_1 _7241_ (.A1(_1735_),
    .A2(_2477_),
    .B1(_2479_),
    .X(_2621_));
 sky130_fd_sc_hd__and2_1 _7242_ (.A(_1738_),
    .B(_2445_),
    .X(_2622_));
 sky130_fd_sc_hd__o22a_1 _7243_ (.A1(_1733_),
    .A2(_2540_),
    .B1(_2621_),
    .B2(_2622_),
    .X(_2623_));
 sky130_fd_sc_hd__mux2_4 _7244_ (.A0(_2623_),
    .A1(_1742_),
    .S(_2574_),
    .X(_2624_));
 sky130_fd_sc_hd__buf_1 _7245_ (.A(_2624_),
    .X(net670));
 sky130_fd_sc_hd__and2_1 _7246_ (.A(_1750_),
    .B(_2478_),
    .X(_2625_));
 sky130_fd_sc_hd__a21o_1 _7247_ (.A1(_1745_),
    .A2(_2477_),
    .B1(_2479_),
    .X(_2626_));
 sky130_fd_sc_hd__o22a_1 _7248_ (.A1(_1753_),
    .A2(_2540_),
    .B1(_2625_),
    .B2(_2626_),
    .X(_2627_));
 sky130_fd_sc_hd__mux2_2 _7249_ (.A0(_2627_),
    .A1(_1756_),
    .S(_2574_),
    .X(_2628_));
 sky130_fd_sc_hd__buf_1 _7250_ (.A(_2628_),
    .X(net671));
 sky130_fd_sc_hd__nor2_1 _7251_ (.A(_0287_),
    .B(_1775_),
    .Y(_2629_));
 sky130_fd_sc_hd__a221o_1 _7252_ (.A1(_2629_),
    .A2(_2429_),
    .B1(_1764_),
    .B2(_2434_),
    .C1(_2436_),
    .X(_2630_));
 sky130_fd_sc_hd__o21ai_1 _7253_ (.A1(_1779_),
    .A2(_2447_),
    .B1(_2630_),
    .Y(_2631_));
 sky130_fd_sc_hd__inv_2 _7254_ (.A(_2631_),
    .Y(_2632_));
 sky130_fd_sc_hd__mux2_2 _7255_ (.A0(_2632_),
    .A1(_1762_),
    .S(_2441_),
    .X(_2633_));
 sky130_fd_sc_hd__buf_1 _7256_ (.A(_2633_),
    .X(net672));
 sky130_fd_sc_hd__a221o_1 _7257_ (.A1(_1768_),
    .A2(_2430_),
    .B1(_1794_),
    .B2(_2500_),
    .C1(_2501_),
    .X(_2634_));
 sky130_fd_sc_hd__o21a_1 _7258_ (.A1(_1801_),
    .A2(_2450_),
    .B1(_2634_),
    .X(_2635_));
 sky130_fd_sc_hd__mux2_2 _7259_ (.A0(_2635_),
    .A1(_1788_),
    .S(_2441_),
    .X(_2636_));
 sky130_fd_sc_hd__buf_1 _7260_ (.A(_2636_),
    .X(net673));
 sky130_fd_sc_hd__a221o_1 _7261_ (.A1(_1807_),
    .A2(_2434_),
    .B1(_2404_),
    .B2(_2429_),
    .C1(_2436_),
    .X(_2637_));
 sky130_fd_sc_hd__o21ai_1 _7262_ (.A1(_1816_),
    .A2(_2447_),
    .B1(_2637_),
    .Y(_2638_));
 sky130_fd_sc_hd__inv_2 _7263_ (.A(_2638_),
    .Y(_2639_));
 sky130_fd_sc_hd__mux2_4 _7264_ (.A0(_2639_),
    .A1(_1784_),
    .S(_2441_),
    .X(_2640_));
 sky130_fd_sc_hd__buf_1 _7265_ (.A(_2640_),
    .X(net675));
 sky130_fd_sc_hd__and2_1 _7266_ (.A(_1809_),
    .B(_0288_),
    .X(_2641_));
 sky130_fd_sc_hd__a221o_1 _7267_ (.A1(_1822_),
    .A2(_2434_),
    .B1(_2641_),
    .B2(_2429_),
    .C1(_2436_),
    .X(_2642_));
 sky130_fd_sc_hd__o21ai_1 _7268_ (.A1(_1826_),
    .A2(_2447_),
    .B1(_2642_),
    .Y(_2643_));
 sky130_fd_sc_hd__inv_2 _7269_ (.A(_2643_),
    .Y(_2644_));
 sky130_fd_sc_hd__mux2_2 _7270_ (.A0(_2644_),
    .A1(_1786_),
    .S(_2441_),
    .X(_2645_));
 sky130_fd_sc_hd__buf_1 _7271_ (.A(_2645_),
    .X(net676));
 sky130_fd_sc_hd__and3_1 _7272_ (.A(_2431_),
    .B(_0229_),
    .C(_2432_),
    .X(_2646_));
 sky130_fd_sc_hd__a21o_1 _7273_ (.A1(_0041_),
    .A2(_2477_),
    .B1(_2479_),
    .X(_2647_));
 sky130_fd_sc_hd__o22a_1 _7274_ (.A1(_0131_),
    .A2(_2540_),
    .B1(_2646_),
    .B2(_2647_),
    .X(_2648_));
 sky130_fd_sc_hd__mux2_1 _7275_ (.A0(_2648_),
    .A1(_0191_),
    .S(_2441_),
    .X(_2649_));
 sky130_fd_sc_hd__buf_1 _7276_ (.A(_2649_),
    .X(net677));
 sky130_fd_sc_hd__a21o_1 _7277_ (.A1(_1836_),
    .A2(_2477_),
    .B1(_2479_),
    .X(_2650_));
 sky130_fd_sc_hd__and2_1 _7278_ (.A(_1839_),
    .B(_2445_),
    .X(_2651_));
 sky130_fd_sc_hd__o22a_1 _7279_ (.A1(_1842_),
    .A2(_2540_),
    .B1(_2650_),
    .B2(_2651_),
    .X(_2652_));
 sky130_fd_sc_hd__mux2_2 _7280_ (.A0(_2652_),
    .A1(_1845_),
    .S(_2441_),
    .X(_2653_));
 sky130_fd_sc_hd__buf_1 _7281_ (.A(_2653_),
    .X(net678));
 sky130_fd_sc_hd__a21o_1 _7282_ (.A1(_1855_),
    .A2(_2477_),
    .B1(_2479_),
    .X(_2654_));
 sky130_fd_sc_hd__and2b_1 _7283_ (.A_N(_1852_),
    .B(_2445_),
    .X(_2655_));
 sky130_fd_sc_hd__o22a_1 _7284_ (.A1(_1850_),
    .A2(_2540_),
    .B1(_2654_),
    .B2(_2655_),
    .X(_2656_));
 sky130_fd_sc_hd__mux2_4 _7285_ (.A0(_2656_),
    .A1(_1848_),
    .S(_2441_),
    .X(_2657_));
 sky130_fd_sc_hd__buf_1 _7286_ (.A(_2657_),
    .X(net679));
 sky130_fd_sc_hd__a21o_1 _7287_ (.A1(_1863_),
    .A2(_2477_),
    .B1(_2479_),
    .X(_2658_));
 sky130_fd_sc_hd__and2b_1 _7288_ (.A_N(_1866_),
    .B(_2445_),
    .X(_2659_));
 sky130_fd_sc_hd__o22a_1 _7289_ (.A1(_1869_),
    .A2(_2447_),
    .B1(_2658_),
    .B2(_2659_),
    .X(_2660_));
 sky130_fd_sc_hd__mux2_2 _7290_ (.A0(_2660_),
    .A1(_1873_),
    .S(_2441_),
    .X(_2661_));
 sky130_fd_sc_hd__buf_1 _7291_ (.A(_2661_),
    .X(net680));
 sky130_fd_sc_hd__a221o_1 _7292_ (.A1(_1879_),
    .A2(_2429_),
    .B1(_1881_),
    .B2(_2434_),
    .C1(_2436_),
    .X(_2662_));
 sky130_fd_sc_hd__o21ai_1 _7293_ (.A1(_1876_),
    .A2(_2447_),
    .B1(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__inv_2 _7294_ (.A(_2663_),
    .Y(_2664_));
 sky130_fd_sc_hd__mux2_2 _7295_ (.A0(_2664_),
    .A1(_1885_),
    .S(_2441_),
    .X(_2665_));
 sky130_fd_sc_hd__buf_1 _7296_ (.A(_2665_),
    .X(net681));
 sky130_fd_sc_hd__nor2_8 _7297_ (.A(_4094_),
    .B(_0056_),
    .Y(_2666_));
 sky130_fd_sc_hd__clkinv_4 _7298_ (.A(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__nand2_8 _7299_ (.A(_0612_),
    .B(_4233_),
    .Y(_2668_));
 sky130_fd_sc_hd__nand2_8 _7300_ (.A(_2667_),
    .B(_2668_),
    .Y(_2669_));
 sky130_fd_sc_hd__buf_6 _7301_ (.A(_2669_),
    .X(_2670_));
 sky130_fd_sc_hd__nor2_8 _7302_ (.A(_4094_),
    .B(_0440_),
    .Y(_2671_));
 sky130_fd_sc_hd__inv_2 _7303_ (.A(_2671_),
    .Y(_2672_));
 sky130_fd_sc_hd__nand2_4 _7304_ (.A(_4186_),
    .B(_0588_),
    .Y(_2673_));
 sky130_fd_sc_hd__nand2_2 _7305_ (.A(_2672_),
    .B(_2673_),
    .Y(_2674_));
 sky130_fd_sc_hd__inv_2 _7306_ (.A(_2674_),
    .Y(_2675_));
 sky130_fd_sc_hd__nor2_8 _7307_ (.A(_2669_),
    .B(_2675_),
    .Y(_2676_));
 sky130_fd_sc_hd__a22o_1 _7308_ (.A1(_0416_),
    .A2(_2670_),
    .B1(_0439_),
    .B2(_2676_),
    .X(_2677_));
 sky130_fd_sc_hd__nor2_8 _7309_ (.A(_4094_),
    .B(_0134_),
    .Y(_2678_));
 sky130_fd_sc_hd__inv_4 _7310_ (.A(_2678_),
    .Y(_2679_));
 sky130_fd_sc_hd__nand2_8 _7311_ (.A(_0111_),
    .B(_4239_),
    .Y(_2680_));
 sky130_fd_sc_hd__nand2_4 _7312_ (.A(_2679_),
    .B(_2680_),
    .Y(_2681_));
 sky130_fd_sc_hd__clkbuf_8 _7313_ (.A(_2681_),
    .X(_2682_));
 sky130_fd_sc_hd__mux2_1 _7314_ (.A0(_2677_),
    .A1(_0459_),
    .S(_2682_),
    .X(_2683_));
 sky130_fd_sc_hd__nand2_2 _7315_ (.A(_0168_),
    .B(_4095_),
    .Y(_2684_));
 sky130_fd_sc_hd__nand2_8 _7316_ (.A(_0766_),
    .B(\arbiter.state[3][1] ),
    .Y(_2685_));
 sky130_fd_sc_hd__nand2_8 _7317_ (.A(_2684_),
    .B(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__mux2_1 _7318_ (.A0(_2683_),
    .A1(_0482_),
    .S(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__clkbuf_2 _7319_ (.A(_2687_),
    .X(net518));
 sky130_fd_sc_hd__a22o_1 _7320_ (.A1(_0494_),
    .A2(_2669_),
    .B1(_0499_),
    .B2(_2676_),
    .X(_2688_));
 sky130_fd_sc_hd__mux2_1 _7321_ (.A0(_2688_),
    .A1(_0502_),
    .S(_2682_),
    .X(_2689_));
 sky130_fd_sc_hd__mux2_1 _7322_ (.A0(_2689_),
    .A1(_0505_),
    .S(_2686_),
    .X(_2690_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _7323_ (.A(_2690_),
    .X(net519));
 sky130_fd_sc_hd__inv_2 _7324_ (.A(_2681_),
    .Y(_2691_));
 sky130_fd_sc_hd__buf_8 _7325_ (.A(_2691_),
    .X(_2692_));
 sky130_fd_sc_hd__buf_6 _7326_ (.A(_2692_),
    .X(_2693_));
 sky130_fd_sc_hd__a221o_1 _7327_ (.A1(_0519_),
    .A2(_2676_),
    .B1(_0508_),
    .B2(_2670_),
    .C1(_2682_),
    .X(_2694_));
 sky130_fd_sc_hd__o21ai_4 _7328_ (.A1(_0530_),
    .A2(_2693_),
    .B1(_2694_),
    .Y(_2695_));
 sky130_fd_sc_hd__inv_2 _7329_ (.A(_2686_),
    .Y(_2696_));
 sky130_fd_sc_hd__clkbuf_8 _7330_ (.A(_2696_),
    .X(_2697_));
 sky130_fd_sc_hd__buf_8 _7331_ (.A(_2697_),
    .X(_2698_));
 sky130_fd_sc_hd__nor2_1 _7332_ (.A(_2698_),
    .B(_0533_),
    .Y(_2699_));
 sky130_fd_sc_hd__a21oi_4 _7333_ (.A1(_2695_),
    .A2(_2698_),
    .B1(_2699_),
    .Y(net520));
 sky130_fd_sc_hd__clkbuf_8 _7334_ (.A(_2691_),
    .X(_2700_));
 sky130_fd_sc_hd__a221o_1 _7335_ (.A1(_0553_),
    .A2(_2670_),
    .B1(_1954_),
    .B2(_2676_),
    .C1(_2681_),
    .X(_2701_));
 sky130_fd_sc_hd__o21a_1 _7336_ (.A1(_0537_),
    .A2(_2700_),
    .B1(_2701_),
    .X(_2702_));
 sky130_fd_sc_hd__mux2_1 _7337_ (.A0(_2702_),
    .A1(_0565_),
    .S(_2686_),
    .X(_2703_));
 sky130_fd_sc_hd__clkbuf_2 _7338_ (.A(_2703_),
    .X(net521));
 sky130_fd_sc_hd__a221o_1 _7339_ (.A1(_0586_),
    .A2(_2676_),
    .B1(_2459_),
    .B2(_2670_),
    .C1(_2682_),
    .X(_2704_));
 sky130_fd_sc_hd__o21ai_1 _7340_ (.A1(_0571_),
    .A2(_2693_),
    .B1(_2704_),
    .Y(_2705_));
 sky130_fd_sc_hd__nor2_1 _7341_ (.A(_2697_),
    .B(_0569_),
    .Y(_2706_));
 sky130_fd_sc_hd__a21oi_2 _7342_ (.A1(_2705_),
    .A2(_2698_),
    .B1(_2706_),
    .Y(net522));
 sky130_fd_sc_hd__a221o_1 _7343_ (.A1(_0609_),
    .A2(_2676_),
    .B1(_2464_),
    .B2(_2670_),
    .C1(_2682_),
    .X(_2707_));
 sky130_fd_sc_hd__o21ai_1 _7344_ (.A1(_0574_),
    .A2(_2693_),
    .B1(_2707_),
    .Y(_2708_));
 sky130_fd_sc_hd__nor2_1 _7345_ (.A(_2697_),
    .B(_0648_),
    .Y(_2709_));
 sky130_fd_sc_hd__a21oi_2 _7346_ (.A1(_2708_),
    .A2(_2698_),
    .B1(_2709_),
    .Y(net523));
 sky130_fd_sc_hd__inv_6 _7347_ (.A(_2669_),
    .Y(_2710_));
 sky130_fd_sc_hd__buf_6 _7348_ (.A(_2710_),
    .X(_2711_));
 sky130_fd_sc_hd__inv_2 _7349_ (.A(_2676_),
    .Y(_2712_));
 sky130_fd_sc_hd__o22a_1 _7350_ (.A1(_0617_),
    .A2(_2711_),
    .B1(_2712_),
    .B2(net730),
    .X(_2713_));
 sky130_fd_sc_hd__mux2_1 _7351_ (.A0(_2713_),
    .A1(_0577_),
    .S(_2682_),
    .X(_2714_));
 sky130_fd_sc_hd__nor2_1 _7352_ (.A(_2697_),
    .B(_0656_),
    .Y(_2715_));
 sky130_fd_sc_hd__a21oi_2 _7353_ (.A1(_2714_),
    .A2(_2698_),
    .B1(_2715_),
    .Y(net525));
 sky130_fd_sc_hd__o22a_1 _7354_ (.A1(_0619_),
    .A2(_2711_),
    .B1(_2712_),
    .B2(_0675_),
    .X(_2716_));
 sky130_fd_sc_hd__mux2_1 _7355_ (.A0(_2716_),
    .A1(_0640_),
    .S(_2682_),
    .X(_2717_));
 sky130_fd_sc_hd__nor2_1 _7356_ (.A(_2697_),
    .B(_0650_),
    .Y(_2718_));
 sky130_fd_sc_hd__a21oi_2 _7357_ (.A1(_2717_),
    .A2(_2698_),
    .B1(_2718_),
    .Y(net526));
 sky130_fd_sc_hd__inv_2 _7358_ (.A(_2685_),
    .Y(_2719_));
 sky130_fd_sc_hd__clkbuf_8 _7359_ (.A(_2719_),
    .X(_2720_));
 sky130_fd_sc_hd__inv_2 _7360_ (.A(_2680_),
    .Y(_2721_));
 sky130_fd_sc_hd__clkbuf_8 _7361_ (.A(_2721_),
    .X(_2722_));
 sky130_fd_sc_hd__inv_2 _7362_ (.A(_2668_),
    .Y(_2723_));
 sky130_fd_sc_hd__buf_6 _7363_ (.A(_2723_),
    .X(_2724_));
 sky130_fd_sc_hd__inv_6 _7364_ (.A(_2673_),
    .Y(_2725_));
 sky130_fd_sc_hd__a22o_1 _7365_ (.A1(_0693_),
    .A2(_2671_),
    .B1(_2013_),
    .B2(_2725_),
    .X(_2726_));
 sky130_fd_sc_hd__nor2_1 _7366_ (.A(_2667_),
    .B(_2001_),
    .Y(_2727_));
 sky130_fd_sc_hd__a221o_1 _7367_ (.A1(_2020_),
    .A2(_2724_),
    .B1(_2726_),
    .B2(_2710_),
    .C1(_2727_),
    .X(_2728_));
 sky130_fd_sc_hd__nor2_1 _7368_ (.A(_2679_),
    .B(_0728_),
    .Y(_2729_));
 sky130_fd_sc_hd__a221o_1 _7369_ (.A1(_2026_),
    .A2(_2722_),
    .B1(_2728_),
    .B2(_2692_),
    .C1(_2729_),
    .X(_2730_));
 sky130_fd_sc_hd__clkbuf_8 _7370_ (.A(_4094_),
    .X(_2731_));
 sky130_fd_sc_hd__o21ai_1 _7371_ (.A1(_2731_),
    .A2(_0688_),
    .B1(_1757_),
    .Y(_2732_));
 sky130_fd_sc_hd__nand2_8 _7372_ (.A(_2685_),
    .B(_0483_),
    .Y(_2733_));
 sky130_fd_sc_hd__buf_4 _7373_ (.A(_2733_),
    .X(_2734_));
 sky130_fd_sc_hd__nand2_1 _7374_ (.A(_2732_),
    .B(_2734_),
    .Y(_2735_));
 sky130_fd_sc_hd__buf_8 _7375_ (.A(_2731_),
    .X(_2736_));
 sky130_fd_sc_hd__nor2_1 _7376_ (.A(_2736_),
    .B(_2732_),
    .Y(_2737_));
 sky130_fd_sc_hd__a221o_2 _7377_ (.A1(_2011_),
    .A2(_2720_),
    .B1(_2730_),
    .B2(_2735_),
    .C1(_2737_),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_8 _7378_ (.A(_4094_),
    .X(_2738_));
 sky130_fd_sc_hd__o21ai_2 _7379_ (.A1(_2738_),
    .A2(_0736_),
    .B1(_0168_),
    .Y(_2739_));
 sky130_fd_sc_hd__nand2_1 _7380_ (.A(_2043_),
    .B(_2720_),
    .Y(_2740_));
 sky130_fd_sc_hd__clkbuf_16 _7381_ (.A(_2667_),
    .X(_2741_));
 sky130_fd_sc_hd__clkbuf_16 _7382_ (.A(_2668_),
    .X(_2742_));
 sky130_fd_sc_hd__nand2_1 _7383_ (.A(_0698_),
    .B(_2671_),
    .Y(_2743_));
 sky130_fd_sc_hd__nand2_2 _7384_ (.A(_4235_),
    .B(_4094_),
    .Y(_2744_));
 sky130_fd_sc_hd__inv_2 _7385_ (.A(_2744_),
    .Y(_2745_));
 sky130_fd_sc_hd__a31o_1 _7386_ (.A1(_2743_),
    .A2(_0056_),
    .A3(_2668_),
    .B1(_2745_),
    .X(_2746_));
 sky130_fd_sc_hd__a21bo_1 _7387_ (.A1(_0705_),
    .A2(_2725_),
    .B1_N(_2746_),
    .X(_2747_));
 sky130_fd_sc_hd__o221ai_4 _7388_ (.A1(_0710_),
    .A2(_2741_),
    .B1(_0720_),
    .B2(_2742_),
    .C1(_2747_),
    .Y(_2748_));
 sky130_fd_sc_hd__clkbuf_8 _7389_ (.A(_2678_),
    .X(_2749_));
 sky130_fd_sc_hd__a22o_1 _7390_ (.A1(_2025_),
    .A2(_2749_),
    .B1(_2739_),
    .B2(_2733_),
    .X(_2750_));
 sky130_fd_sc_hd__a221o_1 _7391_ (.A1(_2037_),
    .A2(_2722_),
    .B1(_2748_),
    .B2(_2700_),
    .C1(_2750_),
    .X(_2751_));
 sky130_fd_sc_hd__o211ai_4 _7392_ (.A1(_2736_),
    .A2(_2739_),
    .B1(_2740_),
    .C1(_2751_),
    .Y(net528));
 sky130_fd_sc_hd__a2bb2o_1 _7393_ (.A1_N(_1007_),
    .A2_N(_0811_),
    .B1(_0701_),
    .B2(_2671_),
    .X(_2752_));
 sky130_fd_sc_hd__nor2_1 _7394_ (.A(_2668_),
    .B(_2046_),
    .Y(_2753_));
 sky130_fd_sc_hd__a221o_1 _7395_ (.A1(_0712_),
    .A2(_2666_),
    .B1(_2752_),
    .B2(_2710_),
    .C1(_2753_),
    .X(_2754_));
 sky130_fd_sc_hd__nor2_1 _7396_ (.A(_2680_),
    .B(_2054_),
    .Y(_2755_));
 sky130_fd_sc_hd__a221o_1 _7397_ (.A1(_0752_),
    .A2(_2749_),
    .B1(_2754_),
    .B2(_2692_),
    .C1(_2755_),
    .X(_2756_));
 sky130_fd_sc_hd__buf_4 _7398_ (.A(_0168_),
    .X(_2757_));
 sky130_fd_sc_hd__o21ai_1 _7399_ (.A1(_2731_),
    .A2(_0746_),
    .B1(_2757_),
    .Y(_2758_));
 sky130_fd_sc_hd__nand2_1 _7400_ (.A(_2758_),
    .B(_2734_),
    .Y(_2759_));
 sky130_fd_sc_hd__nor2_1 _7401_ (.A(_2736_),
    .B(_2758_),
    .Y(_2760_));
 sky130_fd_sc_hd__a221o_2 _7402_ (.A1(_2059_),
    .A2(_2720_),
    .B1(_2756_),
    .B2(_2759_),
    .C1(_2760_),
    .X(net529));
 sky130_fd_sc_hd__o221a_1 _7403_ (.A1(_0797_),
    .A2(_2672_),
    .B1(_1007_),
    .B2(_0820_),
    .C1(_2710_),
    .X(_2761_));
 sky130_fd_sc_hd__o21ai_1 _7404_ (.A1(_2741_),
    .A2(_0780_),
    .B1(_2691_),
    .Y(_2762_));
 sky130_fd_sc_hd__a211oi_2 _7405_ (.A1(_2065_),
    .A2(_2724_),
    .B1(_2761_),
    .C1(_2762_),
    .Y(_2763_));
 sky130_fd_sc_hd__a221o_1 _7406_ (.A1(_0754_),
    .A2(_2749_),
    .B1(_0762_),
    .B2(_2722_),
    .C1(_2763_),
    .X(_2764_));
 sky130_fd_sc_hd__o21ai_1 _7407_ (.A1(_2731_),
    .A2(_0765_),
    .B1(_2757_),
    .Y(_2765_));
 sky130_fd_sc_hd__nand2_1 _7408_ (.A(_2765_),
    .B(_2734_),
    .Y(_2766_));
 sky130_fd_sc_hd__nor2_1 _7409_ (.A(_2736_),
    .B(_2765_),
    .Y(_2767_));
 sky130_fd_sc_hd__a221o_2 _7410_ (.A1(_0858_),
    .A2(_2720_),
    .B1(_2764_),
    .B2(_2766_),
    .C1(_2767_),
    .X(net530));
 sky130_fd_sc_hd__buf_6 _7411_ (.A(_2671_),
    .X(_2768_));
 sky130_fd_sc_hd__a22o_1 _7412_ (.A1(_0808_),
    .A2(_2768_),
    .B1(_0814_),
    .B2(_2725_),
    .X(_2769_));
 sky130_fd_sc_hd__and2_1 _7413_ (.A(_0788_),
    .B(_2666_),
    .X(_2770_));
 sky130_fd_sc_hd__a221o_1 _7414_ (.A1(_0793_),
    .A2(_2724_),
    .B1(_2769_),
    .B2(_2711_),
    .C1(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__nor2_1 _7415_ (.A(_2679_),
    .B(_0851_),
    .Y(_2772_));
 sky130_fd_sc_hd__a221o_1 _7416_ (.A1(_0776_),
    .A2(_2722_),
    .B1(_2771_),
    .B2(_2700_),
    .C1(_2772_),
    .X(_2773_));
 sky130_fd_sc_hd__o21ai_1 _7417_ (.A1(_2738_),
    .A2(_0854_),
    .B1(_2757_),
    .Y(_2774_));
 sky130_fd_sc_hd__nand2_1 _7418_ (.A(_2774_),
    .B(_2734_),
    .Y(_2775_));
 sky130_fd_sc_hd__a2bb2o_1 _7419_ (.A1_N(_2731_),
    .A2_N(_2774_),
    .B1(_2719_),
    .B2(_0891_),
    .X(_2776_));
 sky130_fd_sc_hd__a21o_1 _7420_ (.A1(_2773_),
    .A2(_2775_),
    .B1(_2776_),
    .X(net531));
 sky130_fd_sc_hd__a22o_1 _7421_ (.A1(_0826_),
    .A2(_2671_),
    .B1(_0829_),
    .B2(_2725_),
    .X(_2777_));
 sky130_fd_sc_hd__and2_1 _7422_ (.A(_0784_),
    .B(_2666_),
    .X(_2778_));
 sky130_fd_sc_hd__a221o_1 _7423_ (.A1(_0836_),
    .A2(_2724_),
    .B1(_2777_),
    .B2(_2710_),
    .C1(_2778_),
    .X(_2779_));
 sky130_fd_sc_hd__and2_1 _7424_ (.A(_0848_),
    .B(_2721_),
    .X(_2780_));
 sky130_fd_sc_hd__a221o_1 _7425_ (.A1(_0773_),
    .A2(_2749_),
    .B1(_2779_),
    .B2(_2692_),
    .C1(_2780_),
    .X(_2781_));
 sky130_fd_sc_hd__o21ai_1 _7426_ (.A1(_2738_),
    .A2(_0885_),
    .B1(_2757_),
    .Y(_2782_));
 sky130_fd_sc_hd__nand2_1 _7427_ (.A(_2782_),
    .B(_2734_),
    .Y(_2783_));
 sky130_fd_sc_hd__nor2_1 _7428_ (.A(_2736_),
    .B(_2782_),
    .Y(_2784_));
 sky130_fd_sc_hd__a221o_2 _7429_ (.A1(_2081_),
    .A2(_2720_),
    .B1(_2781_),
    .B2(_2783_),
    .C1(_2784_),
    .X(net532));
 sky130_fd_sc_hd__o221a_1 _7430_ (.A1(_0843_),
    .A2(_2679_),
    .B1(_2680_),
    .B2(_0880_),
    .C1(_2697_),
    .X(_2785_));
 sky130_fd_sc_hd__or3_1 _7431_ (.A(_1007_),
    .B(_1133_),
    .C(_0825_),
    .X(_2786_));
 sky130_fd_sc_hd__nor2_1 _7432_ (.A(_2672_),
    .B(_0825_),
    .Y(_2787_));
 sky130_fd_sc_hd__a21oi_1 _7433_ (.A1(_0629_),
    .A2(_4233_),
    .B1(_0287_),
    .Y(_2788_));
 sky130_fd_sc_hd__o21ai_1 _7434_ (.A1(_2787_),
    .A2(_2788_),
    .B1(_2744_),
    .Y(_2789_));
 sky130_fd_sc_hd__a2bb2o_1 _7435_ (.A1_N(_0628_),
    .A2_N(_2711_),
    .B1(_2786_),
    .B2(_2789_),
    .X(_2790_));
 sky130_fd_sc_hd__nand2_1 _7436_ (.A(_2790_),
    .B(_2693_),
    .Y(_2791_));
 sky130_fd_sc_hd__a22o_1 _7437_ (.A1(_0896_),
    .A2(_2686_),
    .B1(_2785_),
    .B2(_2791_),
    .X(net533));
 sky130_fd_sc_hd__a22o_1 _7438_ (.A1(_2505_),
    .A2(_2671_),
    .B1(_0917_),
    .B2(_0588_),
    .X(_2792_));
 sky130_fd_sc_hd__nor2_1 _7439_ (.A(_2741_),
    .B(_0925_),
    .Y(_2793_));
 sky130_fd_sc_hd__a221o_1 _7440_ (.A1(_2792_),
    .A2(_2711_),
    .B1(_0907_),
    .B2(_2724_),
    .C1(_2793_),
    .X(_2794_));
 sky130_fd_sc_hd__nor2_1 _7441_ (.A(_2679_),
    .B(_2090_),
    .Y(_2795_));
 sky130_fd_sc_hd__a221o_1 _7442_ (.A1(_2103_),
    .A2(_2722_),
    .B1(_2794_),
    .B2(_2700_),
    .C1(_2795_),
    .X(_2796_));
 sky130_fd_sc_hd__o21ai_1 _7443_ (.A1(_2731_),
    .A2(_0893_),
    .B1(_1757_),
    .Y(_2797_));
 sky130_fd_sc_hd__nand2_1 _7444_ (.A(_2797_),
    .B(_2734_),
    .Y(_2798_));
 sky130_fd_sc_hd__o22ai_1 _7445_ (.A1(_2736_),
    .A2(_2797_),
    .B1(_2685_),
    .B2(_2096_),
    .Y(_2799_));
 sky130_fd_sc_hd__a21o_1 _7446_ (.A1(_2796_),
    .A2(_2798_),
    .B1(_2799_),
    .X(net534));
 sky130_fd_sc_hd__inv_2 _7447_ (.A(_2733_),
    .Y(_2800_));
 sky130_fd_sc_hd__o21a_1 _7448_ (.A1(_2731_),
    .A2(_0940_),
    .B1(_1757_),
    .X(_2801_));
 sky130_fd_sc_hd__nor2_1 _7449_ (.A(_2800_),
    .B(_2801_),
    .Y(_2802_));
 sky130_fd_sc_hd__nand2_1 _7450_ (.A(_0931_),
    .B(_2725_),
    .Y(_2803_));
 sky130_fd_sc_hd__nand2_1 _7451_ (.A(_0948_),
    .B(_2768_),
    .Y(_2804_));
 sky130_fd_sc_hd__o221ai_2 _7452_ (.A1(_0904_),
    .A2(_2741_),
    .B1(_2742_),
    .B2(_0971_),
    .C1(_2692_),
    .Y(_2805_));
 sky130_fd_sc_hd__a31o_1 _7453_ (.A1(_2711_),
    .A2(_2803_),
    .A3(_2804_),
    .B1(_2805_),
    .X(_2806_));
 sky130_fd_sc_hd__o221a_1 _7454_ (.A1(_2102_),
    .A2(_2679_),
    .B1(_2109_),
    .B2(_2680_),
    .C1(_2806_),
    .X(_2807_));
 sky130_fd_sc_hd__a2bb2o_1 _7455_ (.A1_N(_2802_),
    .A2_N(_2807_),
    .B1(_0940_),
    .B2(_2686_),
    .X(net536));
 sky130_fd_sc_hd__a22o_1 _7456_ (.A1(_0957_),
    .A2(_2768_),
    .B1(_1008_),
    .B2(_2725_),
    .X(_2808_));
 sky130_fd_sc_hd__a22o_1 _7457_ (.A1(_0944_),
    .A2(_2666_),
    .B1(_2808_),
    .B2(_2711_),
    .X(_2809_));
 sky130_fd_sc_hd__a21o_1 _7458_ (.A1(_0947_),
    .A2(_2724_),
    .B1(_2809_),
    .X(_2810_));
 sky130_fd_sc_hd__nand2_1 _7459_ (.A(_0980_),
    .B(_2749_),
    .Y(_2811_));
 sky130_fd_sc_hd__o21ai_1 _7460_ (.A1(_2680_),
    .A2(_2126_),
    .B1(_2811_),
    .Y(_2812_));
 sky130_fd_sc_hd__a21o_1 _7461_ (.A1(_2810_),
    .A2(_2693_),
    .B1(_2812_),
    .X(_2813_));
 sky130_fd_sc_hd__o21ai_1 _7462_ (.A1(_2731_),
    .A2(_0983_),
    .B1(_1757_),
    .Y(_2814_));
 sky130_fd_sc_hd__nand2_1 _7463_ (.A(_2814_),
    .B(_2734_),
    .Y(_2815_));
 sky130_fd_sc_hd__a22o_1 _7464_ (.A1(_0983_),
    .A2(_2686_),
    .B1(_2813_),
    .B2(_2815_),
    .X(net537));
 sky130_fd_sc_hd__o21ai_1 _7465_ (.A1(_2731_),
    .A2(_0986_),
    .B1(_2757_),
    .Y(_2816_));
 sky130_fd_sc_hd__and2_1 _7466_ (.A(_2816_),
    .B(_2733_),
    .X(_2817_));
 sky130_fd_sc_hd__a22o_1 _7467_ (.A1(_2118_),
    .A2(_2768_),
    .B1(_0969_),
    .B2(_2725_),
    .X(_2818_));
 sky130_fd_sc_hd__nand2_1 _7468_ (.A(_2818_),
    .B(_2711_),
    .Y(_2819_));
 sky130_fd_sc_hd__o221a_1 _7469_ (.A1(_0987_),
    .A2(_2741_),
    .B1(_2742_),
    .B2(_0976_),
    .C1(_2819_),
    .X(_2820_));
 sky130_fd_sc_hd__nand2_1 _7470_ (.A(_1014_),
    .B(_2749_),
    .Y(_2821_));
 sky130_fd_sc_hd__o221a_1 _7471_ (.A1(_2131_),
    .A2(_2680_),
    .B1(_2682_),
    .B2(_2820_),
    .C1(_2821_),
    .X(_2822_));
 sky130_fd_sc_hd__a2bb2o_1 _7472_ (.A1_N(_2817_),
    .A2_N(_2822_),
    .B1(_0986_),
    .B2(_2686_),
    .X(net538));
 sky130_fd_sc_hd__a22o_1 _7473_ (.A1(_1025_),
    .A2(_2671_),
    .B1(_1058_),
    .B2(_0588_),
    .X(_2823_));
 sky130_fd_sc_hd__nor2_1 _7474_ (.A(_2668_),
    .B(_0993_),
    .Y(_2824_));
 sky130_fd_sc_hd__a221o_1 _7475_ (.A1(_0973_),
    .A2(_2666_),
    .B1(_2823_),
    .B2(_2710_),
    .C1(_2824_),
    .X(_2825_));
 sky130_fd_sc_hd__and2_1 _7476_ (.A(_2145_),
    .B(_2721_),
    .X(_2826_));
 sky130_fd_sc_hd__a221o_1 _7477_ (.A1(_1019_),
    .A2(_2749_),
    .B1(_2825_),
    .B2(_2692_),
    .C1(_2826_),
    .X(_2827_));
 sky130_fd_sc_hd__mux2_1 _7478_ (.A0(_2827_),
    .A1(_1017_),
    .S(_2686_),
    .X(_2828_));
 sky130_fd_sc_hd__buf_1 _7479_ (.A(_2828_),
    .X(net539));
 sky130_fd_sc_hd__a22o_1 _7480_ (.A1(_2526_),
    .A2(_2671_),
    .B1(_1037_),
    .B2(_2725_),
    .X(_2829_));
 sky130_fd_sc_hd__a22o_1 _7481_ (.A1(_0990_),
    .A2(_2666_),
    .B1(_1023_),
    .B2(_2723_),
    .X(_2830_));
 sky130_fd_sc_hd__a21o_1 _7482_ (.A1(_2710_),
    .A2(_2829_),
    .B1(_2830_),
    .X(_2831_));
 sky130_fd_sc_hd__nor2_1 _7483_ (.A(_2680_),
    .B(_2151_),
    .Y(_2832_));
 sky130_fd_sc_hd__a221o_1 _7484_ (.A1(_1064_),
    .A2(_2749_),
    .B1(_2831_),
    .B2(_2692_),
    .C1(_2832_),
    .X(_2833_));
 sky130_fd_sc_hd__mux2_1 _7485_ (.A0(_2833_),
    .A1(_1050_),
    .S(_2686_),
    .X(_2834_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _7486_ (.A(_2834_),
    .X(net540));
 sky130_fd_sc_hd__a221o_1 _7487_ (.A1(_1068_),
    .A2(_2768_),
    .B1(_1098_),
    .B2(_2725_),
    .C1(_2670_),
    .X(_2835_));
 sky130_fd_sc_hd__nand2_1 _7488_ (.A(_1054_),
    .B(_2724_),
    .Y(_2836_));
 sky130_fd_sc_hd__o21a_1 _7489_ (.A1(_2741_),
    .A2(_1021_),
    .B1(_2692_),
    .X(_2837_));
 sky130_fd_sc_hd__a22o_1 _7490_ (.A1(_1077_),
    .A2(_2678_),
    .B1(_2161_),
    .B2(_2721_),
    .X(_2838_));
 sky130_fd_sc_hd__a31o_1 _7491_ (.A1(_2835_),
    .A2(_2836_),
    .A3(_2837_),
    .B1(_2838_),
    .X(_2839_));
 sky130_fd_sc_hd__mux2_1 _7492_ (.A0(_2839_),
    .A1(_1067_),
    .S(_2686_),
    .X(_2840_));
 sky130_fd_sc_hd__clkbuf_2 _7493_ (.A(_2840_),
    .X(net541));
 sky130_fd_sc_hd__o21ai_2 _7494_ (.A1(_4094_),
    .A2(_1106_),
    .B1(_0168_),
    .Y(_2841_));
 sky130_fd_sc_hd__a21o_1 _7495_ (.A1(_1052_),
    .A2(_0613_),
    .B1(_4184_),
    .X(_2842_));
 sky130_fd_sc_hd__a22o_1 _7496_ (.A1(_1099_),
    .A2(_2768_),
    .B1(_2842_),
    .B2(_0288_),
    .X(_2843_));
 sky130_fd_sc_hd__nand2_1 _7497_ (.A(_2843_),
    .B(_2744_),
    .Y(_2844_));
 sky130_fd_sc_hd__nand2_1 _7498_ (.A(_1128_),
    .B(_0589_),
    .Y(_2845_));
 sky130_fd_sc_hd__a22o_1 _7499_ (.A1(_1101_),
    .A2(_2670_),
    .B1(_2844_),
    .B2(_2845_),
    .X(_2846_));
 sky130_fd_sc_hd__a2bb2o_1 _7500_ (.A1_N(_1081_),
    .A2_N(_2679_),
    .B1(_2733_),
    .B2(_2841_),
    .X(_2847_));
 sky130_fd_sc_hd__a221o_1 _7501_ (.A1(_1085_),
    .A2(_2722_),
    .B1(_2846_),
    .B2(_2693_),
    .C1(_2847_),
    .X(_2848_));
 sky130_fd_sc_hd__o221ai_4 _7502_ (.A1(_2736_),
    .A2(_2841_),
    .B1(_0138_),
    .B2(_1162_),
    .C1(_2848_),
    .Y(net542));
 sky130_fd_sc_hd__o21ai_1 _7503_ (.A1(_2675_),
    .A2(_1111_),
    .B1(_2711_),
    .Y(_2849_));
 sky130_fd_sc_hd__o221a_1 _7504_ (.A1(_1071_),
    .A2(_2667_),
    .B1(_2742_),
    .B2(_1091_),
    .C1(_2849_),
    .X(_2850_));
 sky130_fd_sc_hd__or2_1 _7505_ (.A(_2682_),
    .B(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__o21a_1 _7506_ (.A1(_2700_),
    .A2(_1083_),
    .B1(_2696_),
    .X(_2852_));
 sky130_fd_sc_hd__nor2_1 _7507_ (.A(_2684_),
    .B(_1161_),
    .Y(_2853_));
 sky130_fd_sc_hd__a221o_1 _7508_ (.A1(_1167_),
    .A2(_2720_),
    .B1(_2851_),
    .B2(_2852_),
    .C1(_2853_),
    .X(net543));
 sky130_fd_sc_hd__nand2_1 _7509_ (.A(_1145_),
    .B(_4239_),
    .Y(_2854_));
 sky130_fd_sc_hd__nand2_1 _7510_ (.A(_4241_),
    .B(_4094_),
    .Y(_2855_));
 sky130_fd_sc_hd__nand2_2 _7511_ (.A(_2855_),
    .B(_0342_),
    .Y(_2856_));
 sky130_fd_sc_hd__inv_2 _7512_ (.A(_2856_),
    .Y(_2857_));
 sky130_fd_sc_hd__o22a_1 _7513_ (.A1(_1090_),
    .A2(_2741_),
    .B1(_2742_),
    .B2(_1137_),
    .X(_2858_));
 sky130_fd_sc_hd__nand2_1 _7514_ (.A(_1174_),
    .B(_2768_),
    .Y(_2859_));
 sky130_fd_sc_hd__a31o_1 _7515_ (.A1(_2859_),
    .A2(_0056_),
    .A3(_2668_),
    .B1(_2745_),
    .X(_2860_));
 sky130_fd_sc_hd__o21ai_1 _7516_ (.A1(_1007_),
    .A2(_1123_),
    .B1(_2860_),
    .Y(_2861_));
 sky130_fd_sc_hd__a22o_1 _7517_ (.A1(_2854_),
    .A2(_2857_),
    .B1(_2858_),
    .B2(_2861_),
    .X(_2862_));
 sky130_fd_sc_hd__o21ai_1 _7518_ (.A1(_4094_),
    .A2(_1158_),
    .B1(_0168_),
    .Y(_2863_));
 sky130_fd_sc_hd__o2bb2a_1 _7519_ (.A1_N(_2733_),
    .A2_N(_2863_),
    .B1(_1144_),
    .B2(_2700_),
    .X(_2864_));
 sky130_fd_sc_hd__nor2_1 _7520_ (.A(_2736_),
    .B(_2863_),
    .Y(_2865_));
 sky130_fd_sc_hd__a221o_2 _7521_ (.A1(_1165_),
    .A2(_2720_),
    .B1(_2862_),
    .B2(_2864_),
    .C1(_2865_),
    .X(net544));
 sky130_fd_sc_hd__o21a_1 _7522_ (.A1(_4094_),
    .A2(_1155_),
    .B1(_0168_),
    .X(_2866_));
 sky130_fd_sc_hd__a22o_1 _7523_ (.A1(_1117_),
    .A2(_2671_),
    .B1(_1183_),
    .B2(_0588_),
    .X(_2867_));
 sky130_fd_sc_hd__and2_1 _7524_ (.A(_0995_),
    .B(_2666_),
    .X(_2868_));
 sky130_fd_sc_hd__a221o_2 _7525_ (.A1(_1190_),
    .A2(_2724_),
    .B1(_2867_),
    .B2(_2710_),
    .C1(_2868_),
    .X(_2869_));
 sky130_fd_sc_hd__nor2_1 _7526_ (.A(_2679_),
    .B(_1142_),
    .Y(_2870_));
 sky130_fd_sc_hd__a221o_1 _7527_ (.A1(_2187_),
    .A2(_2722_),
    .B1(_2869_),
    .B2(_2692_),
    .C1(_2870_),
    .X(_2871_));
 sky130_fd_sc_hd__or2_1 _7528_ (.A(_2800_),
    .B(_2866_),
    .X(_2872_));
 sky130_fd_sc_hd__nor2_1 _7529_ (.A(_0138_),
    .B(_1171_),
    .Y(_2873_));
 sky130_fd_sc_hd__a221o_1 _7530_ (.A1(_4095_),
    .A2(_2866_),
    .B1(_2871_),
    .B2(_2872_),
    .C1(_2873_),
    .X(net545));
 sky130_fd_sc_hd__nand2_1 _7531_ (.A(_1206_),
    .B(_0588_),
    .Y(_2874_));
 sky130_fd_sc_hd__nor2_1 _7532_ (.A(_2672_),
    .B(_1180_),
    .Y(_2875_));
 sky130_fd_sc_hd__a21oi_1 _7533_ (.A1(_1197_),
    .A2(_4233_),
    .B1(_0287_),
    .Y(_2876_));
 sky130_fd_sc_hd__o21ai_1 _7534_ (.A1(_2875_),
    .A2(_2876_),
    .B1(_2744_),
    .Y(_2877_));
 sky130_fd_sc_hd__a2bb2o_2 _7535_ (.A1_N(_0997_),
    .A2_N(_2710_),
    .B1(_2874_),
    .B2(_2877_),
    .X(_2878_));
 sky130_fd_sc_hd__nand2_1 _7536_ (.A(_2857_),
    .B(_0572_),
    .Y(_2879_));
 sky130_fd_sc_hd__a22o_1 _7537_ (.A1(_0572_),
    .A2(_2189_),
    .B1(_2878_),
    .B2(_2879_),
    .X(_2880_));
 sky130_fd_sc_hd__a21o_1 _7538_ (.A1(_2878_),
    .A2(_2856_),
    .B1(_4239_),
    .X(_2881_));
 sky130_fd_sc_hd__a221o_1 _7539_ (.A1(_2189_),
    .A2(_2749_),
    .B1(_2880_),
    .B2(_2881_),
    .C1(_2686_),
    .X(_2882_));
 sky130_fd_sc_hd__o21ai_2 _7540_ (.A1(_1170_),
    .A2(_2698_),
    .B1(_2882_),
    .Y(net547));
 sky130_fd_sc_hd__a22o_1 _7541_ (.A1(_2193_),
    .A2(_2768_),
    .B1(_1225_),
    .B2(_2725_),
    .X(_2883_));
 sky130_fd_sc_hd__nor2_1 _7542_ (.A(_2741_),
    .B(_1196_),
    .Y(_2884_));
 sky130_fd_sc_hd__a221o_2 _7543_ (.A1(_1004_),
    .A2(_2724_),
    .B1(_2883_),
    .B2(_2711_),
    .C1(_2884_),
    .X(_2885_));
 sky130_fd_sc_hd__and2_1 _7544_ (.A(_1215_),
    .B(_2749_),
    .X(_2886_));
 sky130_fd_sc_hd__a221o_1 _7545_ (.A1(_2202_),
    .A2(_2722_),
    .B1(_2885_),
    .B2(_2700_),
    .C1(_2886_),
    .X(_2887_));
 sky130_fd_sc_hd__o21ai_1 _7546_ (.A1(_2738_),
    .A2(_1232_),
    .B1(_2757_),
    .Y(_2888_));
 sky130_fd_sc_hd__nand2_1 _7547_ (.A(_2888_),
    .B(_2734_),
    .Y(_2889_));
 sky130_fd_sc_hd__a2bb2o_1 _7548_ (.A1_N(_2731_),
    .A2_N(_2888_),
    .B1(_2719_),
    .B2(_2201_),
    .X(_2890_));
 sky130_fd_sc_hd__a21o_1 _7549_ (.A1(_2887_),
    .A2(_2889_),
    .B1(_2890_),
    .X(net548));
 sky130_fd_sc_hd__a22o_1 _7550_ (.A1(_1257_),
    .A2(_2671_),
    .B1(_1240_),
    .B2(_0588_),
    .X(_2891_));
 sky130_fd_sc_hd__and2_1 _7551_ (.A(_1002_),
    .B(_2666_),
    .X(_2892_));
 sky130_fd_sc_hd__a221o_2 _7552_ (.A1(_1247_),
    .A2(_2724_),
    .B1(_2891_),
    .B2(_2710_),
    .C1(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__mux2_1 _7553_ (.A0(_2893_),
    .A1(_1277_),
    .S(_2682_),
    .X(_2894_));
 sky130_fd_sc_hd__o21ai_1 _7554_ (.A1(_2738_),
    .A2(_1256_),
    .B1(_2757_),
    .Y(_2895_));
 sky130_fd_sc_hd__nand2_1 _7555_ (.A(_2895_),
    .B(_2734_),
    .Y(_2896_));
 sky130_fd_sc_hd__nor2_1 _7556_ (.A(_2736_),
    .B(_2895_),
    .Y(_2897_));
 sky130_fd_sc_hd__a221o_1 _7557_ (.A1(_2221_),
    .A2(_2720_),
    .B1(_2894_),
    .B2(_2896_),
    .C1(_2897_),
    .X(net549));
 sky130_fd_sc_hd__nand2_1 _7558_ (.A(_2224_),
    .B(_4239_),
    .Y(_2898_));
 sky130_fd_sc_hd__o22a_1 _7559_ (.A1(_1246_),
    .A2(_2741_),
    .B1(_2742_),
    .B2(_1272_),
    .X(_2899_));
 sky130_fd_sc_hd__nand2_1 _7560_ (.A(_1294_),
    .B(_2768_),
    .Y(_2900_));
 sky130_fd_sc_hd__a31o_1 _7561_ (.A1(_2900_),
    .A2(_0056_),
    .A3(_2668_),
    .B1(_2745_),
    .X(_2901_));
 sky130_fd_sc_hd__o21ai_2 _7562_ (.A1(_1007_),
    .A2(_1261_),
    .B1(_2901_),
    .Y(_2902_));
 sky130_fd_sc_hd__a22o_1 _7563_ (.A1(_2857_),
    .A2(_2898_),
    .B1(_2899_),
    .B2(_2902_),
    .X(_2903_));
 sky130_fd_sc_hd__o21ai_1 _7564_ (.A1(_4094_),
    .A2(_1282_),
    .B1(_0168_),
    .Y(_2904_));
 sky130_fd_sc_hd__o2bb2a_1 _7565_ (.A1_N(_2733_),
    .A2_N(_2904_),
    .B1(_1304_),
    .B2(_2700_),
    .X(_2905_));
 sky130_fd_sc_hd__nor2_1 _7566_ (.A(_2736_),
    .B(_2904_),
    .Y(_2906_));
 sky130_fd_sc_hd__a221o_2 _7567_ (.A1(_1285_),
    .A2(_2720_),
    .B1(_2903_),
    .B2(_2905_),
    .C1(_2906_),
    .X(net550));
 sky130_fd_sc_hd__nor2_1 _7568_ (.A(_2667_),
    .B(_1313_),
    .Y(_2907_));
 sky130_fd_sc_hd__a221o_1 _7569_ (.A1(_1260_),
    .A2(_2676_),
    .B1(_2231_),
    .B2(_2724_),
    .C1(_2907_),
    .X(_2908_));
 sky130_fd_sc_hd__nor2_1 _7570_ (.A(_2680_),
    .B(_1308_),
    .Y(_2909_));
 sky130_fd_sc_hd__a221o_1 _7571_ (.A1(_1299_),
    .A2(_2678_),
    .B1(_2908_),
    .B2(_2692_),
    .C1(_2909_),
    .X(_2910_));
 sky130_fd_sc_hd__mux2_1 _7572_ (.A0(_2910_),
    .A1(_1284_),
    .S(_2686_),
    .X(_2911_));
 sky130_fd_sc_hd__buf_1 _7573_ (.A(_2911_),
    .X(net551));
 sky130_fd_sc_hd__a22o_1 _7574_ (.A1(_2566_),
    .A2(_2671_),
    .B1(_1324_),
    .B2(_2725_),
    .X(_2912_));
 sky130_fd_sc_hd__nor2_1 _7575_ (.A(_2668_),
    .B(_2244_),
    .Y(_2913_));
 sky130_fd_sc_hd__a221o_2 _7576_ (.A1(_1335_),
    .A2(_2666_),
    .B1(_2912_),
    .B2(_2710_),
    .C1(_2913_),
    .X(_2914_));
 sky130_fd_sc_hd__nor2_1 _7577_ (.A(_2680_),
    .B(_2250_),
    .Y(_2915_));
 sky130_fd_sc_hd__a221o_1 _7578_ (.A1(_1301_),
    .A2(_2749_),
    .B1(_2914_),
    .B2(_2692_),
    .C1(_2915_),
    .X(_2916_));
 sky130_fd_sc_hd__o21ai_1 _7579_ (.A1(_2738_),
    .A2(_1333_),
    .B1(_2757_),
    .Y(_2917_));
 sky130_fd_sc_hd__nand2_1 _7580_ (.A(_2917_),
    .B(_2734_),
    .Y(_2918_));
 sky130_fd_sc_hd__nor2_1 _7581_ (.A(_2736_),
    .B(_2917_),
    .Y(_2919_));
 sky130_fd_sc_hd__a221o_2 _7582_ (.A1(_2255_),
    .A2(_2720_),
    .B1(_2916_),
    .B2(_2918_),
    .C1(_2919_),
    .X(net552));
 sky130_fd_sc_hd__a221o_1 _7583_ (.A1(_1373_),
    .A2(_2768_),
    .B1(_1412_),
    .B2(_0589_),
    .C1(_2670_),
    .X(_2920_));
 sky130_fd_sc_hd__nand2_1 _7584_ (.A(_1352_),
    .B(_2724_),
    .Y(_2921_));
 sky130_fd_sc_hd__o21a_1 _7585_ (.A1(_2741_),
    .A2(_1347_),
    .B1(_2692_),
    .X(_2922_));
 sky130_fd_sc_hd__a22o_1 _7586_ (.A1(_1390_),
    .A2(_2678_),
    .B1(_2264_),
    .B2(_2722_),
    .X(_2923_));
 sky130_fd_sc_hd__a31o_2 _7587_ (.A1(_2920_),
    .A2(_2921_),
    .A3(_2922_),
    .B1(_2923_),
    .X(_2924_));
 sky130_fd_sc_hd__o21ai_1 _7588_ (.A1(_2738_),
    .A2(_1361_),
    .B1(_2757_),
    .Y(_2925_));
 sky130_fd_sc_hd__nand2_1 _7589_ (.A(_2925_),
    .B(_2734_),
    .Y(_2926_));
 sky130_fd_sc_hd__nor2_1 _7590_ (.A(_2736_),
    .B(_2925_),
    .Y(_2927_));
 sky130_fd_sc_hd__a221o_1 _7591_ (.A1(_2270_),
    .A2(_2720_),
    .B1(_2924_),
    .B2(_2926_),
    .C1(_2927_),
    .X(net553));
 sky130_fd_sc_hd__nand2_1 _7592_ (.A(_1384_),
    .B(_2725_),
    .Y(_2928_));
 sky130_fd_sc_hd__o21a_1 _7593_ (.A1(_2672_),
    .A2(_1382_),
    .B1(_2710_),
    .X(_2929_));
 sky130_fd_sc_hd__o21ai_1 _7594_ (.A1(_2741_),
    .A2(_1345_),
    .B1(_2692_),
    .Y(_2930_));
 sky130_fd_sc_hd__a221o_2 _7595_ (.A1(_2928_),
    .A2(_2929_),
    .B1(_1371_),
    .B2(_2724_),
    .C1(_2930_),
    .X(_2931_));
 sky130_fd_sc_hd__o221ai_4 _7596_ (.A1(_2266_),
    .A2(_2679_),
    .B1(_2279_),
    .B2(_2680_),
    .C1(_2931_),
    .Y(_2932_));
 sky130_fd_sc_hd__o21ai_1 _7597_ (.A1(_2738_),
    .A2(_1393_),
    .B1(_2757_),
    .Y(_2933_));
 sky130_fd_sc_hd__nand2_1 _7598_ (.A(_2933_),
    .B(_2734_),
    .Y(_2934_));
 sky130_fd_sc_hd__nor2_1 _7599_ (.A(_2731_),
    .B(_2933_),
    .Y(_2935_));
 sky130_fd_sc_hd__a221o_1 _7600_ (.A1(_1396_),
    .A2(_2720_),
    .B1(_2932_),
    .B2(_2934_),
    .C1(_2935_),
    .X(net554));
 sky130_fd_sc_hd__o21a_1 _7601_ (.A1(_4094_),
    .A2(_1395_),
    .B1(_0168_),
    .X(_2936_));
 sky130_fd_sc_hd__a221o_1 _7602_ (.A1(_1436_),
    .A2(_2768_),
    .B1(_1479_),
    .B2(_2725_),
    .C1(_2669_),
    .X(_2937_));
 sky130_fd_sc_hd__o21a_1 _7603_ (.A1(_2710_),
    .A2(_1367_),
    .B1(_2691_),
    .X(_2938_));
 sky130_fd_sc_hd__nor2_1 _7604_ (.A(_2680_),
    .B(_2293_),
    .Y(_2939_));
 sky130_fd_sc_hd__a221o_1 _7605_ (.A1(_1435_),
    .A2(_2749_),
    .B1(_2937_),
    .B2(_2938_),
    .C1(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__or2_1 _7606_ (.A(_2800_),
    .B(_2936_),
    .X(_2941_));
 sky130_fd_sc_hd__nor2_1 _7607_ (.A(_0138_),
    .B(_1406_),
    .Y(_2942_));
 sky130_fd_sc_hd__a221o_1 _7608_ (.A1(_4095_),
    .A2(_2936_),
    .B1(_2940_),
    .B2(_2941_),
    .C1(_2942_),
    .X(net555));
 sky130_fd_sc_hd__o21ai_2 _7609_ (.A1(_2738_),
    .A2(_1404_),
    .B1(_0168_),
    .Y(_2943_));
 sky130_fd_sc_hd__nand2_1 _7610_ (.A(_1433_),
    .B(_2720_),
    .Y(_2944_));
 sky130_fd_sc_hd__nand2_1 _7611_ (.A(_1469_),
    .B(_2768_),
    .Y(_2945_));
 sky130_fd_sc_hd__a31o_1 _7612_ (.A1(_2945_),
    .A2(_0056_),
    .A3(_2742_),
    .B1(_2745_),
    .X(_2946_));
 sky130_fd_sc_hd__o21ai_1 _7613_ (.A1(_1007_),
    .A2(_1446_),
    .B1(_2946_),
    .Y(_2947_));
 sky130_fd_sc_hd__o221ai_4 _7614_ (.A1(_1418_),
    .A2(_2741_),
    .B1(_2742_),
    .B2(_1457_),
    .C1(_2947_),
    .Y(_2948_));
 sky130_fd_sc_hd__a22o_1 _7615_ (.A1(_2295_),
    .A2(_2749_),
    .B1(_2305_),
    .B2(_2722_),
    .X(_2949_));
 sky130_fd_sc_hd__a221o_1 _7616_ (.A1(_2733_),
    .A2(_2943_),
    .B1(_2948_),
    .B2(_2700_),
    .C1(_2949_),
    .X(_2950_));
 sky130_fd_sc_hd__o211ai_4 _7617_ (.A1(_2736_),
    .A2(_2943_),
    .B1(_2944_),
    .C1(_2950_),
    .Y(net556));
 sky130_fd_sc_hd__o21ai_2 _7618_ (.A1(_2738_),
    .A2(_1428_),
    .B1(_0168_),
    .Y(_2951_));
 sky130_fd_sc_hd__nand2_1 _7619_ (.A(_1466_),
    .B(_2720_),
    .Y(_2952_));
 sky130_fd_sc_hd__nand2_1 _7620_ (.A(_1502_),
    .B(_2768_),
    .Y(_2953_));
 sky130_fd_sc_hd__a31o_1 _7621_ (.A1(_2953_),
    .A2(_0056_),
    .A3(_2668_),
    .B1(_2745_),
    .X(_2954_));
 sky130_fd_sc_hd__nand2_1 _7622_ (.A(_1476_),
    .B(_0589_),
    .Y(_2955_));
 sky130_fd_sc_hd__nor2_1 _7623_ (.A(_2742_),
    .B(_1488_),
    .Y(_2956_));
 sky130_fd_sc_hd__a221o_2 _7624_ (.A1(_1506_),
    .A2(_2666_),
    .B1(_2954_),
    .B2(_2955_),
    .C1(_2956_),
    .X(_2957_));
 sky130_fd_sc_hd__a22o_1 _7625_ (.A1(_2307_),
    .A2(_2749_),
    .B1(_2951_),
    .B2(_2733_),
    .X(_2958_));
 sky130_fd_sc_hd__a221o_1 _7626_ (.A1(_2316_),
    .A2(_2722_),
    .B1(_2957_),
    .B2(_2700_),
    .C1(_2958_),
    .X(_2959_));
 sky130_fd_sc_hd__o211ai_4 _7627_ (.A1(_2736_),
    .A2(_2951_),
    .B1(_2952_),
    .C1(_2959_),
    .Y(net558));
 sky130_fd_sc_hd__o21ai_2 _7628_ (.A1(_2738_),
    .A2(_1462_),
    .B1(_2757_),
    .Y(_2960_));
 sky130_fd_sc_hd__nand2_1 _7629_ (.A(_1498_),
    .B(_0589_),
    .Y(_2961_));
 sky130_fd_sc_hd__nand2_1 _7630_ (.A(_1474_),
    .B(_2671_),
    .Y(_2962_));
 sky130_fd_sc_hd__a31o_1 _7631_ (.A1(_2962_),
    .A2(_0056_),
    .A3(_2668_),
    .B1(_2745_),
    .X(_2963_));
 sky130_fd_sc_hd__nor2_1 _7632_ (.A(_2742_),
    .B(_1545_),
    .Y(_2964_));
 sky130_fd_sc_hd__a221o_2 _7633_ (.A1(_1531_),
    .A2(_2666_),
    .B1(_2961_),
    .B2(_2963_),
    .C1(_2964_),
    .X(_2965_));
 sky130_fd_sc_hd__a2bb2o_1 _7634_ (.A1_N(_1535_),
    .A2_N(_2679_),
    .B1(_2722_),
    .B2(_2326_),
    .X(_2966_));
 sky130_fd_sc_hd__a221o_1 _7635_ (.A1(_2733_),
    .A2(_2960_),
    .B1(_2965_),
    .B2(_2693_),
    .C1(_2966_),
    .X(_2967_));
 sky130_fd_sc_hd__o221ai_4 _7636_ (.A1(_2736_),
    .A2(_2960_),
    .B1(_0138_),
    .B2(_1561_),
    .C1(_2967_),
    .Y(net559));
 sky130_fd_sc_hd__or2_1 _7637_ (.A(_2742_),
    .B(_1522_),
    .X(_2968_));
 sky130_fd_sc_hd__nand2_1 _7638_ (.A(_1528_),
    .B(_2725_),
    .Y(_2969_));
 sky130_fd_sc_hd__nand2_1 _7639_ (.A(_1548_),
    .B(_2768_),
    .Y(_2970_));
 sky130_fd_sc_hd__nand3_1 _7640_ (.A(_2969_),
    .B(_2711_),
    .C(_2970_),
    .Y(_2971_));
 sky130_fd_sc_hd__o21a_1 _7641_ (.A1(_2741_),
    .A2(_1518_),
    .B1(_2692_),
    .X(_2972_));
 sky130_fd_sc_hd__a22o_1 _7642_ (.A1(_1564_),
    .A2(_2678_),
    .B1(_2337_),
    .B2(_2722_),
    .X(_2973_));
 sky130_fd_sc_hd__a31o_2 _7643_ (.A1(_2968_),
    .A2(_2971_),
    .A3(_2972_),
    .B1(_2973_),
    .X(_2974_));
 sky130_fd_sc_hd__o21ai_1 _7644_ (.A1(_2738_),
    .A2(_1539_),
    .B1(_2757_),
    .Y(_2975_));
 sky130_fd_sc_hd__nand2_1 _7645_ (.A(_2975_),
    .B(_2734_),
    .Y(_2976_));
 sky130_fd_sc_hd__nor2_1 _7646_ (.A(_2731_),
    .B(_2975_),
    .Y(_2977_));
 sky130_fd_sc_hd__a221o_1 _7647_ (.A1(_2347_),
    .A2(_2720_),
    .B1(_2974_),
    .B2(_2976_),
    .C1(_2977_),
    .X(net560));
 sky130_fd_sc_hd__or2_1 _7648_ (.A(_2742_),
    .B(_1547_),
    .X(_2978_));
 sky130_fd_sc_hd__o21ai_1 _7649_ (.A1(_2672_),
    .A2(_1526_),
    .B1(_2710_),
    .Y(_2979_));
 sky130_fd_sc_hd__nor2_1 _7650_ (.A(_1007_),
    .B(_1553_),
    .Y(_2980_));
 sky130_fd_sc_hd__or2_1 _7651_ (.A(_2979_),
    .B(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__o21a_1 _7652_ (.A1(_2741_),
    .A2(_1515_),
    .B1(_2692_),
    .X(_2982_));
 sky130_fd_sc_hd__a22o_1 _7653_ (.A1(_1588_),
    .A2(_2678_),
    .B1(_1609_),
    .B2(_2722_),
    .X(_2983_));
 sky130_fd_sc_hd__a31o_2 _7654_ (.A1(_2978_),
    .A2(_2981_),
    .A3(_2982_),
    .B1(_2983_),
    .X(_2984_));
 sky130_fd_sc_hd__o21ai_1 _7655_ (.A1(_2738_),
    .A2(_1591_),
    .B1(_2757_),
    .Y(_2985_));
 sky130_fd_sc_hd__nand2_1 _7656_ (.A(_2985_),
    .B(_2734_),
    .Y(_2986_));
 sky130_fd_sc_hd__nor2_1 _7657_ (.A(_2731_),
    .B(_2985_),
    .Y(_2987_));
 sky130_fd_sc_hd__a221o_1 _7658_ (.A1(_0209_),
    .A2(_1595_),
    .B1(_2984_),
    .B2(_2986_),
    .C1(_2987_),
    .X(net561));
 sky130_fd_sc_hd__a22o_1 _7659_ (.A1(_2340_),
    .A2(_2768_),
    .B1(_1583_),
    .B2(_2725_),
    .X(_2988_));
 sky130_fd_sc_hd__and2_1 _7660_ (.A(_1541_),
    .B(_2666_),
    .X(_2989_));
 sky130_fd_sc_hd__a221o_1 _7661_ (.A1(_1574_),
    .A2(_2724_),
    .B1(_2988_),
    .B2(_2711_),
    .C1(_2989_),
    .X(_2990_));
 sky130_fd_sc_hd__a22o_1 _7662_ (.A1(_1605_),
    .A2(_2749_),
    .B1(_2357_),
    .B2(_2722_),
    .X(_2991_));
 sky130_fd_sc_hd__a21o_1 _7663_ (.A1(_2990_),
    .A2(_2693_),
    .B1(_2991_),
    .X(_2992_));
 sky130_fd_sc_hd__o21ai_1 _7664_ (.A1(_2731_),
    .A2(_1594_),
    .B1(_1757_),
    .Y(_2993_));
 sky130_fd_sc_hd__nand2_1 _7665_ (.A(_2993_),
    .B(_2734_),
    .Y(_2994_));
 sky130_fd_sc_hd__o22ai_1 _7666_ (.A1(_2736_),
    .A2(_2993_),
    .B1(_2685_),
    .B2(_2349_),
    .Y(_2995_));
 sky130_fd_sc_hd__a21o_1 _7667_ (.A1(_2992_),
    .A2(_2994_),
    .B1(_2995_),
    .X(net562));
 sky130_fd_sc_hd__nand2_1 _7668_ (.A(_2351_),
    .B(_2768_),
    .Y(_2996_));
 sky130_fd_sc_hd__a31o_1 _7669_ (.A1(_2996_),
    .A2(_0056_),
    .A3(_2742_),
    .B1(_2745_),
    .X(_2997_));
 sky130_fd_sc_hd__o21ai_1 _7670_ (.A1(_1007_),
    .A2(_1622_),
    .B1(_2997_),
    .Y(_2998_));
 sky130_fd_sc_hd__o221ai_4 _7671_ (.A1(_1570_),
    .A2(_2741_),
    .B1(_2742_),
    .B2(_1619_),
    .C1(_2998_),
    .Y(_2999_));
 sky130_fd_sc_hd__nand2_1 _7672_ (.A(_2999_),
    .B(_2693_),
    .Y(_3000_));
 sky130_fd_sc_hd__or2_1 _7673_ (.A(_2680_),
    .B(_1611_),
    .X(_3001_));
 sky130_fd_sc_hd__o21a_1 _7674_ (.A1(_2738_),
    .A2(_1636_),
    .B1(_0168_),
    .X(_3002_));
 sky130_fd_sc_hd__o22a_1 _7675_ (.A1(_1601_),
    .A2(_2679_),
    .B1(_2800_),
    .B2(_3002_),
    .X(_3003_));
 sky130_fd_sc_hd__a22o_1 _7676_ (.A1(_4095_),
    .A2(_3002_),
    .B1(_2369_),
    .B2(_2719_),
    .X(_3004_));
 sky130_fd_sc_hd__a31o_1 _7677_ (.A1(_3000_),
    .A2(_3001_),
    .A3(_3003_),
    .B1(_3004_),
    .X(net563));
 sky130_fd_sc_hd__nor2_1 _7678_ (.A(_2675_),
    .B(_1621_),
    .Y(_3005_));
 sky130_fd_sc_hd__o221a_1 _7679_ (.A1(_1614_),
    .A2(_2667_),
    .B1(_2669_),
    .B2(_3005_),
    .C1(_2691_),
    .X(_3006_));
 sky130_fd_sc_hd__nand2_1 _7680_ (.A(_1690_),
    .B(_2724_),
    .Y(_3007_));
 sky130_fd_sc_hd__nor2_1 _7681_ (.A(_2679_),
    .B(_1678_),
    .Y(_3008_));
 sky130_fd_sc_hd__a221o_1 _7682_ (.A1(_1701_),
    .A2(_2722_),
    .B1(_3006_),
    .B2(_3007_),
    .C1(_3008_),
    .X(_3009_));
 sky130_fd_sc_hd__and3_1 _7683_ (.A(_1640_),
    .B(_4095_),
    .C(_2757_),
    .X(_3010_));
 sky130_fd_sc_hd__a221o_1 _7684_ (.A1(_1643_),
    .A2(_2720_),
    .B1(_3009_),
    .B2(_2697_),
    .C1(_3010_),
    .X(net564));
 sky130_fd_sc_hd__a2bb2o_1 _7685_ (.A1_N(_2673_),
    .A2_N(_1665_),
    .B1(_2371_),
    .B2(_2671_),
    .X(_3011_));
 sky130_fd_sc_hd__nor2_1 _7686_ (.A(_2667_),
    .B(_1689_),
    .Y(_3012_));
 sky130_fd_sc_hd__a221o_1 _7687_ (.A1(_1654_),
    .A2(_2724_),
    .B1(_3011_),
    .B2(_2711_),
    .C1(_3012_),
    .X(_3013_));
 sky130_fd_sc_hd__a2bb2o_1 _7688_ (.A1_N(_2680_),
    .A2_N(_1676_),
    .B1(_1673_),
    .B2(_2678_),
    .X(_3014_));
 sky130_fd_sc_hd__a21o_1 _7689_ (.A1(_3013_),
    .A2(_2700_),
    .B1(_3014_),
    .X(_3015_));
 sky130_fd_sc_hd__o21ai_1 _7690_ (.A1(_2738_),
    .A2(_1638_),
    .B1(_2757_),
    .Y(_3016_));
 sky130_fd_sc_hd__nand2_1 _7691_ (.A(_3016_),
    .B(_2734_),
    .Y(_3017_));
 sky130_fd_sc_hd__nor2_1 _7692_ (.A(_2731_),
    .B(_3016_),
    .Y(_3018_));
 sky130_fd_sc_hd__a221o_1 _7693_ (.A1(_1687_),
    .A2(_2719_),
    .B1(_3015_),
    .B2(_3017_),
    .C1(_3018_),
    .X(net565));
 sky130_fd_sc_hd__nor2_1 _7694_ (.A(_2742_),
    .B(_1695_),
    .Y(_3019_));
 sky130_fd_sc_hd__a221o_1 _7695_ (.A1(_1646_),
    .A2(_2666_),
    .B1(_1717_),
    .B2(_2676_),
    .C1(_3019_),
    .X(_3020_));
 sky130_fd_sc_hd__nand2_1 _7696_ (.A(_1670_),
    .B(_2749_),
    .Y(_3021_));
 sky130_fd_sc_hd__o21ai_1 _7697_ (.A1(_2680_),
    .A2(_1707_),
    .B1(_3021_),
    .Y(_3022_));
 sky130_fd_sc_hd__a21o_1 _7698_ (.A1(_3020_),
    .A2(_2700_),
    .B1(_3022_),
    .X(_3023_));
 sky130_fd_sc_hd__o21ai_1 _7699_ (.A1(_2738_),
    .A2(_1681_),
    .B1(_2757_),
    .Y(_3024_));
 sky130_fd_sc_hd__nand2_1 _7700_ (.A(_3024_),
    .B(_2733_),
    .Y(_3025_));
 sky130_fd_sc_hd__nor2_1 _7701_ (.A(_2731_),
    .B(_3024_),
    .Y(_3026_));
 sky130_fd_sc_hd__a221o_1 _7702_ (.A1(_1715_),
    .A2(_2719_),
    .B1(_3023_),
    .B2(_3025_),
    .C1(_3026_),
    .X(net566));
 sky130_fd_sc_hd__a221o_1 _7703_ (.A1(_1692_),
    .A2(_2670_),
    .B1(_2382_),
    .B2(_2676_),
    .C1(_2682_),
    .X(_3027_));
 sky130_fd_sc_hd__o21ai_2 _7704_ (.A1(_1703_),
    .A2(_2693_),
    .B1(_3027_),
    .Y(_3028_));
 sky130_fd_sc_hd__nor2_1 _7705_ (.A(_2697_),
    .B(_1711_),
    .Y(_3029_));
 sky130_fd_sc_hd__a21oi_2 _7706_ (.A1(_3028_),
    .A2(_2698_),
    .B1(_3029_),
    .Y(net567));
 sky130_fd_sc_hd__or4_1 _7707_ (.A(_0083_),
    .B(_0771_),
    .C(_0096_),
    .D(_1733_),
    .X(_3030_));
 sky130_fd_sc_hd__a221o_1 _7708_ (.A1(_1735_),
    .A2(_2669_),
    .B1(_1738_),
    .B2(_2676_),
    .C1(_2681_),
    .X(_3031_));
 sky130_fd_sc_hd__o211a_1 _7709_ (.A1(_1733_),
    .A2(_2679_),
    .B1(_3030_),
    .C1(_3031_),
    .X(_3032_));
 sky130_fd_sc_hd__mux2_1 _7710_ (.A0(_3032_),
    .A1(_1742_),
    .S(_2686_),
    .X(_3033_));
 sky130_fd_sc_hd__buf_1 _7711_ (.A(_3033_),
    .X(net569));
 sky130_fd_sc_hd__o21ai_1 _7712_ (.A1(_2672_),
    .A2(_1749_),
    .B1(_2710_),
    .Y(_3034_));
 sky130_fd_sc_hd__a31o_1 _7713_ (.A1(_0588_),
    .A2(_0694_),
    .A3(_1750_),
    .B1(_3034_),
    .X(_3035_));
 sky130_fd_sc_hd__o21a_1 _7714_ (.A1(_1745_),
    .A2(_2711_),
    .B1(_3035_),
    .X(_3036_));
 sky130_fd_sc_hd__mux2_1 _7715_ (.A0(_3036_),
    .A1(_1753_),
    .S(_2681_),
    .X(_3037_));
 sky130_fd_sc_hd__mux2_1 _7716_ (.A0(_3037_),
    .A1(_1756_),
    .S(_2686_),
    .X(_3038_));
 sky130_fd_sc_hd__buf_1 _7717_ (.A(_3038_),
    .X(net570));
 sky130_fd_sc_hd__a221o_1 _7718_ (.A1(_2629_),
    .A2(_2670_),
    .B1(_1764_),
    .B2(_2676_),
    .C1(_2682_),
    .X(_3039_));
 sky130_fd_sc_hd__o21ai_1 _7719_ (.A1(_1779_),
    .A2(_2693_),
    .B1(_3039_),
    .Y(_3040_));
 sky130_fd_sc_hd__nor2_1 _7720_ (.A(_2697_),
    .B(_1762_),
    .Y(_3041_));
 sky130_fd_sc_hd__a21oi_2 _7721_ (.A1(_3040_),
    .A2(_2698_),
    .B1(_3041_),
    .Y(net571));
 sky130_fd_sc_hd__o22a_1 _7722_ (.A1(_2712_),
    .A2(_1793_),
    .B1(_2711_),
    .B2(_1769_),
    .X(_3042_));
 sky130_fd_sc_hd__nand2_1 _7723_ (.A(_3042_),
    .B(_2693_),
    .Y(_3043_));
 sky130_fd_sc_hd__o21ai_1 _7724_ (.A1(_1801_),
    .A2(_2693_),
    .B1(_3043_),
    .Y(_3044_));
 sky130_fd_sc_hd__nor2_1 _7725_ (.A(_2697_),
    .B(_1788_),
    .Y(_3045_));
 sky130_fd_sc_hd__a21oi_2 _7726_ (.A1(_3044_),
    .A2(_2698_),
    .B1(_3045_),
    .Y(net572));
 sky130_fd_sc_hd__a221o_1 _7727_ (.A1(_1807_),
    .A2(_2676_),
    .B1(_2404_),
    .B2(_2670_),
    .C1(_2682_),
    .X(_3046_));
 sky130_fd_sc_hd__o21ai_1 _7728_ (.A1(_1816_),
    .A2(_2693_),
    .B1(_3046_),
    .Y(_3047_));
 sky130_fd_sc_hd__nor2_1 _7729_ (.A(_2697_),
    .B(_1784_),
    .Y(_3048_));
 sky130_fd_sc_hd__a21oi_2 _7730_ (.A1(_3047_),
    .A2(_2698_),
    .B1(_3048_),
    .Y(net573));
 sky130_fd_sc_hd__a221o_1 _7731_ (.A1(_1822_),
    .A2(_2676_),
    .B1(_2641_),
    .B2(_2670_),
    .C1(_2682_),
    .X(_3049_));
 sky130_fd_sc_hd__o21ai_1 _7732_ (.A1(_1826_),
    .A2(_2693_),
    .B1(_3049_),
    .Y(_3050_));
 sky130_fd_sc_hd__nor2_1 _7733_ (.A(_2697_),
    .B(_1786_),
    .Y(_3051_));
 sky130_fd_sc_hd__a21oi_2 _7734_ (.A1(_3050_),
    .A2(_2698_),
    .B1(_3051_),
    .Y(net574));
 sky130_fd_sc_hd__a221o_1 _7735_ (.A1(_0229_),
    .A2(_2676_),
    .B1(_2411_),
    .B2(_2670_),
    .C1(_2682_),
    .X(_3052_));
 sky130_fd_sc_hd__o21ai_2 _7736_ (.A1(_0131_),
    .A2(_2693_),
    .B1(_3052_),
    .Y(_3053_));
 sky130_fd_sc_hd__nor2_1 _7737_ (.A(_2697_),
    .B(_0191_),
    .Y(_3054_));
 sky130_fd_sc_hd__a21oi_2 _7738_ (.A1(_3053_),
    .A2(_2698_),
    .B1(_3054_),
    .Y(net575));
 sky130_fd_sc_hd__a221o_1 _7739_ (.A1(_1836_),
    .A2(_2670_),
    .B1(_1839_),
    .B2(_2676_),
    .C1(_2681_),
    .X(_3055_));
 sky130_fd_sc_hd__o21a_1 _7740_ (.A1(_1842_),
    .A2(_2700_),
    .B1(_3055_),
    .X(_3056_));
 sky130_fd_sc_hd__mux2_1 _7741_ (.A0(_3056_),
    .A1(_1845_),
    .S(_2686_),
    .X(_3057_));
 sky130_fd_sc_hd__buf_1 _7742_ (.A(_3057_),
    .X(net576));
 sky130_fd_sc_hd__nand2_1 _7743_ (.A(_1855_),
    .B(_2670_),
    .Y(_3058_));
 sky130_fd_sc_hd__o21a_1 _7744_ (.A1(_2712_),
    .A2(_1852_),
    .B1(_2692_),
    .X(_3059_));
 sky130_fd_sc_hd__a2bb2o_1 _7745_ (.A1_N(_1850_),
    .A2_N(_2700_),
    .B1(_3058_),
    .B2(_3059_),
    .X(_3060_));
 sky130_fd_sc_hd__nor2_1 _7746_ (.A(_2697_),
    .B(_1848_),
    .Y(_3061_));
 sky130_fd_sc_hd__a21oi_2 _7747_ (.A1(_3060_),
    .A2(_2698_),
    .B1(_3061_),
    .Y(net577));
 sky130_fd_sc_hd__o22a_1 _7748_ (.A1(_2711_),
    .A2(_1864_),
    .B1(_2712_),
    .B2(_1866_),
    .X(_3062_));
 sky130_fd_sc_hd__mux2_1 _7749_ (.A0(_3062_),
    .A1(_1870_),
    .S(_2682_),
    .X(_3063_));
 sky130_fd_sc_hd__nor2_1 _7750_ (.A(_2697_),
    .B(_1873_),
    .Y(_3064_));
 sky130_fd_sc_hd__a21oi_2 _7751_ (.A1(_3063_),
    .A2(_2698_),
    .B1(_3064_),
    .Y(net578));
 sky130_fd_sc_hd__o2111ai_1 _7752_ (.A1(_2742_),
    .A2(_1878_),
    .B1(_2741_),
    .C1(_2674_),
    .D1(_1881_),
    .Y(_3065_));
 sky130_fd_sc_hd__nand2_1 _7753_ (.A(_1879_),
    .B(_2670_),
    .Y(_3066_));
 sky130_fd_sc_hd__nor2_1 _7754_ (.A(_2700_),
    .B(_1876_),
    .Y(_3067_));
 sky130_fd_sc_hd__a31o_1 _7755_ (.A1(_3065_),
    .A2(_2700_),
    .A3(_3066_),
    .B1(_3067_),
    .X(_3068_));
 sky130_fd_sc_hd__nor2_1 _7756_ (.A(_2697_),
    .B(_1885_),
    .Y(_3069_));
 sky130_fd_sc_hd__a21oi_2 _7757_ (.A1(_3068_),
    .A2(_2698_),
    .B1(_3069_),
    .Y(net580));
 sky130_fd_sc_hd__nor2_2 _7758_ (.A(_0138_),
    .B(_0469_),
    .Y(_3070_));
 sky130_fd_sc_hd__clkbuf_8 _7759_ (.A(_3070_),
    .X(_3071_));
 sky130_fd_sc_hd__clkbuf_8 _7760_ (.A(_3071_),
    .X(_3072_));
 sky130_fd_sc_hd__nand2_1 _7761_ (.A(_2439_),
    .B(_0104_),
    .Y(_3073_));
 sky130_fd_sc_hd__a32o_1 _7762_ (.A1(_3073_),
    .A2(_0651_),
    .A3(net293),
    .B1(net230),
    .B2(_2439_),
    .X(_3074_));
 sky130_fd_sc_hd__a221o_4 _7763_ (.A1(net233),
    .A2(_0194_),
    .B1(net330),
    .B2(_0766_),
    .C1(_3074_),
    .X(_3075_));
 sky130_fd_sc_hd__a22o_1 _7764_ (.A1(_0538_),
    .A2(net230),
    .B1(_1894_),
    .B2(net293),
    .X(_3076_));
 sky130_fd_sc_hd__a221o_4 _7765_ (.A1(net233),
    .A2(_0590_),
    .B1(net330),
    .B2(_0694_),
    .C1(_3076_),
    .X(_3077_));
 sky130_fd_sc_hd__nor2_2 _7766_ (.A(_4184_),
    .B(_0615_),
    .Y(_3078_));
 sky130_fd_sc_hd__nor3_2 _7767_ (.A(_1007_),
    .B(_0427_),
    .C(_3078_),
    .Y(_3079_));
 sky130_fd_sc_hd__clkbuf_8 _7768_ (.A(_3079_),
    .X(_3080_));
 sky130_fd_sc_hd__buf_12 _7769_ (.A(_4278_),
    .X(_3081_));
 sky130_fd_sc_hd__a22o_1 _7770_ (.A1(_4268_),
    .A2(net233),
    .B1(net330),
    .B2(_0613_),
    .X(_3082_));
 sky130_fd_sc_hd__a221o_4 _7771_ (.A1(net230),
    .A2(_3081_),
    .B1(_4273_),
    .B2(_1977_),
    .C1(_3082_),
    .X(_3083_));
 sky130_fd_sc_hd__clkbuf_8 _7772_ (.A(_3078_),
    .X(_3084_));
 sky130_fd_sc_hd__nor2_8 _7773_ (.A(_0083_),
    .B(_0451_),
    .Y(_3085_));
 sky130_fd_sc_hd__clkbuf_8 _7774_ (.A(_3085_),
    .X(_3086_));
 sky130_fd_sc_hd__a221o_1 _7775_ (.A1(_3077_),
    .A2(_3080_),
    .B1(_3083_),
    .B2(_3084_),
    .C1(_3086_),
    .X(_3087_));
 sky130_fd_sc_hd__inv_2 _7776_ (.A(_3085_),
    .Y(_3088_));
 sky130_fd_sc_hd__clkbuf_8 _7777_ (.A(_3088_),
    .X(_3089_));
 sky130_fd_sc_hd__nand2_1 _7778_ (.A(_0759_),
    .B(_0104_),
    .Y(_3090_));
 sky130_fd_sc_hd__a32o_1 _7779_ (.A1(_3090_),
    .A2(_0143_),
    .A3(net293),
    .B1(net230),
    .B2(_0759_),
    .X(_3091_));
 sky130_fd_sc_hd__a221o_4 _7780_ (.A1(net233),
    .A2(_0108_),
    .B1(net330),
    .B2(_0729_),
    .C1(_3091_),
    .X(_3092_));
 sky130_fd_sc_hd__o21ba_1 _7781_ (.A1(_3089_),
    .A2(_3092_),
    .B1_N(_3071_),
    .X(_3093_));
 sky130_fd_sc_hd__a22o_2 _7782_ (.A1(_3072_),
    .A2(_3075_),
    .B1(_3087_),
    .B2(_3093_),
    .X(net366));
 sky130_fd_sc_hd__a22o_1 _7783_ (.A1(_2439_),
    .A2(net277),
    .B1(_0766_),
    .B2(net331),
    .X(_3094_));
 sky130_fd_sc_hd__a221o_4 _7784_ (.A1(net294),
    .A2(_0651_),
    .B1(net234),
    .B2(_0194_),
    .C1(_3094_),
    .X(_3095_));
 sky130_fd_sc_hd__a22o_1 _7785_ (.A1(_0910_),
    .A2(net277),
    .B1(_4186_),
    .B2(net331),
    .X(_3096_));
 sky130_fd_sc_hd__a221o_2 _7786_ (.A1(net294),
    .A2(_1894_),
    .B1(net234),
    .B2(_0590_),
    .C1(_3096_),
    .X(_3097_));
 sky130_fd_sc_hd__a22o_1 _7787_ (.A1(_4268_),
    .A2(net234),
    .B1(_4280_),
    .B2(net294),
    .X(_3098_));
 sky130_fd_sc_hd__a221o_2 _7788_ (.A1(net331),
    .A2(_0612_),
    .B1(net277),
    .B2(_4278_),
    .C1(_3098_),
    .X(_3099_));
 sky130_fd_sc_hd__a221o_1 _7789_ (.A1(_3097_),
    .A2(_3080_),
    .B1(_3099_),
    .B2(_3084_),
    .C1(_3086_),
    .X(_3100_));
 sky130_fd_sc_hd__a22o_1 _7790_ (.A1(_0759_),
    .A2(net277),
    .B1(_0111_),
    .B2(net331),
    .X(_3101_));
 sky130_fd_sc_hd__a221o_2 _7791_ (.A1(net294),
    .A2(_0143_),
    .B1(net234),
    .B2(_0108_),
    .C1(_3101_),
    .X(_3102_));
 sky130_fd_sc_hd__buf_4 _7792_ (.A(_3070_),
    .X(_3103_));
 sky130_fd_sc_hd__o21ba_1 _7793_ (.A1(_3089_),
    .A2(_3102_),
    .B1_N(_3103_),
    .X(_3104_));
 sky130_fd_sc_hd__a22o_2 _7794_ (.A1(_3072_),
    .A2(_3095_),
    .B1(_3100_),
    .B2(_3104_),
    .X(net413));
 sky130_fd_sc_hd__a22o_1 _7795_ (.A1(_2439_),
    .A2(net288),
    .B1(_0652_),
    .B2(net295),
    .X(_3105_));
 sky130_fd_sc_hd__a221o_4 _7796_ (.A1(net333),
    .A2(_0767_),
    .B1(net235),
    .B2(_0194_),
    .C1(_3105_),
    .X(_3106_));
 sky130_fd_sc_hd__a22o_1 _7797_ (.A1(_0539_),
    .A2(net288),
    .B1(_1989_),
    .B2(net295),
    .X(_3107_));
 sky130_fd_sc_hd__a221o_4 _7798_ (.A1(net333),
    .A2(_0694_),
    .B1(net235),
    .B2(_0590_),
    .C1(_3107_),
    .X(_3108_));
 sky130_fd_sc_hd__a22o_1 _7799_ (.A1(_4268_),
    .A2(net235),
    .B1(net333),
    .B2(_0613_),
    .X(_3109_));
 sky130_fd_sc_hd__a221o_4 _7800_ (.A1(net295),
    .A2(_4280_),
    .B1(net288),
    .B2(_3081_),
    .C1(_3109_),
    .X(_3110_));
 sky130_fd_sc_hd__a221o_1 _7801_ (.A1(_3108_),
    .A2(_3080_),
    .B1(_3110_),
    .B2(_3084_),
    .C1(_3086_),
    .X(_3111_));
 sky130_fd_sc_hd__a22o_1 _7802_ (.A1(_0759_),
    .A2(net288),
    .B1(_0143_),
    .B2(net295),
    .X(_3112_));
 sky130_fd_sc_hd__a221oi_4 _7803_ (.A1(net333),
    .A2(_0729_),
    .B1(net235),
    .B2(_0108_),
    .C1(_3112_),
    .Y(_3113_));
 sky130_fd_sc_hd__a21oi_1 _7804_ (.A1(_3113_),
    .A2(_3086_),
    .B1(_3071_),
    .Y(_3114_));
 sky130_fd_sc_hd__a22o_2 _7805_ (.A1(_3072_),
    .A2(_3106_),
    .B1(_3111_),
    .B2(_3114_),
    .X(net424));
 sky130_fd_sc_hd__a22o_1 _7806_ (.A1(_2439_),
    .A2(net299),
    .B1(_0651_),
    .B2(net296),
    .X(_3115_));
 sky130_fd_sc_hd__a221o_4 _7807_ (.A1(net236),
    .A2(_0194_),
    .B1(net334),
    .B2(_0766_),
    .C1(_3115_),
    .X(_3116_));
 sky130_fd_sc_hd__a22o_1 _7808_ (.A1(_0538_),
    .A2(net299),
    .B1(_1894_),
    .B2(net296),
    .X(_3117_));
 sky130_fd_sc_hd__a221o_4 _7809_ (.A1(net236),
    .A2(_0590_),
    .B1(net334),
    .B2(_0694_),
    .C1(_3117_),
    .X(_3118_));
 sky130_fd_sc_hd__a22o_1 _7810_ (.A1(_4280_),
    .A2(net296),
    .B1(net299),
    .B2(_4278_),
    .X(_3119_));
 sky130_fd_sc_hd__a221o_4 _7811_ (.A1(net236),
    .A2(_4268_),
    .B1(net334),
    .B2(_0612_),
    .C1(_3119_),
    .X(_3120_));
 sky130_fd_sc_hd__a221o_1 _7812_ (.A1(_3118_),
    .A2(_3080_),
    .B1(_3120_),
    .B2(_3084_),
    .C1(_3086_),
    .X(_3121_));
 sky130_fd_sc_hd__a22o_1 _7813_ (.A1(_0759_),
    .A2(net299),
    .B1(_0143_),
    .B2(net296),
    .X(_3122_));
 sky130_fd_sc_hd__a221oi_4 _7814_ (.A1(net236),
    .A2(_0108_),
    .B1(net334),
    .B2(_0729_),
    .C1(_3122_),
    .Y(_3123_));
 sky130_fd_sc_hd__a21oi_1 _7815_ (.A1(_3123_),
    .A2(_3086_),
    .B1(_3071_),
    .Y(_3124_));
 sky130_fd_sc_hd__a22o_2 _7816_ (.A1(_3072_),
    .A2(_3116_),
    .B1(_3121_),
    .B2(_3124_),
    .X(net435));
 sky130_fd_sc_hd__nor2_1 _7817_ (.A(net310),
    .B(_0198_),
    .Y(_3125_));
 sky130_fd_sc_hd__nor2_1 _7818_ (.A(net297),
    .B(_0855_),
    .Y(_3126_));
 sky130_fd_sc_hd__o21ai_2 _7819_ (.A1(_3125_),
    .A2(_3126_),
    .B1(_0199_),
    .Y(_3127_));
 sky130_fd_sc_hd__o221ai_4 _7820_ (.A1(net237),
    .A2(_0486_),
    .B1(net335),
    .B2(_0654_),
    .C1(_3127_),
    .Y(_3128_));
 sky130_fd_sc_hd__inv_2 _7821_ (.A(_3128_),
    .Y(_3129_));
 sky130_fd_sc_hd__inv_2 _7822_ (.A(net310),
    .Y(_3130_));
 sky130_fd_sc_hd__nand2_1 _7823_ (.A(_3130_),
    .B(_0555_),
    .Y(_3131_));
 sky130_fd_sc_hd__a21o_1 _7824_ (.A1(_3131_),
    .A2(_4275_),
    .B1(\arbiter.slave_sel[1][1] ),
    .X(_3132_));
 sky130_fd_sc_hd__o221a_4 _7825_ (.A1(net237),
    .A2(_1291_),
    .B1(net335),
    .B2(_0614_),
    .C1(_3132_),
    .X(_3133_));
 sky130_fd_sc_hd__clkbuf_8 _7826_ (.A(_3078_),
    .X(_3134_));
 sky130_fd_sc_hd__inv_2 _7827_ (.A(net237),
    .Y(_3135_));
 sky130_fd_sc_hd__inv_2 _7828_ (.A(net335),
    .Y(_3136_));
 sky130_fd_sc_hd__nand2_1 _7829_ (.A(_0800_),
    .B(net310),
    .Y(_3137_));
 sky130_fd_sc_hd__a21o_1 _7830_ (.A1(_3137_),
    .A2(_4131_),
    .B1(_4118_),
    .X(_3138_));
 sky130_fd_sc_hd__o221a_1 _7831_ (.A1(_3135_),
    .A2(_0678_),
    .B1(_3136_),
    .B2(_1133_),
    .C1(_3138_),
    .X(_3139_));
 sky130_fd_sc_hd__clkinv_4 _7832_ (.A(_3139_),
    .Y(_3140_));
 sky130_fd_sc_hd__a221o_1 _7833_ (.A1(_3133_),
    .A2(_3134_),
    .B1(_3140_),
    .B2(_3080_),
    .C1(_3086_),
    .X(_3141_));
 sky130_fd_sc_hd__mux2_1 _7834_ (.A0(_3130_),
    .A1(_4274_),
    .S(_0088_),
    .X(_3142_));
 sky130_fd_sc_hd__buf_8 _7835_ (.A(_0160_),
    .X(_3143_));
 sky130_fd_sc_hd__nor2_1 _7836_ (.A(net335),
    .B(_3143_),
    .Y(_3144_));
 sky130_fd_sc_hd__a221o_4 _7837_ (.A1(_3135_),
    .A2(_0108_),
    .B1(_3142_),
    .B2(_0096_),
    .C1(_3144_),
    .X(_3145_));
 sky130_fd_sc_hd__a21oi_1 _7838_ (.A1(_3145_),
    .A2(_3086_),
    .B1(_3071_),
    .Y(_3146_));
 sky130_fd_sc_hd__a22o_2 _7839_ (.A1(_3072_),
    .A2(_3129_),
    .B1(_3141_),
    .B2(_3146_),
    .X(net446));
 sky130_fd_sc_hd__inv_2 _7840_ (.A(net238),
    .Y(_3147_));
 sky130_fd_sc_hd__inv_2 _7841_ (.A(net336),
    .Y(_3148_));
 sky130_fd_sc_hd__nand2_1 _7842_ (.A(_0090_),
    .B(net321),
    .Y(_3149_));
 sky130_fd_sc_hd__nand2_1 _7843_ (.A(_0088_),
    .B(net298),
    .Y(_3150_));
 sky130_fd_sc_hd__a21o_1 _7844_ (.A1(_3149_),
    .A2(_3150_),
    .B1(\arbiter.slave_sel[2][1] ),
    .X(_3151_));
 sky130_fd_sc_hd__o221a_4 _7845_ (.A1(_3147_),
    .A2(_0107_),
    .B1(_3148_),
    .B2(_0160_),
    .C1(_3151_),
    .X(_3152_));
 sky130_fd_sc_hd__a21o_1 _7846_ (.A1(_3152_),
    .A2(_3085_),
    .B1(_3071_),
    .X(_3153_));
 sky130_fd_sc_hd__nand2_1 _7847_ (.A(_4114_),
    .B(net321),
    .Y(_3154_));
 sky130_fd_sc_hd__nand2_1 _7848_ (.A(_4127_),
    .B(net298),
    .Y(_3155_));
 sky130_fd_sc_hd__a21o_1 _7849_ (.A1(_3154_),
    .A2(_3155_),
    .B1(_4118_),
    .X(_3156_));
 sky130_fd_sc_hd__o221a_2 _7850_ (.A1(_3147_),
    .A2(_0678_),
    .B1(_3148_),
    .B2(_1133_),
    .C1(_3156_),
    .X(_3157_));
 sky130_fd_sc_hd__inv_2 _7851_ (.A(_3157_),
    .Y(_3158_));
 sky130_fd_sc_hd__nand2_1 _7852_ (.A(_4253_),
    .B(net321),
    .Y(_3159_));
 sky130_fd_sc_hd__nand2_1 _7853_ (.A(_4252_),
    .B(net298),
    .Y(_3160_));
 sky130_fd_sc_hd__a21o_1 _7854_ (.A1(_3159_),
    .A2(_3160_),
    .B1(\arbiter.slave_sel[1][1] ),
    .X(_3161_));
 sky130_fd_sc_hd__o221a_2 _7855_ (.A1(_3147_),
    .A2(_4263_),
    .B1(_3148_),
    .B2(_4287_),
    .C1(_3161_),
    .X(_3162_));
 sky130_fd_sc_hd__inv_2 _7856_ (.A(_3162_),
    .Y(_3163_));
 sky130_fd_sc_hd__a221oi_1 _7857_ (.A1(_3158_),
    .A2(_3080_),
    .B1(_3084_),
    .B2(_3163_),
    .C1(_3086_),
    .Y(_3164_));
 sky130_fd_sc_hd__nand2_1 _7858_ (.A(_0195_),
    .B(net321),
    .Y(_3165_));
 sky130_fd_sc_hd__nand2_1 _7859_ (.A(_0198_),
    .B(net298),
    .Y(_3166_));
 sky130_fd_sc_hd__a21o_1 _7860_ (.A1(_3165_),
    .A2(_3166_),
    .B1(\arbiter.slave_sel[3][1] ),
    .X(_3167_));
 sky130_fd_sc_hd__o221a_4 _7861_ (.A1(_3147_),
    .A2(_0486_),
    .B1(_3148_),
    .B2(_0654_),
    .C1(_3167_),
    .X(_3168_));
 sky130_fd_sc_hd__inv_2 _7862_ (.A(_3168_),
    .Y(_3169_));
 sky130_fd_sc_hd__a2bb2o_2 _7863_ (.A1_N(_3153_),
    .A2_N(_3164_),
    .B1(_3072_),
    .B2(_3169_),
    .X(net457));
 sky130_fd_sc_hd__inv_2 _7864_ (.A(net332),
    .Y(_3170_));
 sky130_fd_sc_hd__inv_2 _7865_ (.A(net300),
    .Y(_3171_));
 sky130_fd_sc_hd__o22ai_2 _7866_ (.A1(net239),
    .A2(_0486_),
    .B1(net337),
    .B2(_0654_),
    .Y(_3172_));
 sky130_fd_sc_hd__a221oi_4 _7867_ (.A1(_3170_),
    .A2(_2439_),
    .B1(_3171_),
    .B2(_0652_),
    .C1(_3172_),
    .Y(_3173_));
 sky130_fd_sc_hd__o22ai_2 _7868_ (.A1(net239),
    .A2(_0678_),
    .B1(net337),
    .B2(_1133_),
    .Y(_3174_));
 sky130_fd_sc_hd__a221oi_4 _7869_ (.A1(_3170_),
    .A2(_0539_),
    .B1(_3171_),
    .B2(_1989_),
    .C1(_3174_),
    .Y(_3175_));
 sky130_fd_sc_hd__o22ai_2 _7870_ (.A1(net239),
    .A2(_1291_),
    .B1(net337),
    .B2(_0614_),
    .Y(_3176_));
 sky130_fd_sc_hd__a221oi_4 _7871_ (.A1(_3170_),
    .A2(_3081_),
    .B1(_3171_),
    .B2(_1977_),
    .C1(_3176_),
    .Y(_3177_));
 sky130_fd_sc_hd__clkbuf_8 _7872_ (.A(_3085_),
    .X(_3178_));
 sky130_fd_sc_hd__a221o_1 _7873_ (.A1(_3175_),
    .A2(_3080_),
    .B1(_3177_),
    .B2(_3084_),
    .C1(_3178_),
    .X(_3179_));
 sky130_fd_sc_hd__buf_12 _7874_ (.A(_0759_),
    .X(_3180_));
 sky130_fd_sc_hd__buf_12 _7875_ (.A(_0143_),
    .X(_3181_));
 sky130_fd_sc_hd__buf_8 _7876_ (.A(_0107_),
    .X(_3182_));
 sky130_fd_sc_hd__o22ai_2 _7877_ (.A1(net239),
    .A2(_3182_),
    .B1(net337),
    .B2(_3143_),
    .Y(_3183_));
 sky130_fd_sc_hd__a221oi_4 _7878_ (.A1(_3170_),
    .A2(_3180_),
    .B1(_3171_),
    .B2(_3181_),
    .C1(_3183_),
    .Y(_3184_));
 sky130_fd_sc_hd__o21ba_1 _7879_ (.A1(_3089_),
    .A2(_3184_),
    .B1_N(_3103_),
    .X(_3185_));
 sky130_fd_sc_hd__a22o_2 _7880_ (.A1(_3072_),
    .A2(_3173_),
    .B1(_3179_),
    .B2(_3185_),
    .X(net468));
 sky130_fd_sc_hd__inv_2 _7881_ (.A(net338),
    .Y(_3186_));
 sky130_fd_sc_hd__inv_2 _7882_ (.A(net240),
    .Y(_3187_));
 sky130_fd_sc_hd__inv_2 _7883_ (.A(net343),
    .Y(_3188_));
 sky130_fd_sc_hd__inv_2 _7884_ (.A(net301),
    .Y(_3189_));
 sky130_fd_sc_hd__a22o_1 _7885_ (.A1(_2439_),
    .A2(_3188_),
    .B1(_0652_),
    .B2(_3189_),
    .X(_3190_));
 sky130_fd_sc_hd__a221oi_4 _7886_ (.A1(_3186_),
    .A2(_0767_),
    .B1(_3187_),
    .B2(_0194_),
    .C1(_3190_),
    .Y(_3191_));
 sky130_fd_sc_hd__a22o_1 _7887_ (.A1(_0539_),
    .A2(_3188_),
    .B1(_1989_),
    .B2(_3189_),
    .X(_3192_));
 sky130_fd_sc_hd__a221oi_4 _7888_ (.A1(_3186_),
    .A2(_0694_),
    .B1(_3187_),
    .B2(_0590_),
    .C1(_3192_),
    .Y(_3193_));
 sky130_fd_sc_hd__a22o_1 _7889_ (.A1(_4268_),
    .A2(_3187_),
    .B1(_3186_),
    .B2(_0613_),
    .X(_3194_));
 sky130_fd_sc_hd__a221oi_4 _7890_ (.A1(_3189_),
    .A2(_1977_),
    .B1(_3188_),
    .B2(_3081_),
    .C1(_3194_),
    .Y(_3195_));
 sky130_fd_sc_hd__a221o_1 _7891_ (.A1(_3193_),
    .A2(_3080_),
    .B1(_3195_),
    .B2(_3084_),
    .C1(_3178_),
    .X(_3196_));
 sky130_fd_sc_hd__a22o_1 _7892_ (.A1(_0759_),
    .A2(_3188_),
    .B1(_0109_),
    .B2(_3189_),
    .X(_3197_));
 sky130_fd_sc_hd__a221o_4 _7893_ (.A1(_3186_),
    .A2(_0111_),
    .B1(_3187_),
    .B2(_0108_),
    .C1(_3197_),
    .X(_3198_));
 sky130_fd_sc_hd__a21oi_1 _7894_ (.A1(_3198_),
    .A2(_3086_),
    .B1(_3071_),
    .Y(_3199_));
 sky130_fd_sc_hd__a22o_2 _7895_ (.A1(_3072_),
    .A2(_3191_),
    .B1(_3196_),
    .B2(_3199_),
    .X(net479));
 sky130_fd_sc_hd__inv_2 _7896_ (.A(net354),
    .Y(_3200_));
 sky130_fd_sc_hd__inv_2 _7897_ (.A(net302),
    .Y(_3201_));
 sky130_fd_sc_hd__o22ai_4 _7898_ (.A1(net242),
    .A2(_0193_),
    .B1(net339),
    .B2(_0653_),
    .Y(_3202_));
 sky130_fd_sc_hd__a221oi_4 _7899_ (.A1(_3200_),
    .A2(_0741_),
    .B1(_3201_),
    .B2(_0651_),
    .C1(_3202_),
    .Y(_3203_));
 sky130_fd_sc_hd__o22ai_2 _7900_ (.A1(net242),
    .A2(_0678_),
    .B1(net339),
    .B2(_1133_),
    .Y(_3204_));
 sky130_fd_sc_hd__a221oi_4 _7901_ (.A1(_3200_),
    .A2(_0539_),
    .B1(_3201_),
    .B2(_1989_),
    .C1(_3204_),
    .Y(_3205_));
 sky130_fd_sc_hd__o22ai_2 _7902_ (.A1(net242),
    .A2(_1291_),
    .B1(net339),
    .B2(_0614_),
    .Y(_3206_));
 sky130_fd_sc_hd__a221oi_4 _7903_ (.A1(_3200_),
    .A2(_3081_),
    .B1(_3201_),
    .B2(_1977_),
    .C1(_3206_),
    .Y(_3207_));
 sky130_fd_sc_hd__a221o_1 _7904_ (.A1(_3205_),
    .A2(_3080_),
    .B1(_3207_),
    .B2(_3084_),
    .C1(_3178_),
    .X(_3208_));
 sky130_fd_sc_hd__o22ai_2 _7905_ (.A1(net242),
    .A2(_3182_),
    .B1(net339),
    .B2(_3143_),
    .Y(_3209_));
 sky130_fd_sc_hd__a221oi_4 _7906_ (.A1(_3200_),
    .A2(_0759_),
    .B1(_3201_),
    .B2(_0143_),
    .C1(_3209_),
    .Y(_3210_));
 sky130_fd_sc_hd__o21ba_1 _7907_ (.A1(_3089_),
    .A2(_3210_),
    .B1_N(_3103_),
    .X(_3211_));
 sky130_fd_sc_hd__a22o_2 _7908_ (.A1(_3072_),
    .A2(_3203_),
    .B1(_3208_),
    .B2(_3211_),
    .X(net490));
 sky130_fd_sc_hd__inv_2 _7909_ (.A(net365),
    .Y(_3212_));
 sky130_fd_sc_hd__inv_2 _7910_ (.A(net303),
    .Y(_3213_));
 sky130_fd_sc_hd__o22ai_2 _7911_ (.A1(net243),
    .A2(_0486_),
    .B1(net340),
    .B2(_0654_),
    .Y(_3214_));
 sky130_fd_sc_hd__a221oi_4 _7912_ (.A1(_3212_),
    .A2(_2439_),
    .B1(_3213_),
    .B2(_0652_),
    .C1(_3214_),
    .Y(_3215_));
 sky130_fd_sc_hd__o22ai_2 _7913_ (.A1(net243),
    .A2(_0678_),
    .B1(net340),
    .B2(_1133_),
    .Y(_3216_));
 sky130_fd_sc_hd__a221oi_4 _7914_ (.A1(_3212_),
    .A2(_0539_),
    .B1(_3213_),
    .B2(_1989_),
    .C1(_3216_),
    .Y(_3217_));
 sky130_fd_sc_hd__o22ai_2 _7915_ (.A1(net243),
    .A2(_1291_),
    .B1(net340),
    .B2(_0614_),
    .Y(_3218_));
 sky130_fd_sc_hd__a221oi_4 _7916_ (.A1(_3212_),
    .A2(_4278_),
    .B1(_3213_),
    .B2(_4280_),
    .C1(_3218_),
    .Y(_3219_));
 sky130_fd_sc_hd__a221o_1 _7917_ (.A1(_3217_),
    .A2(_3080_),
    .B1(_3219_),
    .B2(_3084_),
    .C1(_3178_),
    .X(_3220_));
 sky130_fd_sc_hd__o22ai_2 _7918_ (.A1(net243),
    .A2(_0107_),
    .B1(net340),
    .B2(_0160_),
    .Y(_3221_));
 sky130_fd_sc_hd__a221oi_4 _7919_ (.A1(_3212_),
    .A2(_0759_),
    .B1(_3213_),
    .B2(_0143_),
    .C1(_3221_),
    .Y(_3222_));
 sky130_fd_sc_hd__o21ba_1 _7920_ (.A1(_3089_),
    .A2(_3222_),
    .B1_N(_3103_),
    .X(_3223_));
 sky130_fd_sc_hd__a22o_2 _7921_ (.A1(_3072_),
    .A2(_3215_),
    .B1(_3220_),
    .B2(_3223_),
    .X(net501));
 sky130_fd_sc_hd__inv_2 _7922_ (.A(net241),
    .Y(_3224_));
 sky130_fd_sc_hd__clkinv_4 _7923_ (.A(net304),
    .Y(_3225_));
 sky130_fd_sc_hd__o22ai_2 _7924_ (.A1(net244),
    .A2(_0193_),
    .B1(net341),
    .B2(_0653_),
    .Y(_3226_));
 sky130_fd_sc_hd__a221oi_4 _7925_ (.A1(_3224_),
    .A2(_0741_),
    .B1(_3225_),
    .B2(_0196_),
    .C1(_3226_),
    .Y(_3227_));
 sky130_fd_sc_hd__o22ai_4 _7926_ (.A1(net244),
    .A2(_4223_),
    .B1(net341),
    .B2(_1132_),
    .Y(_3228_));
 sky130_fd_sc_hd__a221oi_4 _7927_ (.A1(_3224_),
    .A2(_4204_),
    .B1(_3225_),
    .B2(_4213_),
    .C1(_3228_),
    .Y(_3229_));
 sky130_fd_sc_hd__o22ai_2 _7928_ (.A1(net244),
    .A2(_1291_),
    .B1(net341),
    .B2(_0614_),
    .Y(_3230_));
 sky130_fd_sc_hd__a221oi_4 _7929_ (.A1(_3224_),
    .A2(_3081_),
    .B1(_3225_),
    .B2(_1977_),
    .C1(_3230_),
    .Y(_3231_));
 sky130_fd_sc_hd__a221o_1 _7930_ (.A1(_3229_),
    .A2(_3080_),
    .B1(_3231_),
    .B2(_3084_),
    .C1(_3178_),
    .X(_3232_));
 sky130_fd_sc_hd__o22ai_2 _7931_ (.A1(net244),
    .A2(_3182_),
    .B1(net341),
    .B2(_3143_),
    .Y(_3233_));
 sky130_fd_sc_hd__a221oi_4 _7932_ (.A1(_3224_),
    .A2(_3180_),
    .B1(_3225_),
    .B2(_3181_),
    .C1(_3233_),
    .Y(_3234_));
 sky130_fd_sc_hd__o21ba_1 _7933_ (.A1(_3089_),
    .A2(_3234_),
    .B1_N(_3103_),
    .X(_3235_));
 sky130_fd_sc_hd__a22o_2 _7934_ (.A1(_3072_),
    .A2(_3227_),
    .B1(_3232_),
    .B2(_3235_),
    .X(net377));
 sky130_fd_sc_hd__inv_2 _7935_ (.A(net252),
    .Y(_3236_));
 sky130_fd_sc_hd__clkinv_4 _7936_ (.A(net305),
    .Y(_3237_));
 sky130_fd_sc_hd__o22ai_2 _7937_ (.A1(net245),
    .A2(_0486_),
    .B1(net342),
    .B2(_0654_),
    .Y(_3238_));
 sky130_fd_sc_hd__a221oi_4 _7938_ (.A1(_3236_),
    .A2(_0741_),
    .B1(_3237_),
    .B2(_0651_),
    .C1(_3238_),
    .Y(_3239_));
 sky130_fd_sc_hd__o22ai_2 _7939_ (.A1(net245),
    .A2(_0678_),
    .B1(net342),
    .B2(_1133_),
    .Y(_3240_));
 sky130_fd_sc_hd__a221oi_4 _7940_ (.A1(_3236_),
    .A2(_0539_),
    .B1(_3237_),
    .B2(_1989_),
    .C1(_3240_),
    .Y(_3241_));
 sky130_fd_sc_hd__o22ai_2 _7941_ (.A1(net245),
    .A2(_1291_),
    .B1(net342),
    .B2(_0614_),
    .Y(_3242_));
 sky130_fd_sc_hd__a221oi_4 _7942_ (.A1(_3236_),
    .A2(_3081_),
    .B1(_3237_),
    .B2(_1977_),
    .C1(_3242_),
    .Y(_3243_));
 sky130_fd_sc_hd__a221o_1 _7943_ (.A1(_3241_),
    .A2(_3080_),
    .B1(_3243_),
    .B2(_3084_),
    .C1(_3178_),
    .X(_3244_));
 sky130_fd_sc_hd__o22ai_2 _7944_ (.A1(net245),
    .A2(_3182_),
    .B1(net342),
    .B2(_3143_),
    .Y(_3245_));
 sky130_fd_sc_hd__a221oi_4 _7945_ (.A1(_3236_),
    .A2(_3180_),
    .B1(_3237_),
    .B2(_3181_),
    .C1(_3245_),
    .Y(_3246_));
 sky130_fd_sc_hd__o21ba_1 _7946_ (.A1(_3089_),
    .A2(_3246_),
    .B1_N(_3103_),
    .X(_3247_));
 sky130_fd_sc_hd__a22o_4 _7947_ (.A1(_3072_),
    .A2(_3239_),
    .B1(_3244_),
    .B2(_3247_),
    .X(net388));
 sky130_fd_sc_hd__inv_2 _7948_ (.A(net263),
    .Y(_3248_));
 sky130_fd_sc_hd__inv_2 _7949_ (.A(net306),
    .Y(_3249_));
 sky130_fd_sc_hd__o22ai_2 _7950_ (.A1(net246),
    .A2(_0193_),
    .B1(net344),
    .B2(_0653_),
    .Y(_3250_));
 sky130_fd_sc_hd__a221oi_4 _7951_ (.A1(_3248_),
    .A2(_0741_),
    .B1(_3249_),
    .B2(_0651_),
    .C1(_3250_),
    .Y(_3251_));
 sky130_fd_sc_hd__o22ai_2 _7952_ (.A1(net246),
    .A2(_4223_),
    .B1(net344),
    .B2(_1132_),
    .Y(_3252_));
 sky130_fd_sc_hd__a221oi_4 _7953_ (.A1(_3248_),
    .A2(_4204_),
    .B1(_3249_),
    .B2(_1894_),
    .C1(_3252_),
    .Y(_3253_));
 sky130_fd_sc_hd__clkbuf_8 _7954_ (.A(_3079_),
    .X(_3254_));
 sky130_fd_sc_hd__o22ai_2 _7955_ (.A1(net246),
    .A2(_1291_),
    .B1(net344),
    .B2(_0614_),
    .Y(_3255_));
 sky130_fd_sc_hd__a221oi_4 _7956_ (.A1(_3248_),
    .A2(_3081_),
    .B1(_3249_),
    .B2(_1977_),
    .C1(_3255_),
    .Y(_3256_));
 sky130_fd_sc_hd__a221o_1 _7957_ (.A1(_3253_),
    .A2(_3254_),
    .B1(_3256_),
    .B2(_3084_),
    .C1(_3178_),
    .X(_3257_));
 sky130_fd_sc_hd__o22ai_2 _7958_ (.A1(net246),
    .A2(_3182_),
    .B1(net344),
    .B2(_3143_),
    .Y(_3258_));
 sky130_fd_sc_hd__a221oi_4 _7959_ (.A1(_3248_),
    .A2(_3180_),
    .B1(_3249_),
    .B2(_3181_),
    .C1(_3258_),
    .Y(_3259_));
 sky130_fd_sc_hd__o21ba_1 _7960_ (.A1(_3089_),
    .A2(_3259_),
    .B1_N(_3103_),
    .X(_3260_));
 sky130_fd_sc_hd__a22o_2 _7961_ (.A1(_3072_),
    .A2(_3251_),
    .B1(_3257_),
    .B2(_3260_),
    .X(net399));
 sky130_fd_sc_hd__inv_2 _7962_ (.A(net270),
    .Y(_3261_));
 sky130_fd_sc_hd__inv_2 _7963_ (.A(net307),
    .Y(_3262_));
 sky130_fd_sc_hd__o22ai_2 _7964_ (.A1(net247),
    .A2(_0486_),
    .B1(net345),
    .B2(_0654_),
    .Y(_3263_));
 sky130_fd_sc_hd__a221oi_4 _7965_ (.A1(_3261_),
    .A2(_0741_),
    .B1(_3262_),
    .B2(_0651_),
    .C1(_3263_),
    .Y(_3264_));
 sky130_fd_sc_hd__o22ai_2 _7966_ (.A1(net247),
    .A2(_0678_),
    .B1(net345),
    .B2(_1133_),
    .Y(_3265_));
 sky130_fd_sc_hd__a221oi_4 _7967_ (.A1(_3261_),
    .A2(_0538_),
    .B1(_3262_),
    .B2(_1894_),
    .C1(_3265_),
    .Y(_3266_));
 sky130_fd_sc_hd__o22ai_2 _7968_ (.A1(net247),
    .A2(_1291_),
    .B1(net345),
    .B2(_0614_),
    .Y(_3267_));
 sky130_fd_sc_hd__a221oi_4 _7969_ (.A1(_3261_),
    .A2(_3081_),
    .B1(_3262_),
    .B2(_1977_),
    .C1(_3267_),
    .Y(_3268_));
 sky130_fd_sc_hd__a221o_1 _7970_ (.A1(_3266_),
    .A2(_3254_),
    .B1(_3268_),
    .B2(_3084_),
    .C1(_3178_),
    .X(_3269_));
 sky130_fd_sc_hd__o22ai_4 _7971_ (.A1(net247),
    .A2(_3182_),
    .B1(net345),
    .B2(_3143_),
    .Y(_3270_));
 sky130_fd_sc_hd__a221oi_4 _7972_ (.A1(_3261_),
    .A2(_3180_),
    .B1(_3262_),
    .B2(_3181_),
    .C1(_3270_),
    .Y(_3271_));
 sky130_fd_sc_hd__o21ba_1 _7973_ (.A1(_3089_),
    .A2(_3271_),
    .B1_N(_3103_),
    .X(_3272_));
 sky130_fd_sc_hd__a22o_2 _7974_ (.A1(_3072_),
    .A2(_3264_),
    .B1(_3269_),
    .B2(_3272_),
    .X(net406));
 sky130_fd_sc_hd__buf_6 _7975_ (.A(_3071_),
    .X(_3273_));
 sky130_fd_sc_hd__clkinv_4 _7976_ (.A(net308),
    .Y(_3274_));
 sky130_fd_sc_hd__inv_2 _7977_ (.A(net271),
    .Y(_3275_));
 sky130_fd_sc_hd__o22ai_2 _7978_ (.A1(net248),
    .A2(_0486_),
    .B1(net346),
    .B2(_0654_),
    .Y(_3276_));
 sky130_fd_sc_hd__a221oi_4 _7979_ (.A1(_3274_),
    .A2(_0651_),
    .B1(_3275_),
    .B2(_0741_),
    .C1(_3276_),
    .Y(_3277_));
 sky130_fd_sc_hd__o22ai_2 _7980_ (.A1(net248),
    .A2(_0678_),
    .B1(net346),
    .B2(_1133_),
    .Y(_3278_));
 sky130_fd_sc_hd__a221oi_4 _7981_ (.A1(_3274_),
    .A2(_1894_),
    .B1(_3275_),
    .B2(_0538_),
    .C1(_3278_),
    .Y(_3279_));
 sky130_fd_sc_hd__o22ai_2 _7982_ (.A1(net248),
    .A2(_1291_),
    .B1(net346),
    .B2(_0614_),
    .Y(_3280_));
 sky130_fd_sc_hd__a221oi_4 _7983_ (.A1(_3274_),
    .A2(_1977_),
    .B1(_3275_),
    .B2(_3081_),
    .C1(_3280_),
    .Y(_3281_));
 sky130_fd_sc_hd__a221o_1 _7984_ (.A1(_3279_),
    .A2(_3254_),
    .B1(_3281_),
    .B2(_3084_),
    .C1(_3178_),
    .X(_3282_));
 sky130_fd_sc_hd__o22ai_2 _7985_ (.A1(net248),
    .A2(_3182_),
    .B1(net346),
    .B2(_3143_),
    .Y(_3283_));
 sky130_fd_sc_hd__a221oi_4 _7986_ (.A1(_3274_),
    .A2(_3181_),
    .B1(_3275_),
    .B2(_3180_),
    .C1(_3283_),
    .Y(_3284_));
 sky130_fd_sc_hd__o21ba_1 _7987_ (.A1(_3089_),
    .A2(_3284_),
    .B1_N(_3103_),
    .X(_3285_));
 sky130_fd_sc_hd__a22o_2 _7988_ (.A1(_3273_),
    .A2(_3277_),
    .B1(_3282_),
    .B2(_3285_),
    .X(net407));
 sky130_fd_sc_hd__inv_2 _7989_ (.A(net309),
    .Y(_3286_));
 sky130_fd_sc_hd__inv_2 _7990_ (.A(net272),
    .Y(_3287_));
 sky130_fd_sc_hd__o22ai_2 _7991_ (.A1(net249),
    .A2(_0193_),
    .B1(net347),
    .B2(_0653_),
    .Y(_3288_));
 sky130_fd_sc_hd__a221oi_4 _7992_ (.A1(_3286_),
    .A2(_0651_),
    .B1(_3287_),
    .B2(_0741_),
    .C1(_3288_),
    .Y(_3289_));
 sky130_fd_sc_hd__o22ai_2 _7993_ (.A1(net249),
    .A2(_0678_),
    .B1(net347),
    .B2(_1133_),
    .Y(_3290_));
 sky130_fd_sc_hd__a221oi_4 _7994_ (.A1(_3286_),
    .A2(_1894_),
    .B1(_3287_),
    .B2(_0538_),
    .C1(_3290_),
    .Y(_3291_));
 sky130_fd_sc_hd__o22ai_4 _7995_ (.A1(net249),
    .A2(_4263_),
    .B1(net347),
    .B2(_4287_),
    .Y(_3292_));
 sky130_fd_sc_hd__a221oi_4 _7996_ (.A1(_3286_),
    .A2(_4280_),
    .B1(_3287_),
    .B2(_4278_),
    .C1(_3292_),
    .Y(_3293_));
 sky130_fd_sc_hd__a221o_1 _7997_ (.A1(_3291_),
    .A2(_3254_),
    .B1(_3293_),
    .B2(_3134_),
    .C1(_3178_),
    .X(_3294_));
 sky130_fd_sc_hd__o22ai_2 _7998_ (.A1(net249),
    .A2(_3182_),
    .B1(net347),
    .B2(_3143_),
    .Y(_3295_));
 sky130_fd_sc_hd__a221oi_4 _7999_ (.A1(_3286_),
    .A2(_3181_),
    .B1(_3287_),
    .B2(_3180_),
    .C1(_3295_),
    .Y(_3296_));
 sky130_fd_sc_hd__o21ba_1 _8000_ (.A1(_3089_),
    .A2(_3296_),
    .B1_N(_3103_),
    .X(_3297_));
 sky130_fd_sc_hd__a22o_4 _8001_ (.A1(_3273_),
    .A2(_3289_),
    .B1(_3294_),
    .B2(_3297_),
    .X(net408));
 sky130_fd_sc_hd__inv_2 _8002_ (.A(net273),
    .Y(_3298_));
 sky130_fd_sc_hd__inv_2 _8003_ (.A(net311),
    .Y(_3299_));
 sky130_fd_sc_hd__o22ai_2 _8004_ (.A1(net250),
    .A2(_0193_),
    .B1(net348),
    .B2(_0653_),
    .Y(_3300_));
 sky130_fd_sc_hd__a221oi_4 _8005_ (.A1(_3298_),
    .A2(_0741_),
    .B1(_3299_),
    .B2(_0196_),
    .C1(_3300_),
    .Y(_3301_));
 sky130_fd_sc_hd__o22ai_2 _8006_ (.A1(net250),
    .A2(_0678_),
    .B1(net348),
    .B2(_1133_),
    .Y(_3302_));
 sky130_fd_sc_hd__a221oi_4 _8007_ (.A1(_3298_),
    .A2(_0538_),
    .B1(_3299_),
    .B2(_1894_),
    .C1(_3302_),
    .Y(_3303_));
 sky130_fd_sc_hd__o22ai_2 _8008_ (.A1(net250),
    .A2(_1291_),
    .B1(net348),
    .B2(_0614_),
    .Y(_3304_));
 sky130_fd_sc_hd__a221oi_4 _8009_ (.A1(_3298_),
    .A2(_3081_),
    .B1(_3299_),
    .B2(_1977_),
    .C1(_3304_),
    .Y(_3305_));
 sky130_fd_sc_hd__a221o_1 _8010_ (.A1(_3303_),
    .A2(_3254_),
    .B1(_3305_),
    .B2(_3134_),
    .C1(_3178_),
    .X(_3306_));
 sky130_fd_sc_hd__o22ai_2 _8011_ (.A1(net250),
    .A2(_3182_),
    .B1(net348),
    .B2(_3143_),
    .Y(_3307_));
 sky130_fd_sc_hd__a221oi_4 _8012_ (.A1(_3298_),
    .A2(_3180_),
    .B1(_3299_),
    .B2(_3181_),
    .C1(_3307_),
    .Y(_3308_));
 sky130_fd_sc_hd__o21ba_1 _8013_ (.A1(_3089_),
    .A2(_3308_),
    .B1_N(_3103_),
    .X(_3309_));
 sky130_fd_sc_hd__a22o_2 _8014_ (.A1(_3273_),
    .A2(_3301_),
    .B1(_3306_),
    .B2(_3309_),
    .X(net409));
 sky130_fd_sc_hd__inv_2 _8015_ (.A(net274),
    .Y(_3310_));
 sky130_fd_sc_hd__inv_2 _8016_ (.A(net312),
    .Y(_3311_));
 sky130_fd_sc_hd__o22ai_2 _8017_ (.A1(net251),
    .A2(_0486_),
    .B1(net349),
    .B2(_0654_),
    .Y(_3312_));
 sky130_fd_sc_hd__a221oi_4 _8018_ (.A1(_3310_),
    .A2(_0741_),
    .B1(_3311_),
    .B2(_0651_),
    .C1(_3312_),
    .Y(_3313_));
 sky130_fd_sc_hd__o22ai_4 _8019_ (.A1(net251),
    .A2(_4223_),
    .B1(net349),
    .B2(_1132_),
    .Y(_3314_));
 sky130_fd_sc_hd__a221oi_4 _8020_ (.A1(_3310_),
    .A2(_0910_),
    .B1(_3311_),
    .B2(_1894_),
    .C1(_3314_),
    .Y(_3315_));
 sky130_fd_sc_hd__o22ai_2 _8021_ (.A1(net251),
    .A2(_4263_),
    .B1(net349),
    .B2(_4287_),
    .Y(_3316_));
 sky130_fd_sc_hd__a221oi_4 _8022_ (.A1(_3310_),
    .A2(_4278_),
    .B1(_3311_),
    .B2(_4280_),
    .C1(_3316_),
    .Y(_3317_));
 sky130_fd_sc_hd__a221o_1 _8023_ (.A1(_3315_),
    .A2(_3254_),
    .B1(_3317_),
    .B2(_3134_),
    .C1(_3178_),
    .X(_3318_));
 sky130_fd_sc_hd__o22ai_2 _8024_ (.A1(net251),
    .A2(_3182_),
    .B1(net349),
    .B2(_3143_),
    .Y(_3319_));
 sky130_fd_sc_hd__a221oi_4 _8025_ (.A1(_3310_),
    .A2(_3180_),
    .B1(_3311_),
    .B2(_3181_),
    .C1(_3319_),
    .Y(_3320_));
 sky130_fd_sc_hd__o21ba_1 _8026_ (.A1(_3089_),
    .A2(_3320_),
    .B1_N(_3103_),
    .X(_3321_));
 sky130_fd_sc_hd__a22o_4 _8027_ (.A1(_3273_),
    .A2(_3313_),
    .B1(_3318_),
    .B2(_3321_),
    .X(net410));
 sky130_fd_sc_hd__inv_2 _8028_ (.A(net253),
    .Y(_3322_));
 sky130_fd_sc_hd__inv_2 _8029_ (.A(net350),
    .Y(_3323_));
 sky130_fd_sc_hd__inv_2 _8030_ (.A(net275),
    .Y(_3324_));
 sky130_fd_sc_hd__inv_2 _8031_ (.A(net313),
    .Y(_3325_));
 sky130_fd_sc_hd__a22o_1 _8032_ (.A1(_0192_),
    .A2(_3324_),
    .B1(_0196_),
    .B2(_3325_),
    .X(_3326_));
 sky130_fd_sc_hd__a221oi_4 _8033_ (.A1(_3322_),
    .A2(_0194_),
    .B1(_3323_),
    .B2(_0200_),
    .C1(_3326_),
    .Y(_3327_));
 sky130_fd_sc_hd__a22o_1 _8034_ (.A1(_4204_),
    .A2(_3324_),
    .B1(_4213_),
    .B2(_3325_),
    .X(_3328_));
 sky130_fd_sc_hd__a221o_1 _8035_ (.A1(_3322_),
    .A2(_0590_),
    .B1(_3323_),
    .B2(_4186_),
    .C1(_3328_),
    .X(_3329_));
 sky130_fd_sc_hd__inv_2 _8036_ (.A(_3329_),
    .Y(_3330_));
 sky130_fd_sc_hd__a22o_1 _8037_ (.A1(_4280_),
    .A2(_3325_),
    .B1(_3324_),
    .B2(_4278_),
    .X(_3331_));
 sky130_fd_sc_hd__a221o_2 _8038_ (.A1(_3322_),
    .A2(_4268_),
    .B1(_3323_),
    .B2(_4265_),
    .C1(_3331_),
    .X(_3332_));
 sky130_fd_sc_hd__inv_2 _8039_ (.A(_3332_),
    .Y(_3333_));
 sky130_fd_sc_hd__a221o_1 _8040_ (.A1(_3330_),
    .A2(_3254_),
    .B1(_3333_),
    .B2(_3134_),
    .C1(_3178_),
    .X(_3334_));
 sky130_fd_sc_hd__a22o_1 _8041_ (.A1(_3180_),
    .A2(_3324_),
    .B1(_3181_),
    .B2(_3325_),
    .X(_3335_));
 sky130_fd_sc_hd__a221oi_4 _8042_ (.A1(_3322_),
    .A2(_0108_),
    .B1(_3323_),
    .B2(_0572_),
    .C1(_3335_),
    .Y(_3336_));
 sky130_fd_sc_hd__o21ba_1 _8043_ (.A1(_3089_),
    .A2(_3336_),
    .B1_N(_3103_),
    .X(_3337_));
 sky130_fd_sc_hd__a22o_4 _8044_ (.A1(_3273_),
    .A2(_3327_),
    .B1(_3334_),
    .B2(_3337_),
    .X(net411));
 sky130_fd_sc_hd__inv_2 _8045_ (.A(net276),
    .Y(_3338_));
 sky130_fd_sc_hd__inv_2 _8046_ (.A(net314),
    .Y(_3339_));
 sky130_fd_sc_hd__o22ai_2 _8047_ (.A1(net254),
    .A2(_0486_),
    .B1(net351),
    .B2(_0654_),
    .Y(_3340_));
 sky130_fd_sc_hd__a221oi_4 _8048_ (.A1(_3338_),
    .A2(_0741_),
    .B1(_3339_),
    .B2(_0651_),
    .C1(_3340_),
    .Y(_3341_));
 sky130_fd_sc_hd__o22ai_2 _8049_ (.A1(net254),
    .A2(_4223_),
    .B1(net351),
    .B2(_1132_),
    .Y(_3342_));
 sky130_fd_sc_hd__a221oi_4 _8050_ (.A1(_3338_),
    .A2(_0910_),
    .B1(_3339_),
    .B2(_1894_),
    .C1(_3342_),
    .Y(_3343_));
 sky130_fd_sc_hd__o22ai_2 _8051_ (.A1(net254),
    .A2(_1291_),
    .B1(net351),
    .B2(_0614_),
    .Y(_3344_));
 sky130_fd_sc_hd__a221oi_4 _8052_ (.A1(_3338_),
    .A2(_4278_),
    .B1(_3339_),
    .B2(_4280_),
    .C1(_3344_),
    .Y(_3345_));
 sky130_fd_sc_hd__a221o_1 _8053_ (.A1(_3343_),
    .A2(_3254_),
    .B1(_3345_),
    .B2(_3134_),
    .C1(_3178_),
    .X(_3346_));
 sky130_fd_sc_hd__o22ai_2 _8054_ (.A1(net254),
    .A2(_3182_),
    .B1(net351),
    .B2(_3143_),
    .Y(_3347_));
 sky130_fd_sc_hd__a221oi_4 _8055_ (.A1(_3338_),
    .A2(_3180_),
    .B1(_3339_),
    .B2(_3181_),
    .C1(_3347_),
    .Y(_3348_));
 sky130_fd_sc_hd__o21ba_1 _8056_ (.A1(_3089_),
    .A2(_3348_),
    .B1_N(_3103_),
    .X(_3349_));
 sky130_fd_sc_hd__a22o_4 _8057_ (.A1(_3273_),
    .A2(_3341_),
    .B1(_3346_),
    .B2(_3349_),
    .X(net412));
 sky130_fd_sc_hd__inv_2 _8058_ (.A(net278),
    .Y(_3350_));
 sky130_fd_sc_hd__inv_2 _8059_ (.A(net315),
    .Y(_3351_));
 sky130_fd_sc_hd__o22ai_2 _8060_ (.A1(net255),
    .A2(_0193_),
    .B1(net352),
    .B2(_0653_),
    .Y(_3352_));
 sky130_fd_sc_hd__a221oi_4 _8061_ (.A1(_3350_),
    .A2(_0741_),
    .B1(_3351_),
    .B2(_0196_),
    .C1(_3352_),
    .Y(_3353_));
 sky130_fd_sc_hd__o22ai_2 _8062_ (.A1(net255),
    .A2(_0678_),
    .B1(net352),
    .B2(_1133_),
    .Y(_3354_));
 sky130_fd_sc_hd__a221oi_4 _8063_ (.A1(_3350_),
    .A2(_0539_),
    .B1(_3351_),
    .B2(_1989_),
    .C1(_3354_),
    .Y(_3355_));
 sky130_fd_sc_hd__o22ai_4 _8064_ (.A1(net255),
    .A2(_4263_),
    .B1(net352),
    .B2(_4287_),
    .Y(_3356_));
 sky130_fd_sc_hd__a221oi_4 _8065_ (.A1(_3350_),
    .A2(_4278_),
    .B1(_3351_),
    .B2(_4280_),
    .C1(_3356_),
    .Y(_3357_));
 sky130_fd_sc_hd__a221o_1 _8066_ (.A1(_3355_),
    .A2(_3254_),
    .B1(_3357_),
    .B2(_3134_),
    .C1(_3178_),
    .X(_3358_));
 sky130_fd_sc_hd__o22ai_2 _8067_ (.A1(net255),
    .A2(_3182_),
    .B1(net352),
    .B2(_3143_),
    .Y(_3359_));
 sky130_fd_sc_hd__a221oi_4 _8068_ (.A1(_3350_),
    .A2(_3180_),
    .B1(_3351_),
    .B2(_3181_),
    .C1(_3359_),
    .Y(_3360_));
 sky130_fd_sc_hd__o21ba_1 _8069_ (.A1(_3089_),
    .A2(_3360_),
    .B1_N(_3103_),
    .X(_3361_));
 sky130_fd_sc_hd__a22o_2 _8070_ (.A1(_3273_),
    .A2(_3353_),
    .B1(_3358_),
    .B2(_3361_),
    .X(net414));
 sky130_fd_sc_hd__inv_2 _8071_ (.A(net279),
    .Y(_3362_));
 sky130_fd_sc_hd__inv_2 _8072_ (.A(net316),
    .Y(_3363_));
 sky130_fd_sc_hd__o22ai_2 _8073_ (.A1(net256),
    .A2(_0486_),
    .B1(net353),
    .B2(_0654_),
    .Y(_3364_));
 sky130_fd_sc_hd__a221oi_4 _8074_ (.A1(_3362_),
    .A2(_0741_),
    .B1(_3363_),
    .B2(_0651_),
    .C1(_3364_),
    .Y(_3365_));
 sky130_fd_sc_hd__o22ai_2 _8075_ (.A1(net256),
    .A2(_4223_),
    .B1(net353),
    .B2(_1132_),
    .Y(_3366_));
 sky130_fd_sc_hd__a221oi_4 _8076_ (.A1(_3362_),
    .A2(_0910_),
    .B1(_3363_),
    .B2(_1894_),
    .C1(_3366_),
    .Y(_3367_));
 sky130_fd_sc_hd__o22ai_2 _8077_ (.A1(net256),
    .A2(_4263_),
    .B1(net353),
    .B2(_4287_),
    .Y(_3368_));
 sky130_fd_sc_hd__a221oi_4 _8078_ (.A1(_3362_),
    .A2(_4278_),
    .B1(_3363_),
    .B2(_4280_),
    .C1(_3368_),
    .Y(_3369_));
 sky130_fd_sc_hd__a221o_1 _8079_ (.A1(_3367_),
    .A2(_3254_),
    .B1(_3369_),
    .B2(_3134_),
    .C1(_3178_),
    .X(_3370_));
 sky130_fd_sc_hd__o22ai_2 _8080_ (.A1(net256),
    .A2(_3182_),
    .B1(net353),
    .B2(_3143_),
    .Y(_3371_));
 sky130_fd_sc_hd__a221oi_4 _8081_ (.A1(_3362_),
    .A2(_3180_),
    .B1(_3363_),
    .B2(_3181_),
    .C1(_3371_),
    .Y(_3372_));
 sky130_fd_sc_hd__o21ba_1 _8082_ (.A1(_3088_),
    .A2(_3372_),
    .B1_N(_3103_),
    .X(_3373_));
 sky130_fd_sc_hd__a22o_4 _8083_ (.A1(_3273_),
    .A2(_3365_),
    .B1(_3370_),
    .B2(_3373_),
    .X(net415));
 sky130_fd_sc_hd__inv_2 _8084_ (.A(net317),
    .Y(_3374_));
 sky130_fd_sc_hd__inv_2 _8085_ (.A(net280),
    .Y(_3375_));
 sky130_fd_sc_hd__o22ai_2 _8086_ (.A1(net257),
    .A2(_0193_),
    .B1(net355),
    .B2(_0653_),
    .Y(_3376_));
 sky130_fd_sc_hd__a221oi_4 _8087_ (.A1(_3374_),
    .A2(_0196_),
    .B1(_3375_),
    .B2(_0741_),
    .C1(_3376_),
    .Y(_3377_));
 sky130_fd_sc_hd__o22ai_2 _8088_ (.A1(net257),
    .A2(_0678_),
    .B1(net355),
    .B2(_1133_),
    .Y(_3378_));
 sky130_fd_sc_hd__a221oi_4 _8089_ (.A1(_3374_),
    .A2(_1894_),
    .B1(_3375_),
    .B2(_0538_),
    .C1(_3378_),
    .Y(_3379_));
 sky130_fd_sc_hd__o22ai_2 _8090_ (.A1(net257),
    .A2(_1291_),
    .B1(net355),
    .B2(_0614_),
    .Y(_3380_));
 sky130_fd_sc_hd__a221oi_4 _8091_ (.A1(_3374_),
    .A2(_1977_),
    .B1(_3375_),
    .B2(_3081_),
    .C1(_3380_),
    .Y(_3381_));
 sky130_fd_sc_hd__a221o_1 _8092_ (.A1(_3379_),
    .A2(_3254_),
    .B1(_3381_),
    .B2(_3134_),
    .C1(_3085_),
    .X(_3382_));
 sky130_fd_sc_hd__o22ai_1 _8093_ (.A1(net257),
    .A2(_3182_),
    .B1(net355),
    .B2(_0160_),
    .Y(_3383_));
 sky130_fd_sc_hd__a221oi_1 _8094_ (.A1(_3374_),
    .A2(_0143_),
    .B1(_3375_),
    .B2(_0759_),
    .C1(_3383_),
    .Y(_3384_));
 sky130_fd_sc_hd__o21ba_1 _8095_ (.A1(_3088_),
    .A2(net731),
    .B1_N(_3070_),
    .X(_3385_));
 sky130_fd_sc_hd__a22o_2 _8096_ (.A1(_3273_),
    .A2(_3377_),
    .B1(_3382_),
    .B2(_3385_),
    .X(net416));
 sky130_fd_sc_hd__inv_2 _8097_ (.A(net318),
    .Y(_3386_));
 sky130_fd_sc_hd__inv_2 _8098_ (.A(net281),
    .Y(_3387_));
 sky130_fd_sc_hd__o22ai_4 _8099_ (.A1(net258),
    .A2(_0486_),
    .B1(net356),
    .B2(_0654_),
    .Y(_3388_));
 sky130_fd_sc_hd__a221oi_4 _8100_ (.A1(_3386_),
    .A2(_0651_),
    .B1(_3387_),
    .B2(_0741_),
    .C1(_3388_),
    .Y(_3389_));
 sky130_fd_sc_hd__o22ai_4 _8101_ (.A1(net258),
    .A2(_0678_),
    .B1(net356),
    .B2(_1132_),
    .Y(_3390_));
 sky130_fd_sc_hd__a221oi_4 _8102_ (.A1(_3386_),
    .A2(_1894_),
    .B1(_3387_),
    .B2(_0538_),
    .C1(_3390_),
    .Y(_3391_));
 sky130_fd_sc_hd__o22ai_2 _8103_ (.A1(net258),
    .A2(_1291_),
    .B1(net356),
    .B2(_0614_),
    .Y(_3392_));
 sky130_fd_sc_hd__a221oi_4 _8104_ (.A1(_3386_),
    .A2(_1977_),
    .B1(_3387_),
    .B2(_3081_),
    .C1(_3392_),
    .Y(_3393_));
 sky130_fd_sc_hd__a221o_1 _8105_ (.A1(_3391_),
    .A2(_3254_),
    .B1(_3393_),
    .B2(_3134_),
    .C1(_3085_),
    .X(_3394_));
 sky130_fd_sc_hd__o22ai_4 _8106_ (.A1(net258),
    .A2(_3182_),
    .B1(net356),
    .B2(_3143_),
    .Y(_3395_));
 sky130_fd_sc_hd__a221oi_4 _8107_ (.A1(_3386_),
    .A2(_3181_),
    .B1(_3387_),
    .B2(_3180_),
    .C1(_3395_),
    .Y(_3396_));
 sky130_fd_sc_hd__o21ba_1 _8108_ (.A1(_3088_),
    .A2(_3396_),
    .B1_N(_3070_),
    .X(_3397_));
 sky130_fd_sc_hd__a22o_2 _8109_ (.A1(_3273_),
    .A2(_3389_),
    .B1(_3394_),
    .B2(_3397_),
    .X(net417));
 sky130_fd_sc_hd__inv_2 _8110_ (.A(net282),
    .Y(_3398_));
 sky130_fd_sc_hd__clkinv_4 _8111_ (.A(net319),
    .Y(_3399_));
 sky130_fd_sc_hd__o22ai_2 _8112_ (.A1(net259),
    .A2(_0486_),
    .B1(net357),
    .B2(_0654_),
    .Y(_3400_));
 sky130_fd_sc_hd__a221oi_4 _8113_ (.A1(_3398_),
    .A2(_2439_),
    .B1(_3399_),
    .B2(_0652_),
    .C1(_3400_),
    .Y(_3401_));
 sky130_fd_sc_hd__o22ai_2 _8114_ (.A1(net259),
    .A2(_0678_),
    .B1(net357),
    .B2(_1133_),
    .Y(_3402_));
 sky130_fd_sc_hd__a221oi_4 _8115_ (.A1(_3398_),
    .A2(_0539_),
    .B1(_3399_),
    .B2(_1989_),
    .C1(_3402_),
    .Y(_3403_));
 sky130_fd_sc_hd__o22ai_2 _8116_ (.A1(net259),
    .A2(_1291_),
    .B1(net357),
    .B2(_0614_),
    .Y(_3404_));
 sky130_fd_sc_hd__a221oi_4 _8117_ (.A1(_3398_),
    .A2(_3081_),
    .B1(_3399_),
    .B2(_1977_),
    .C1(_3404_),
    .Y(_3405_));
 sky130_fd_sc_hd__a221o_1 _8118_ (.A1(_3403_),
    .A2(_3254_),
    .B1(_3405_),
    .B2(_3134_),
    .C1(_3085_),
    .X(_3406_));
 sky130_fd_sc_hd__o22ai_2 _8119_ (.A1(net259),
    .A2(_3182_),
    .B1(net357),
    .B2(_3143_),
    .Y(_3407_));
 sky130_fd_sc_hd__a221oi_4 _8120_ (.A1(_3398_),
    .A2(_0759_),
    .B1(_3399_),
    .B2(_0143_),
    .C1(_3407_),
    .Y(_3408_));
 sky130_fd_sc_hd__o21ba_1 _8121_ (.A1(_3088_),
    .A2(_3408_),
    .B1_N(_3070_),
    .X(_3409_));
 sky130_fd_sc_hd__a22o_2 _8122_ (.A1(_3273_),
    .A2(_3401_),
    .B1(_3406_),
    .B2(_3409_),
    .X(net418));
 sky130_fd_sc_hd__inv_2 _8123_ (.A(net283),
    .Y(_3410_));
 sky130_fd_sc_hd__inv_2 _8124_ (.A(net320),
    .Y(_3411_));
 sky130_fd_sc_hd__o22ai_2 _8125_ (.A1(net260),
    .A2(_0486_),
    .B1(net358),
    .B2(_0654_),
    .Y(_3412_));
 sky130_fd_sc_hd__a221oi_4 _8126_ (.A1(_3410_),
    .A2(_2439_),
    .B1(_3411_),
    .B2(_0651_),
    .C1(_3412_),
    .Y(_3413_));
 sky130_fd_sc_hd__o22ai_2 _8127_ (.A1(net260),
    .A2(_0678_),
    .B1(net358),
    .B2(_1133_),
    .Y(_3414_));
 sky130_fd_sc_hd__a221oi_4 _8128_ (.A1(_3410_),
    .A2(_0539_),
    .B1(_3411_),
    .B2(_1989_),
    .C1(_3414_),
    .Y(_3415_));
 sky130_fd_sc_hd__o22ai_2 _8129_ (.A1(net260),
    .A2(_1291_),
    .B1(net358),
    .B2(_0614_),
    .Y(_3416_));
 sky130_fd_sc_hd__a221oi_4 _8130_ (.A1(_3410_),
    .A2(_4278_),
    .B1(_3411_),
    .B2(_4280_),
    .C1(_3416_),
    .Y(_3417_));
 sky130_fd_sc_hd__a221o_1 _8131_ (.A1(_3415_),
    .A2(_3254_),
    .B1(_3417_),
    .B2(_3134_),
    .C1(_3085_),
    .X(_3418_));
 sky130_fd_sc_hd__o22ai_2 _8132_ (.A1(net260),
    .A2(_0107_),
    .B1(net358),
    .B2(_0160_),
    .Y(_3419_));
 sky130_fd_sc_hd__a221oi_4 _8133_ (.A1(_3410_),
    .A2(_0759_),
    .B1(_3411_),
    .B2(_0143_),
    .C1(_3419_),
    .Y(_3420_));
 sky130_fd_sc_hd__o21ba_1 _8134_ (.A1(_3088_),
    .A2(_3420_),
    .B1_N(_3070_),
    .X(_3421_));
 sky130_fd_sc_hd__a22o_2 _8135_ (.A1(_3273_),
    .A2(_3413_),
    .B1(_3418_),
    .B2(_3421_),
    .X(net419));
 sky130_fd_sc_hd__o22a_1 _8136_ (.A1(net261),
    .A2(_0486_),
    .B1(net359),
    .B2(_0654_),
    .X(_3422_));
 sky130_fd_sc_hd__o221a_4 _8137_ (.A1(net284),
    .A2(_0888_),
    .B1(net322),
    .B2(_0197_),
    .C1(_3422_),
    .X(_3423_));
 sky130_fd_sc_hd__inv_2 _8138_ (.A(net359),
    .Y(_3424_));
 sky130_fd_sc_hd__nor2_1 _8139_ (.A(_0522_),
    .B(_3424_),
    .Y(_3425_));
 sky130_fd_sc_hd__nand2_1 _8140_ (.A(_0522_),
    .B(net261),
    .Y(_3426_));
 sky130_fd_sc_hd__nand2_1 _8141_ (.A(_3426_),
    .B(_4118_),
    .Y(_3427_));
 sky130_fd_sc_hd__inv_2 _8142_ (.A(net322),
    .Y(_3428_));
 sky130_fd_sc_hd__nand2_1 _8143_ (.A(_1989_),
    .B(_3428_),
    .Y(_3429_));
 sky130_fd_sc_hd__o221ai_2 _8144_ (.A1(net284),
    .A2(_0520_),
    .B1(_3425_),
    .B2(_3427_),
    .C1(_3429_),
    .Y(_3430_));
 sky130_fd_sc_hd__inv_2 _8145_ (.A(_3430_),
    .Y(_3431_));
 sky130_fd_sc_hd__nor2_1 _8146_ (.A(_0558_),
    .B(_3424_),
    .Y(_3432_));
 sky130_fd_sc_hd__a211o_1 _8147_ (.A1(net261),
    .A2(_0558_),
    .B1(_4245_),
    .C1(_3432_),
    .X(_3433_));
 sky130_fd_sc_hd__o221a_4 _8148_ (.A1(net284),
    .A2(_0785_),
    .B1(net322),
    .B2(_4271_),
    .C1(_3433_),
    .X(_3434_));
 sky130_fd_sc_hd__a221o_1 _8149_ (.A1(_3431_),
    .A2(_3254_),
    .B1(_3434_),
    .B2(_3134_),
    .C1(_3085_),
    .X(_3435_));
 sky130_fd_sc_hd__nand2_1 _8150_ (.A(_0090_),
    .B(net359),
    .Y(_3436_));
 sky130_fd_sc_hd__nand2_1 _8151_ (.A(net261),
    .B(_0730_),
    .Y(_3437_));
 sky130_fd_sc_hd__a2bb2o_1 _8152_ (.A1_N(net284),
    .A2_N(_0844_),
    .B1(_3428_),
    .B2(_0143_),
    .X(_3438_));
 sky130_fd_sc_hd__a31o_4 _8153_ (.A1(\arbiter.slave_sel[2][1] ),
    .A2(_3436_),
    .A3(_3437_),
    .B1(_3438_),
    .X(_3439_));
 sky130_fd_sc_hd__a21oi_1 _8154_ (.A1(_3439_),
    .A2(_3086_),
    .B1(_3071_),
    .Y(_3440_));
 sky130_fd_sc_hd__a22o_2 _8155_ (.A1(_3273_),
    .A2(_3423_),
    .B1(_3435_),
    .B2(_3440_),
    .X(net420));
 sky130_fd_sc_hd__o22a_1 _8156_ (.A1(net262),
    .A2(_0486_),
    .B1(net360),
    .B2(_0654_),
    .X(_3441_));
 sky130_fd_sc_hd__o221a_4 _8157_ (.A1(net285),
    .A2(_0888_),
    .B1(net323),
    .B2(_0197_),
    .C1(_3441_),
    .X(_3442_));
 sky130_fd_sc_hd__inv_2 _8158_ (.A(net360),
    .Y(_3443_));
 sky130_fd_sc_hd__nor2_1 _8159_ (.A(_4127_),
    .B(_3443_),
    .Y(_3444_));
 sky130_fd_sc_hd__nand2_1 _8160_ (.A(_4127_),
    .B(net262),
    .Y(_3445_));
 sky130_fd_sc_hd__nand2_1 _8161_ (.A(_3445_),
    .B(_4118_),
    .Y(_3446_));
 sky130_fd_sc_hd__inv_2 _8162_ (.A(net323),
    .Y(_3447_));
 sky130_fd_sc_hd__nand2_1 _8163_ (.A(_1989_),
    .B(_3447_),
    .Y(_3448_));
 sky130_fd_sc_hd__o221ai_2 _8164_ (.A1(net285),
    .A2(_0520_),
    .B1(_3444_),
    .B2(_3446_),
    .C1(_3448_),
    .Y(_3449_));
 sky130_fd_sc_hd__inv_2 _8165_ (.A(_3449_),
    .Y(_3450_));
 sky130_fd_sc_hd__nor2_1 _8166_ (.A(_4252_),
    .B(_3443_),
    .Y(_3451_));
 sky130_fd_sc_hd__a211o_1 _8167_ (.A1(_0510_),
    .A2(net262),
    .B1(_4245_),
    .C1(_3451_),
    .X(_3452_));
 sky130_fd_sc_hd__o221ai_2 _8168_ (.A1(net285),
    .A2(_4272_),
    .B1(net323),
    .B2(_4271_),
    .C1(_3452_),
    .Y(_3453_));
 sky130_fd_sc_hd__inv_2 _8169_ (.A(_3453_),
    .Y(_3454_));
 sky130_fd_sc_hd__a221o_1 _8170_ (.A1(_3080_),
    .A2(_3450_),
    .B1(_3454_),
    .B2(_3134_),
    .C1(_3085_),
    .X(_3455_));
 sky130_fd_sc_hd__nor2_1 _8171_ (.A(_0088_),
    .B(_3443_),
    .Y(_3456_));
 sky130_fd_sc_hd__nand2_1 _8172_ (.A(_0088_),
    .B(net262),
    .Y(_3457_));
 sky130_fd_sc_hd__nand2_1 _8173_ (.A(_3457_),
    .B(\arbiter.slave_sel[2][1] ),
    .Y(_3458_));
 sky130_fd_sc_hd__nand2_1 _8174_ (.A(_0143_),
    .B(_3447_),
    .Y(_3459_));
 sky130_fd_sc_hd__o221ai_4 _8175_ (.A1(net285),
    .A2(_0152_),
    .B1(_3456_),
    .B2(_3458_),
    .C1(_3459_),
    .Y(_3460_));
 sky130_fd_sc_hd__a21oi_1 _8176_ (.A1(_3460_),
    .A2(_3086_),
    .B1(_3071_),
    .Y(_3461_));
 sky130_fd_sc_hd__a22o_2 _8177_ (.A1(_3273_),
    .A2(_3442_),
    .B1(_3455_),
    .B2(_3461_),
    .X(net421));
 sky130_fd_sc_hd__nand2_1 _8178_ (.A(net264),
    .B(_0088_),
    .Y(_3462_));
 sky130_fd_sc_hd__inv_2 _8179_ (.A(_3462_),
    .Y(_3463_));
 sky130_fd_sc_hd__inv_2 _8180_ (.A(net361),
    .Y(_3464_));
 sky130_fd_sc_hd__nor2_1 _8181_ (.A(_0088_),
    .B(_3464_),
    .Y(_3465_));
 sky130_fd_sc_hd__o21a_1 _8182_ (.A1(_3463_),
    .A2(_3465_),
    .B1(\arbiter.slave_sel[2][1] ),
    .X(_3466_));
 sky130_fd_sc_hd__a221oi_4 _8183_ (.A1(net286),
    .A2(_0759_),
    .B1(net324),
    .B2(_0143_),
    .C1(_3466_),
    .Y(_3467_));
 sky130_fd_sc_hd__a21o_1 _8184_ (.A1(_3467_),
    .A2(_3085_),
    .B1(_3071_),
    .X(_3468_));
 sky130_fd_sc_hd__nand2_1 _8185_ (.A(_4115_),
    .B(_4118_),
    .Y(_3469_));
 sky130_fd_sc_hd__a21o_1 _8186_ (.A1(_0523_),
    .A2(net264),
    .B1(_3469_),
    .X(_3470_));
 sky130_fd_sc_hd__o221a_4 _8187_ (.A1(net286),
    .A2(_0520_),
    .B1(net324),
    .B2(_1971_),
    .C1(_3470_),
    .X(_3471_));
 sky130_fd_sc_hd__mux2_1 _8188_ (.A0(net361),
    .A1(net264),
    .S(_0558_),
    .X(_3472_));
 sky130_fd_sc_hd__and3_1 _8189_ (.A(_0555_),
    .B(_4245_),
    .C(net286),
    .X(_3473_));
 sky130_fd_sc_hd__a221o_4 _8190_ (.A1(net324),
    .A2(_1977_),
    .B1(_3472_),
    .B2(\arbiter.slave_sel[1][1] ),
    .C1(_3473_),
    .X(_3474_));
 sky130_fd_sc_hd__a221oi_1 _8191_ (.A1(_3471_),
    .A2(_3080_),
    .B1(_3474_),
    .B2(_3084_),
    .C1(_3086_),
    .Y(_3475_));
 sky130_fd_sc_hd__nand2_1 _8192_ (.A(net264),
    .B(_0198_),
    .Y(_3476_));
 sky130_fd_sc_hd__inv_2 _8193_ (.A(_3476_),
    .Y(_3477_));
 sky130_fd_sc_hd__nor2_1 _8194_ (.A(_0198_),
    .B(_3464_),
    .Y(_3478_));
 sky130_fd_sc_hd__o21a_1 _8195_ (.A1(_3477_),
    .A2(_3478_),
    .B1(\arbiter.slave_sel[3][1] ),
    .X(_3479_));
 sky130_fd_sc_hd__a221o_4 _8196_ (.A1(net286),
    .A2(_2439_),
    .B1(net324),
    .B2(_0652_),
    .C1(_3479_),
    .X(_3480_));
 sky130_fd_sc_hd__a2bb2o_2 _8197_ (.A1_N(_3468_),
    .A2_N(_3475_),
    .B1(_3072_),
    .B2(_3480_),
    .X(net422));
 sky130_fd_sc_hd__and2_1 _8198_ (.A(_0195_),
    .B(net362),
    .X(_3481_));
 sky130_fd_sc_hd__a211o_1 _8199_ (.A1(_0198_),
    .A2(net265),
    .B1(_0199_),
    .C1(_3481_),
    .X(_3482_));
 sky130_fd_sc_hd__o221a_2 _8200_ (.A1(net287),
    .A2(_0888_),
    .B1(net325),
    .B2(_0197_),
    .C1(_3482_),
    .X(_3483_));
 sky130_fd_sc_hd__a21o_1 _8201_ (.A1(_0799_),
    .A2(net362),
    .B1(_4119_),
    .X(_3484_));
 sky130_fd_sc_hd__a21o_1 _8202_ (.A1(_0522_),
    .A2(net265),
    .B1(_3484_),
    .X(_3485_));
 sky130_fd_sc_hd__o221a_2 _8203_ (.A1(net287),
    .A2(_0520_),
    .B1(net325),
    .B2(_1971_),
    .C1(_3485_),
    .X(_3486_));
 sky130_fd_sc_hd__a21o_1 _8204_ (.A1(_4253_),
    .A2(net362),
    .B1(_4245_),
    .X(_3487_));
 sky130_fd_sc_hd__a21o_1 _8205_ (.A1(_0510_),
    .A2(net265),
    .B1(_3487_),
    .X(_3488_));
 sky130_fd_sc_hd__o221a_2 _8206_ (.A1(net287),
    .A2(_0785_),
    .B1(net325),
    .B2(_4271_),
    .C1(_3488_),
    .X(_3489_));
 sky130_fd_sc_hd__a221o_1 _8207_ (.A1(_3486_),
    .A2(_3254_),
    .B1(_3489_),
    .B2(_3134_),
    .C1(_3085_),
    .X(_3490_));
 sky130_fd_sc_hd__a21o_1 _8208_ (.A1(_0090_),
    .A2(net362),
    .B1(_0096_),
    .X(_3491_));
 sky130_fd_sc_hd__a21o_1 _8209_ (.A1(_0088_),
    .A2(net265),
    .B1(_3491_),
    .X(_3492_));
 sky130_fd_sc_hd__o221a_2 _8210_ (.A1(net287),
    .A2(_0152_),
    .B1(net325),
    .B2(_0110_),
    .C1(_3492_),
    .X(_3493_));
 sky130_fd_sc_hd__inv_2 _8211_ (.A(_3493_),
    .Y(_3494_));
 sky130_fd_sc_hd__a21oi_1 _8212_ (.A1(_3494_),
    .A2(_3086_),
    .B1(_3071_),
    .Y(_3495_));
 sky130_fd_sc_hd__a22o_2 _8213_ (.A1(_3273_),
    .A2(_3483_),
    .B1(_3490_),
    .B2(_3495_),
    .X(net423));
 sky130_fd_sc_hd__a22o_1 _8214_ (.A1(_2439_),
    .A2(net289),
    .B1(_0651_),
    .B2(net326),
    .X(_3496_));
 sky130_fd_sc_hd__a221o_4 _8215_ (.A1(net363),
    .A2(_0766_),
    .B1(net266),
    .B2(_0194_),
    .C1(_3496_),
    .X(_3497_));
 sky130_fd_sc_hd__a22o_1 _8216_ (.A1(_0539_),
    .A2(net289),
    .B1(_1989_),
    .B2(net326),
    .X(_3498_));
 sky130_fd_sc_hd__a221o_4 _8217_ (.A1(net363),
    .A2(_0694_),
    .B1(net266),
    .B2(_0590_),
    .C1(_3498_),
    .X(_3499_));
 sky130_fd_sc_hd__a22o_1 _8218_ (.A1(_4268_),
    .A2(net266),
    .B1(net363),
    .B2(_0613_),
    .X(_3500_));
 sky130_fd_sc_hd__a221o_4 _8219_ (.A1(net326),
    .A2(_1977_),
    .B1(net289),
    .B2(_3081_),
    .C1(_3500_),
    .X(_3501_));
 sky130_fd_sc_hd__a221o_1 _8220_ (.A1(_3499_),
    .A2(_3079_),
    .B1(_3501_),
    .B2(_3134_),
    .C1(_3085_),
    .X(_3502_));
 sky130_fd_sc_hd__a22o_1 _8221_ (.A1(_0759_),
    .A2(net289),
    .B1(_0143_),
    .B2(net326),
    .X(_3503_));
 sky130_fd_sc_hd__a221o_4 _8222_ (.A1(net363),
    .A2(_0729_),
    .B1(net266),
    .B2(_0108_),
    .C1(_3503_),
    .X(_3504_));
 sky130_fd_sc_hd__o21ba_1 _8223_ (.A1(_3088_),
    .A2(_3504_),
    .B1_N(_3070_),
    .X(_3505_));
 sky130_fd_sc_hd__a22o_2 _8224_ (.A1(_3273_),
    .A2(_3497_),
    .B1(_3502_),
    .B2(_3505_),
    .X(net425));
 sky130_fd_sc_hd__a22o_1 _8225_ (.A1(_2439_),
    .A2(net290),
    .B1(_0652_),
    .B2(net327),
    .X(_3506_));
 sky130_fd_sc_hd__a221o_4 _8226_ (.A1(net364),
    .A2(_0767_),
    .B1(net267),
    .B2(_0194_),
    .C1(_3506_),
    .X(_3507_));
 sky130_fd_sc_hd__a22o_1 _8227_ (.A1(_4268_),
    .A2(net267),
    .B1(net364),
    .B2(_0612_),
    .X(_3508_));
 sky130_fd_sc_hd__a22o_1 _8228_ (.A1(_4280_),
    .A2(net327),
    .B1(net290),
    .B2(_4278_),
    .X(_3509_));
 sky130_fd_sc_hd__nor2_2 _8229_ (.A(_3508_),
    .B(_3509_),
    .Y(_3510_));
 sky130_fd_sc_hd__inv_2 _8230_ (.A(_3510_),
    .Y(_3511_));
 sky130_fd_sc_hd__a22o_1 _8231_ (.A1(_0539_),
    .A2(net290),
    .B1(_1989_),
    .B2(net327),
    .X(_3512_));
 sky130_fd_sc_hd__a221o_4 _8232_ (.A1(net364),
    .A2(_0694_),
    .B1(net267),
    .B2(_0590_),
    .C1(_3512_),
    .X(_3513_));
 sky130_fd_sc_hd__a221o_1 _8233_ (.A1(_3084_),
    .A2(_3511_),
    .B1(_3513_),
    .B2(_3080_),
    .C1(_3085_),
    .X(_3514_));
 sky130_fd_sc_hd__a22o_1 _8234_ (.A1(_3180_),
    .A2(net290),
    .B1(_3181_),
    .B2(net327),
    .X(_3515_));
 sky130_fd_sc_hd__a221oi_4 _8235_ (.A1(net364),
    .A2(_0572_),
    .B1(net267),
    .B2(_0108_),
    .C1(_3515_),
    .Y(_3516_));
 sky130_fd_sc_hd__a21oi_1 _8236_ (.A1(_3516_),
    .A2(_3086_),
    .B1(_3071_),
    .Y(_3517_));
 sky130_fd_sc_hd__a22o_2 _8237_ (.A1(_3071_),
    .A2(_3507_),
    .B1(_3514_),
    .B2(_3517_),
    .X(net426));
 sky130_fd_sc_hd__a21oi_1 _8238_ (.A1(_0118_),
    .A2(_3086_),
    .B1(_3071_),
    .Y(_3518_));
 sky130_fd_sc_hd__inv_2 _8239_ (.A(_4145_),
    .Y(_3519_));
 sky130_fd_sc_hd__inv_2 _8240_ (.A(_4286_),
    .Y(_3520_));
 sky130_fd_sc_hd__a221o_1 _8241_ (.A1(_3519_),
    .A2(_3079_),
    .B1(_3520_),
    .B2(_3078_),
    .C1(_3085_),
    .X(_3521_));
 sky130_fd_sc_hd__a22o_2 _8242_ (.A1(_3518_),
    .A2(_3521_),
    .B1(_0206_),
    .B2(_3072_),
    .X(net427));
 sky130_fd_sc_hd__a22o_1 _8243_ (.A1(_2439_),
    .A2(net292),
    .B1(_0767_),
    .B2(net232),
    .X(_3522_));
 sky130_fd_sc_hd__a221o_4 _8244_ (.A1(net329),
    .A2(_0652_),
    .B1(net269),
    .B2(_0194_),
    .C1(_3522_),
    .X(_3523_));
 sky130_fd_sc_hd__a22o_1 _8245_ (.A1(_4268_),
    .A2(net269),
    .B1(_4280_),
    .B2(net329),
    .X(_3524_));
 sky130_fd_sc_hd__a221oi_4 _8246_ (.A1(net292),
    .A2(_3081_),
    .B1(net232),
    .B2(_0613_),
    .C1(_3524_),
    .Y(_3525_));
 sky130_fd_sc_hd__inv_2 _8247_ (.A(_3525_),
    .Y(_3526_));
 sky130_fd_sc_hd__a22o_1 _8248_ (.A1(_0539_),
    .A2(net292),
    .B1(_0694_),
    .B2(net232),
    .X(_3527_));
 sky130_fd_sc_hd__a221o_4 _8249_ (.A1(net329),
    .A2(_1989_),
    .B1(net269),
    .B2(_0590_),
    .C1(_3527_),
    .X(_3528_));
 sky130_fd_sc_hd__a221o_1 _8250_ (.A1(_3526_),
    .A2(_3078_),
    .B1(_3528_),
    .B2(_3080_),
    .C1(_3085_),
    .X(_3529_));
 sky130_fd_sc_hd__a22o_1 _8251_ (.A1(_3180_),
    .A2(net292),
    .B1(_3181_),
    .B2(net329),
    .X(_3530_));
 sky130_fd_sc_hd__a221o_4 _8252_ (.A1(net232),
    .A2(_0572_),
    .B1(net269),
    .B2(_0108_),
    .C1(_3530_),
    .X(_3531_));
 sky130_fd_sc_hd__o21ba_1 _8253_ (.A1(_3088_),
    .A2(_3531_),
    .B1_N(_3070_),
    .X(_3532_));
 sky130_fd_sc_hd__a22o_2 _8254_ (.A1(_3071_),
    .A2(_3523_),
    .B1(_3529_),
    .B2(_3532_),
    .X(net428));
 sky130_fd_sc_hd__a22o_1 _8255_ (.A1(_0121_),
    .A2(_3504_),
    .B1(_3092_),
    .B2(_0126_),
    .X(_3533_));
 sky130_fd_sc_hd__nand2_2 _8256_ (.A(_0298_),
    .B(_4233_),
    .Y(_3534_));
 sky130_fd_sc_hd__and3_2 _8257_ (.A(_3534_),
    .B(_0588_),
    .C(_0664_),
    .X(_3535_));
 sky130_fd_sc_hd__buf_6 _8258_ (.A(_3535_),
    .X(_3536_));
 sky130_fd_sc_hd__inv_6 _8259_ (.A(_3534_),
    .Y(_3537_));
 sky130_fd_sc_hd__a22o_1 _8260_ (.A1(_3077_),
    .A2(_3536_),
    .B1(_3083_),
    .B2(_3537_),
    .X(_3538_));
 sky130_fd_sc_hd__nand2_8 _8261_ (.A(_0126_),
    .B(_4239_),
    .Y(_3539_));
 sky130_fd_sc_hd__mux2_1 _8262_ (.A0(_3533_),
    .A1(_3538_),
    .S(_3539_),
    .X(_3540_));
 sky130_fd_sc_hd__a22o_1 _8263_ (.A1(_0188_),
    .A2(_3497_),
    .B1(_3075_),
    .B2(_0184_),
    .X(_3541_));
 sky130_fd_sc_hd__nand2_8 _8264_ (.A(_0184_),
    .B(_0209_),
    .Y(_3542_));
 sky130_fd_sc_hd__inv_6 _8265_ (.A(_3542_),
    .Y(_3543_));
 sky130_fd_sc_hd__mux2_1 _8266_ (.A0(_3540_),
    .A1(_3541_),
    .S(_3543_),
    .X(_3544_));
 sky130_fd_sc_hd__buf_1 _8267_ (.A(_3544_),
    .X(net429));
 sky130_fd_sc_hd__inv_2 _8268_ (.A(_3539_),
    .Y(_3545_));
 sky130_fd_sc_hd__buf_6 _8269_ (.A(_3545_),
    .X(_3546_));
 sky130_fd_sc_hd__clkbuf_8 _8270_ (.A(_3546_),
    .X(_3547_));
 sky130_fd_sc_hd__nand2_4 _8271_ (.A(_0637_),
    .B(_0454_),
    .Y(_3548_));
 sky130_fd_sc_hd__nand2_1 _8272_ (.A(_3102_),
    .B(_0119_),
    .Y(_3549_));
 sky130_fd_sc_hd__o22a_1 _8273_ (.A1(_0457_),
    .A2(_3516_),
    .B1(_3548_),
    .B2(_3549_),
    .X(_3550_));
 sky130_fd_sc_hd__a21o_1 _8274_ (.A1(_0319_),
    .A2(_3511_),
    .B1(_3099_),
    .X(_3551_));
 sky130_fd_sc_hd__a22o_1 _8275_ (.A1(_3097_),
    .A2(_0664_),
    .B1(_0436_),
    .B2(_3513_),
    .X(_3552_));
 sky130_fd_sc_hd__a221oi_1 _8276_ (.A1(_3537_),
    .A2(_3551_),
    .B1(_3552_),
    .B2(_3536_),
    .C1(_3546_),
    .Y(_3553_));
 sky130_fd_sc_hd__a21oi_1 _8277_ (.A1(_3547_),
    .A2(_3550_),
    .B1(_3553_),
    .Y(_3554_));
 sky130_fd_sc_hd__mux2_1 _8278_ (.A0(_3554_),
    .A1(_3095_),
    .S(_3543_),
    .X(_3555_));
 sky130_fd_sc_hd__buf_1 _8279_ (.A(_3555_),
    .X(net430));
 sky130_fd_sc_hd__a221o_1 _8280_ (.A1(_3108_),
    .A2(_3535_),
    .B1(_3110_),
    .B2(_3537_),
    .C1(_3545_),
    .X(_3556_));
 sky130_fd_sc_hd__a21boi_1 _8281_ (.A1(_3113_),
    .A2(_3546_),
    .B1_N(_3556_),
    .Y(_3557_));
 sky130_fd_sc_hd__mux2_1 _8282_ (.A0(_3557_),
    .A1(_3106_),
    .S(_3543_),
    .X(_3558_));
 sky130_fd_sc_hd__buf_1 _8283_ (.A(_3558_),
    .X(net431));
 sky130_fd_sc_hd__nor2_1 _8284_ (.A(_0127_),
    .B(_3123_),
    .Y(_3559_));
 sky130_fd_sc_hd__a221o_1 _8285_ (.A1(_3118_),
    .A2(_3536_),
    .B1(_3120_),
    .B2(_3537_),
    .C1(_3546_),
    .X(_3560_));
 sky130_fd_sc_hd__o21a_1 _8286_ (.A1(_3539_),
    .A2(_3559_),
    .B1(_3560_),
    .X(_3561_));
 sky130_fd_sc_hd__mux2_1 _8287_ (.A0(_3561_),
    .A1(_3116_),
    .S(_3543_),
    .X(_3562_));
 sky130_fd_sc_hd__buf_1 _8288_ (.A(_3562_),
    .X(net432));
 sky130_fd_sc_hd__clkbuf_8 _8289_ (.A(_3542_),
    .X(_3563_));
 sky130_fd_sc_hd__nand2_8 _8290_ (.A(_0646_),
    .B(_0475_),
    .Y(_3564_));
 sky130_fd_sc_hd__clkinv_4 _8291_ (.A(_3564_),
    .Y(_3565_));
 sky130_fd_sc_hd__a21o_1 _8292_ (.A1(_3075_),
    .A2(\arbiter.master_sel[3][0] ),
    .B1(_3565_),
    .X(_3566_));
 sky130_fd_sc_hd__o221a_2 _8293_ (.A1(_0473_),
    .A2(_3129_),
    .B1(_0480_),
    .B2(_3106_),
    .C1(_3566_),
    .X(_3567_));
 sky130_fd_sc_hd__clkbuf_8 _8294_ (.A(_3539_),
    .X(_3568_));
 sky130_fd_sc_hd__nand2_1 _8295_ (.A(_3092_),
    .B(_0119_),
    .Y(_3569_));
 sky130_fd_sc_hd__a22o_1 _8296_ (.A1(_0121_),
    .A2(_3113_),
    .B1(_3145_),
    .B2(_0126_),
    .X(_3570_));
 sky130_fd_sc_hd__a21o_2 _8297_ (.A1(_3569_),
    .A2(_3548_),
    .B1(_3570_),
    .X(_3571_));
 sky130_fd_sc_hd__o21ai_1 _8298_ (.A1(_3568_),
    .A2(_3571_),
    .B1(_3563_),
    .Y(_3572_));
 sky130_fd_sc_hd__clkbuf_8 _8299_ (.A(_3537_),
    .X(_3573_));
 sky130_fd_sc_hd__nand2_4 _8300_ (.A(_0426_),
    .B(_0262_),
    .Y(_3574_));
 sky130_fd_sc_hd__inv_2 _8301_ (.A(_3574_),
    .Y(_3575_));
 sky130_fd_sc_hd__a21o_1 _8302_ (.A1(_3077_),
    .A2(\arbiter.master_sel[0][0] ),
    .B1(_3575_),
    .X(_3576_));
 sky130_fd_sc_hd__o221a_2 _8303_ (.A1(_0431_),
    .A2(_3140_),
    .B1(_0253_),
    .B2(_3108_),
    .C1(_3576_),
    .X(_3577_));
 sky130_fd_sc_hd__clkbuf_8 _8304_ (.A(_3536_),
    .X(_3578_));
 sky130_fd_sc_hd__a22o_1 _8305_ (.A1(_3133_),
    .A2(_3573_),
    .B1(_3577_),
    .B2(_3578_),
    .X(_3579_));
 sky130_fd_sc_hd__and2_1 _8306_ (.A(_3579_),
    .B(_3568_),
    .X(_3580_));
 sky130_fd_sc_hd__o22a_2 _8307_ (.A1(_3563_),
    .A2(_3567_),
    .B1(_3572_),
    .B2(_3580_),
    .X(net433));
 sky130_fd_sc_hd__a21o_1 _8308_ (.A1(_3097_),
    .A2(\arbiter.master_sel[0][0] ),
    .B1(_3575_),
    .X(_3581_));
 sky130_fd_sc_hd__o221a_2 _8309_ (.A1(_0431_),
    .A2(_3158_),
    .B1(_0253_),
    .B2(_3118_),
    .C1(_3581_),
    .X(_3582_));
 sky130_fd_sc_hd__nand2_2 _8310_ (.A(_0615_),
    .B(_0412_),
    .Y(_3583_));
 sky130_fd_sc_hd__inv_2 _8311_ (.A(_3583_),
    .Y(_3584_));
 sky130_fd_sc_hd__a21o_1 _8312_ (.A1(_3099_),
    .A2(\arbiter.master_sel[1][0] ),
    .B1(_3584_),
    .X(_3585_));
 sky130_fd_sc_hd__o221a_2 _8313_ (.A1(_0410_),
    .A2(_3163_),
    .B1(_0414_),
    .B2(_3120_),
    .C1(_3585_),
    .X(_3586_));
 sky130_fd_sc_hd__a22o_1 _8314_ (.A1(_3582_),
    .A2(_3536_),
    .B1(_3586_),
    .B2(_3537_),
    .X(_3587_));
 sky130_fd_sc_hd__inv_2 _8315_ (.A(_3152_),
    .Y(_3588_));
 sky130_fd_sc_hd__nand2_1 _8316_ (.A(_3549_),
    .B(_3548_),
    .Y(_3589_));
 sky130_fd_sc_hd__o221a_2 _8317_ (.A1(_0453_),
    .A2(_3588_),
    .B1(_0119_),
    .B2(_3559_),
    .C1(_3589_),
    .X(_3590_));
 sky130_fd_sc_hd__mux2_1 _8318_ (.A0(_3587_),
    .A1(_3590_),
    .S(_3546_),
    .X(_3591_));
 sky130_fd_sc_hd__a21o_1 _8319_ (.A1(_3095_),
    .A2(\arbiter.master_sel[3][0] ),
    .B1(_3565_),
    .X(_3592_));
 sky130_fd_sc_hd__o221a_2 _8320_ (.A1(_0473_),
    .A2(_3169_),
    .B1(_0480_),
    .B2(_3116_),
    .C1(_3592_),
    .X(_3593_));
 sky130_fd_sc_hd__mux2_1 _8321_ (.A0(_3591_),
    .A1(_3593_),
    .S(_3543_),
    .X(_3594_));
 sky130_fd_sc_hd__buf_1 _8322_ (.A(_3594_),
    .X(net434));
 sky130_fd_sc_hd__clkbuf_8 _8323_ (.A(_3543_),
    .X(_3595_));
 sky130_fd_sc_hd__a221o_1 _8324_ (.A1(_3175_),
    .A2(_3578_),
    .B1(_3177_),
    .B2(_3573_),
    .C1(_3547_),
    .X(_3596_));
 sky130_fd_sc_hd__o21a_1 _8325_ (.A1(_3568_),
    .A2(_3184_),
    .B1(_3563_),
    .X(_3597_));
 sky130_fd_sc_hd__a22o_1 _8326_ (.A1(_3173_),
    .A2(_3595_),
    .B1(_3596_),
    .B2(_3597_),
    .X(net436));
 sky130_fd_sc_hd__a221o_1 _8327_ (.A1(_3193_),
    .A2(_3578_),
    .B1(_3195_),
    .B2(_3573_),
    .C1(_3547_),
    .X(_3598_));
 sky130_fd_sc_hd__a21oi_1 _8328_ (.A1(_3198_),
    .A2(_3547_),
    .B1(_3595_),
    .Y(_3599_));
 sky130_fd_sc_hd__a22o_1 _8329_ (.A1(_3191_),
    .A2(_3595_),
    .B1(_3598_),
    .B2(_3599_),
    .X(net437));
 sky130_fd_sc_hd__a221o_1 _8330_ (.A1(_3205_),
    .A2(_3578_),
    .B1(_3207_),
    .B2(_3573_),
    .C1(_3547_),
    .X(_3600_));
 sky130_fd_sc_hd__o21a_1 _8331_ (.A1(_3568_),
    .A2(_3210_),
    .B1(_3563_),
    .X(_3601_));
 sky130_fd_sc_hd__a22o_2 _8332_ (.A1(_3203_),
    .A2(_3595_),
    .B1(_3600_),
    .B2(_3601_),
    .X(net438));
 sky130_fd_sc_hd__inv_2 _8333_ (.A(_3198_),
    .Y(_3602_));
 sky130_fd_sc_hd__nand2_1 _8334_ (.A(_3602_),
    .B(_0450_),
    .Y(_3603_));
 sky130_fd_sc_hd__nand2_1 _8335_ (.A(_3222_),
    .B(_0450_),
    .Y(_3604_));
 sky130_fd_sc_hd__mux2_1 _8336_ (.A0(_3603_),
    .A1(_3604_),
    .S(_0119_),
    .X(_3605_));
 sky130_fd_sc_hd__inv_2 _8337_ (.A(_3605_),
    .Y(_3606_));
 sky130_fd_sc_hd__a221o_1 _8338_ (.A1(_3217_),
    .A2(_3536_),
    .B1(_3219_),
    .B2(_3537_),
    .C1(_3545_),
    .X(_3607_));
 sky130_fd_sc_hd__o21a_1 _8339_ (.A1(_3539_),
    .A2(_3606_),
    .B1(_3607_),
    .X(_3608_));
 sky130_fd_sc_hd__o21a_1 _8340_ (.A1(_0480_),
    .A2(_3191_),
    .B1(_3215_),
    .X(_3609_));
 sky130_fd_sc_hd__mux2_1 _8341_ (.A0(_3608_),
    .A1(_3609_),
    .S(_3543_),
    .X(_3610_));
 sky130_fd_sc_hd__buf_1 _8342_ (.A(_3610_),
    .X(net439));
 sky130_fd_sc_hd__a221o_1 _8343_ (.A1(_3229_),
    .A2(_3536_),
    .B1(_3231_),
    .B2(_3537_),
    .C1(_3546_),
    .X(_3611_));
 sky130_fd_sc_hd__o21ai_2 _8344_ (.A1(_3234_),
    .A2(_3568_),
    .B1(_3611_),
    .Y(_3612_));
 sky130_fd_sc_hd__nand2_1 _8345_ (.A(_3227_),
    .B(_0646_),
    .Y(_3613_));
 sky130_fd_sc_hd__nand2_1 _8346_ (.A(_3203_),
    .B(_0469_),
    .Y(_3614_));
 sky130_fd_sc_hd__mux2_1 _8347_ (.A0(_3613_),
    .A1(_3614_),
    .S(_0183_),
    .X(_3615_));
 sky130_fd_sc_hd__inv_2 _8348_ (.A(_3615_),
    .Y(_3616_));
 sky130_fd_sc_hd__nor2_1 _8349_ (.A(_3563_),
    .B(_3616_),
    .Y(_3617_));
 sky130_fd_sc_hd__a21oi_4 _8350_ (.A1(_3612_),
    .A2(_3563_),
    .B1(_3617_),
    .Y(net440));
 sky130_fd_sc_hd__nand2_1 _8351_ (.A(_3241_),
    .B(_0427_),
    .Y(_3618_));
 sky130_fd_sc_hd__nand2_1 _8352_ (.A(_3217_),
    .B(_0427_),
    .Y(_3619_));
 sky130_fd_sc_hd__mux2_1 _8353_ (.A0(_3618_),
    .A1(_3619_),
    .S(_4153_),
    .X(_3620_));
 sky130_fd_sc_hd__nand2_1 _8354_ (.A(_3620_),
    .B(_3575_),
    .Y(_3621_));
 sky130_fd_sc_hd__a221o_1 _8355_ (.A1(_3243_),
    .A2(_3573_),
    .B1(_3621_),
    .B2(_3578_),
    .C1(_3547_),
    .X(_3622_));
 sky130_fd_sc_hd__o21a_1 _8356_ (.A1(_3568_),
    .A2(_3246_),
    .B1(_3563_),
    .X(_3623_));
 sky130_fd_sc_hd__a22o_2 _8357_ (.A1(_3239_),
    .A2(_3595_),
    .B1(_3622_),
    .B2(_3623_),
    .X(net441));
 sky130_fd_sc_hd__nand2_1 _8358_ (.A(_3253_),
    .B(_0426_),
    .Y(_3624_));
 sky130_fd_sc_hd__nand2_1 _8359_ (.A(_3229_),
    .B(_0426_),
    .Y(_3625_));
 sky130_fd_sc_hd__mux2_1 _8360_ (.A0(_3624_),
    .A1(_3625_),
    .S(_4153_),
    .X(_3626_));
 sky130_fd_sc_hd__inv_2 _8361_ (.A(_3626_),
    .Y(_3627_));
 sky130_fd_sc_hd__a22o_2 _8362_ (.A1(_0433_),
    .A2(_3205_),
    .B1(_3627_),
    .B2(_3575_),
    .X(_3628_));
 sky130_fd_sc_hd__a22o_1 _8363_ (.A1(_3256_),
    .A2(_3537_),
    .B1(_3628_),
    .B2(_3536_),
    .X(_3629_));
 sky130_fd_sc_hd__inv_2 _8364_ (.A(_3548_),
    .Y(_3630_));
 sky130_fd_sc_hd__a21o_1 _8365_ (.A1(_3210_),
    .A2(_0119_),
    .B1(_3630_),
    .X(_3631_));
 sky130_fd_sc_hd__o221a_2 _8366_ (.A1(_0453_),
    .A2(_3259_),
    .B1(_0457_),
    .B2(_3234_),
    .C1(_3631_),
    .X(_3632_));
 sky130_fd_sc_hd__mux2_1 _8367_ (.A0(_3629_),
    .A1(_3632_),
    .S(_3546_),
    .X(_3633_));
 sky130_fd_sc_hd__inv_2 _8368_ (.A(_0475_),
    .Y(_3634_));
 sky130_fd_sc_hd__nand2_1 _8369_ (.A(_3251_),
    .B(_0646_),
    .Y(_3635_));
 sky130_fd_sc_hd__mux2_1 _8370_ (.A0(_3635_),
    .A1(_3613_),
    .S(_0183_),
    .X(_3636_));
 sky130_fd_sc_hd__inv_2 _8371_ (.A(_3636_),
    .Y(_3637_));
 sky130_fd_sc_hd__a22o_1 _8372_ (.A1(_3634_),
    .A2(_3203_),
    .B1(_3637_),
    .B2(_3565_),
    .X(_3638_));
 sky130_fd_sc_hd__mux2_1 _8373_ (.A0(_3633_),
    .A1(_3638_),
    .S(_3543_),
    .X(_3639_));
 sky130_fd_sc_hd__buf_1 _8374_ (.A(_3639_),
    .X(net442));
 sky130_fd_sc_hd__nand2_1 _8375_ (.A(_3264_),
    .B(_0469_),
    .Y(_3640_));
 sky130_fd_sc_hd__nand2_1 _8376_ (.A(_3239_),
    .B(_0469_),
    .Y(_3641_));
 sky130_fd_sc_hd__mux2_1 _8377_ (.A0(_3640_),
    .A1(_3641_),
    .S(_0183_),
    .X(_3642_));
 sky130_fd_sc_hd__inv_2 _8378_ (.A(_3642_),
    .Y(_3643_));
 sky130_fd_sc_hd__a22o_2 _8379_ (.A1(_3634_),
    .A2(_3215_),
    .B1(_3643_),
    .B2(_3565_),
    .X(_3644_));
 sky130_fd_sc_hd__o22a_1 _8380_ (.A1(_0453_),
    .A2(_3271_),
    .B1(_0457_),
    .B2(_3246_),
    .X(_3645_));
 sky130_fd_sc_hd__o21ai_2 _8381_ (.A1(_3630_),
    .A2(_3606_),
    .B1(_3645_),
    .Y(_3646_));
 sky130_fd_sc_hd__o21ai_1 _8382_ (.A1(_3568_),
    .A2(_3646_),
    .B1(_3563_),
    .Y(_3647_));
 sky130_fd_sc_hd__a21o_1 _8383_ (.A1(_3219_),
    .A2(\arbiter.master_sel[1][0] ),
    .B1(_3584_),
    .X(_3648_));
 sky130_fd_sc_hd__o221a_2 _8384_ (.A1(_0410_),
    .A2(_3268_),
    .B1(_0414_),
    .B2(_3243_),
    .C1(_3648_),
    .X(_3649_));
 sky130_fd_sc_hd__o21a_1 _8385_ (.A1(_0262_),
    .A2(_3217_),
    .B1(_0427_),
    .X(_3650_));
 sky130_fd_sc_hd__o221a_2 _8386_ (.A1(_0253_),
    .A2(_3241_),
    .B1(_0431_),
    .B2(_3266_),
    .C1(_3650_),
    .X(_3651_));
 sky130_fd_sc_hd__a22o_1 _8387_ (.A1(_3649_),
    .A2(_3573_),
    .B1(_3578_),
    .B2(_3651_),
    .X(_3652_));
 sky130_fd_sc_hd__and2_1 _8388_ (.A(_3652_),
    .B(_3568_),
    .X(_3653_));
 sky130_fd_sc_hd__o22a_2 _8389_ (.A1(_3563_),
    .A2(_3644_),
    .B1(_3647_),
    .B2(_3653_),
    .X(net443));
 sky130_fd_sc_hd__nand2_1 _8390_ (.A(_3277_),
    .B(_0469_),
    .Y(_3654_));
 sky130_fd_sc_hd__mux2_1 _8391_ (.A0(_3654_),
    .A1(_3635_),
    .S(_0183_),
    .X(_3655_));
 sky130_fd_sc_hd__inv_2 _8392_ (.A(_3655_),
    .Y(_3656_));
 sky130_fd_sc_hd__mux2_1 _8393_ (.A0(_3656_),
    .A1(_3616_),
    .S(_3564_),
    .X(_3657_));
 sky130_fd_sc_hd__nand2_1 _8394_ (.A(_3279_),
    .B(_0427_),
    .Y(_3658_));
 sky130_fd_sc_hd__mux2_1 _8395_ (.A0(_3658_),
    .A1(_3624_),
    .S(_4153_),
    .X(_3659_));
 sky130_fd_sc_hd__a2bb2o_1 _8396_ (.A1_N(_3574_),
    .A2_N(_3659_),
    .B1(_0433_),
    .B2(_3229_),
    .X(_3660_));
 sky130_fd_sc_hd__a221o_1 _8397_ (.A1(_3281_),
    .A2(_3573_),
    .B1(_3660_),
    .B2(_3578_),
    .C1(_3547_),
    .X(_3661_));
 sky130_fd_sc_hd__o21a_1 _8398_ (.A1(_3568_),
    .A2(_3284_),
    .B1(_3542_),
    .X(_3662_));
 sky130_fd_sc_hd__a22o_2 _8399_ (.A1(_3595_),
    .A2(_3657_),
    .B1(_3661_),
    .B2(_3662_),
    .X(net444));
 sky130_fd_sc_hd__nand2_1 _8400_ (.A(_3289_),
    .B(_0646_),
    .Y(_3663_));
 sky130_fd_sc_hd__mux2_1 _8401_ (.A0(_3663_),
    .A1(_3640_),
    .S(_0183_),
    .X(_3664_));
 sky130_fd_sc_hd__a2bb2o_1 _8402_ (.A1_N(_3564_),
    .A2_N(_3664_),
    .B1(_3634_),
    .B2(_3239_),
    .X(_3665_));
 sky130_fd_sc_hd__nand2_1 _8403_ (.A(_3291_),
    .B(_0427_),
    .Y(_3666_));
 sky130_fd_sc_hd__nand2_1 _8404_ (.A(_3266_),
    .B(_0427_),
    .Y(_3667_));
 sky130_fd_sc_hd__mux2_1 _8405_ (.A0(_3666_),
    .A1(_3667_),
    .S(_4153_),
    .X(_3668_));
 sky130_fd_sc_hd__inv_2 _8406_ (.A(_3668_),
    .Y(_3669_));
 sky130_fd_sc_hd__nand2_1 _8407_ (.A(_3669_),
    .B(_3575_),
    .Y(_3670_));
 sky130_fd_sc_hd__o21ai_2 _8408_ (.A1(_0262_),
    .A2(_3620_),
    .B1(_3670_),
    .Y(_3671_));
 sky130_fd_sc_hd__a221o_1 _8409_ (.A1(_3293_),
    .A2(_3573_),
    .B1(_3671_),
    .B2(_3578_),
    .C1(_3547_),
    .X(_3672_));
 sky130_fd_sc_hd__o21a_1 _8410_ (.A1(_3568_),
    .A2(_3296_),
    .B1(_3542_),
    .X(_3673_));
 sky130_fd_sc_hd__a22o_2 _8411_ (.A1(_3595_),
    .A2(_3665_),
    .B1(_3672_),
    .B2(_3673_),
    .X(net445));
 sky130_fd_sc_hd__nand2_1 _8412_ (.A(_3301_),
    .B(_0646_),
    .Y(_3674_));
 sky130_fd_sc_hd__mux2_1 _8413_ (.A0(_3674_),
    .A1(_3654_),
    .S(_0183_),
    .X(_3675_));
 sky130_fd_sc_hd__nand2_1 _8414_ (.A(_3637_),
    .B(_3634_),
    .Y(_3676_));
 sky130_fd_sc_hd__o21ai_1 _8415_ (.A1(_3564_),
    .A2(_3675_),
    .B1(_3676_),
    .Y(_3677_));
 sky130_fd_sc_hd__nand2_1 _8416_ (.A(_3303_),
    .B(_0427_),
    .Y(_3678_));
 sky130_fd_sc_hd__mux2_1 _8417_ (.A0(_3678_),
    .A1(_3658_),
    .S(_4153_),
    .X(_3679_));
 sky130_fd_sc_hd__inv_2 _8418_ (.A(_3679_),
    .Y(_3680_));
 sky130_fd_sc_hd__mux2_1 _8419_ (.A0(_3680_),
    .A1(_3627_),
    .S(_3574_),
    .X(_3681_));
 sky130_fd_sc_hd__a221o_1 _8420_ (.A1(_3305_),
    .A2(_3573_),
    .B1(_3681_),
    .B2(_3578_),
    .C1(_3547_),
    .X(_3682_));
 sky130_fd_sc_hd__o21a_1 _8421_ (.A1(_3568_),
    .A2(_3308_),
    .B1(_3542_),
    .X(_3683_));
 sky130_fd_sc_hd__a22o_2 _8422_ (.A1(_3595_),
    .A2(_3677_),
    .B1(_3682_),
    .B2(_3683_),
    .X(net447));
 sky130_fd_sc_hd__nand2_1 _8423_ (.A(_3317_),
    .B(_0615_),
    .Y(_3684_));
 sky130_fd_sc_hd__nand2_1 _8424_ (.A(_3293_),
    .B(_0615_),
    .Y(_3685_));
 sky130_fd_sc_hd__mux2_1 _8425_ (.A0(_3684_),
    .A1(_3685_),
    .S(_4288_),
    .X(_3686_));
 sky130_fd_sc_hd__inv_2 _8426_ (.A(_3686_),
    .Y(_3687_));
 sky130_fd_sc_hd__nand2_1 _8427_ (.A(_3315_),
    .B(_0426_),
    .Y(_3688_));
 sky130_fd_sc_hd__mux2_1 _8428_ (.A0(_3688_),
    .A1(_3666_),
    .S(_4153_),
    .X(_3689_));
 sky130_fd_sc_hd__inv_2 _8429_ (.A(_3535_),
    .Y(_3690_));
 sky130_fd_sc_hd__a21oi_1 _8430_ (.A1(_3689_),
    .A2(_3575_),
    .B1(_3690_),
    .Y(_3691_));
 sky130_fd_sc_hd__a41o_1 _8431_ (.A1(_3687_),
    .A2(_4233_),
    .A3(\arbiter.master_sel[1][0] ),
    .A4(_0037_),
    .B1(_3691_),
    .X(_3692_));
 sky130_fd_sc_hd__mux2_1 _8432_ (.A0(_3692_),
    .A1(_3320_),
    .S(_3546_),
    .X(_3693_));
 sky130_fd_sc_hd__nand2_1 _8433_ (.A(_3313_),
    .B(_0646_),
    .Y(_3694_));
 sky130_fd_sc_hd__mux2_1 _8434_ (.A0(_3694_),
    .A1(_3663_),
    .S(_0183_),
    .X(_3695_));
 sky130_fd_sc_hd__nand2_1 _8435_ (.A(_3643_),
    .B(_3634_),
    .Y(_3696_));
 sky130_fd_sc_hd__o21ai_2 _8436_ (.A1(_3564_),
    .A2(_3695_),
    .B1(_3696_),
    .Y(_3697_));
 sky130_fd_sc_hd__mux2_2 _8437_ (.A0(_3693_),
    .A1(_3697_),
    .S(_3543_),
    .X(_3698_));
 sky130_fd_sc_hd__buf_1 _8438_ (.A(_3698_),
    .X(net448));
 sky130_fd_sc_hd__nand2_1 _8439_ (.A(_3327_),
    .B(_0646_),
    .Y(_3699_));
 sky130_fd_sc_hd__mux2_1 _8440_ (.A0(_3699_),
    .A1(_3674_),
    .S(_0183_),
    .X(_3700_));
 sky130_fd_sc_hd__nand2_1 _8441_ (.A(_3656_),
    .B(_3634_),
    .Y(_3701_));
 sky130_fd_sc_hd__o21ai_1 _8442_ (.A1(_3564_),
    .A2(_3700_),
    .B1(_3701_),
    .Y(_3702_));
 sky130_fd_sc_hd__a21o_1 _8443_ (.A1(_3336_),
    .A2(_3547_),
    .B1(_3543_),
    .X(_3703_));
 sky130_fd_sc_hd__nor2_2 _8444_ (.A(_0663_),
    .B(_3329_),
    .Y(_3704_));
 sky130_fd_sc_hd__inv_2 _8445_ (.A(_3704_),
    .Y(_3705_));
 sky130_fd_sc_hd__mux2_1 _8446_ (.A0(_3705_),
    .A1(_3678_),
    .S(_4153_),
    .X(_3706_));
 sky130_fd_sc_hd__mux2_1 _8447_ (.A0(_3706_),
    .A1(_3659_),
    .S(_3574_),
    .X(_3707_));
 sky130_fd_sc_hd__o22a_1 _8448_ (.A1(_3332_),
    .A2(_3534_),
    .B1(_3690_),
    .B2(_3707_),
    .X(_3708_));
 sky130_fd_sc_hd__nor2_1 _8449_ (.A(_3547_),
    .B(_3708_),
    .Y(_3709_));
 sky130_fd_sc_hd__o22a_2 _8450_ (.A1(_3563_),
    .A2(_3702_),
    .B1(_3703_),
    .B2(_3709_),
    .X(net449));
 sky130_fd_sc_hd__nand2_1 _8451_ (.A(_3341_),
    .B(_0469_),
    .Y(_3710_));
 sky130_fd_sc_hd__mux2_1 _8452_ (.A0(_3710_),
    .A1(_3694_),
    .S(_0183_),
    .X(_3711_));
 sky130_fd_sc_hd__nand2_1 _8453_ (.A(_3711_),
    .B(_3565_),
    .Y(_3712_));
 sky130_fd_sc_hd__nand2_1 _8454_ (.A(_3664_),
    .B(_3564_),
    .Y(_3713_));
 sky130_fd_sc_hd__nand2_1 _8455_ (.A(_3343_),
    .B(_0426_),
    .Y(_3714_));
 sky130_fd_sc_hd__mux2_1 _8456_ (.A0(_3714_),
    .A1(_3688_),
    .S(_4153_),
    .X(_3715_));
 sky130_fd_sc_hd__nand2_1 _8457_ (.A(_3715_),
    .B(_3575_),
    .Y(_3716_));
 sky130_fd_sc_hd__nand2_1 _8458_ (.A(_3345_),
    .B(_0615_),
    .Y(_3717_));
 sky130_fd_sc_hd__mux2_1 _8459_ (.A0(_3717_),
    .A1(_3684_),
    .S(_4288_),
    .X(_3718_));
 sky130_fd_sc_hd__nand2_1 _8460_ (.A(_3718_),
    .B(_3584_),
    .Y(_3719_));
 sky130_fd_sc_hd__a221o_1 _8461_ (.A1(_3716_),
    .A2(_3536_),
    .B1(_3719_),
    .B2(_3537_),
    .C1(_3546_),
    .X(_3720_));
 sky130_fd_sc_hd__o211a_1 _8462_ (.A1(_3348_),
    .A2(_3539_),
    .B1(_3542_),
    .C1(_3720_),
    .X(_3721_));
 sky130_fd_sc_hd__a31o_2 _8463_ (.A1(_3595_),
    .A2(_3712_),
    .A3(_3713_),
    .B1(_3721_),
    .X(net450));
 sky130_fd_sc_hd__nand2_1 _8464_ (.A(_3355_),
    .B(_0427_),
    .Y(_3722_));
 sky130_fd_sc_hd__mux2_1 _8465_ (.A0(_3705_),
    .A1(_3722_),
    .S(\arbiter.master_sel[0][0] ),
    .X(_3723_));
 sky130_fd_sc_hd__nand2_1 _8466_ (.A(_3723_),
    .B(_3575_),
    .Y(_3724_));
 sky130_fd_sc_hd__o211a_1 _8467_ (.A1(_3575_),
    .A2(_3680_),
    .B1(_3536_),
    .C1(_3724_),
    .X(_3725_));
 sky130_fd_sc_hd__nand2_1 _8468_ (.A(_3333_),
    .B(_0615_),
    .Y(_3726_));
 sky130_fd_sc_hd__nand2_1 _8469_ (.A(_3357_),
    .B(_0615_),
    .Y(_3727_));
 sky130_fd_sc_hd__mux2_1 _8470_ (.A0(_3726_),
    .A1(_3727_),
    .S(\arbiter.master_sel[1][0] ),
    .X(_3728_));
 sky130_fd_sc_hd__inv_2 _8471_ (.A(_3728_),
    .Y(_3729_));
 sky130_fd_sc_hd__a41o_1 _8472_ (.A1(_3729_),
    .A2(_4233_),
    .A3(\arbiter.master_sel[1][0] ),
    .A4(_0037_),
    .B1(_3546_),
    .X(_3730_));
 sky130_fd_sc_hd__o22a_1 _8473_ (.A1(_3360_),
    .A2(_3539_),
    .B1(_3725_),
    .B2(_3730_),
    .X(_3731_));
 sky130_fd_sc_hd__mux2_2 _8474_ (.A0(_3731_),
    .A1(_3353_),
    .S(_3543_),
    .X(_3732_));
 sky130_fd_sc_hd__buf_1 _8475_ (.A(_3732_),
    .X(net451));
 sky130_fd_sc_hd__nand2_1 _8476_ (.A(_3365_),
    .B(_0469_),
    .Y(_3733_));
 sky130_fd_sc_hd__mux2_1 _8477_ (.A0(_3733_),
    .A1(_3710_),
    .S(_0183_),
    .X(_3734_));
 sky130_fd_sc_hd__mux2_1 _8478_ (.A0(_3734_),
    .A1(_3695_),
    .S(_3564_),
    .X(_3735_));
 sky130_fd_sc_hd__inv_2 _8479_ (.A(_3735_),
    .Y(_3736_));
 sky130_fd_sc_hd__nand2_1 _8480_ (.A(_3369_),
    .B(_0615_),
    .Y(_3737_));
 sky130_fd_sc_hd__mux2_1 _8481_ (.A0(_3737_),
    .A1(_3717_),
    .S(_4288_),
    .X(_3738_));
 sky130_fd_sc_hd__nand2_1 _8482_ (.A(_3738_),
    .B(_3584_),
    .Y(_3739_));
 sky130_fd_sc_hd__nand2_1 _8483_ (.A(_3367_),
    .B(_0427_),
    .Y(_3740_));
 sky130_fd_sc_hd__mux2_1 _8484_ (.A0(_3740_),
    .A1(_3714_),
    .S(_4153_),
    .X(_3741_));
 sky130_fd_sc_hd__mux2_1 _8485_ (.A0(_3741_),
    .A1(_3689_),
    .S(_3574_),
    .X(_3742_));
 sky130_fd_sc_hd__inv_2 _8486_ (.A(_3742_),
    .Y(_3743_));
 sky130_fd_sc_hd__a221o_1 _8487_ (.A1(_3573_),
    .A2(_3739_),
    .B1(_3743_),
    .B2(_3578_),
    .C1(_3547_),
    .X(_3744_));
 sky130_fd_sc_hd__o21a_1 _8488_ (.A1(_3568_),
    .A2(_3372_),
    .B1(_3542_),
    .X(_3745_));
 sky130_fd_sc_hd__a22o_2 _8489_ (.A1(_3595_),
    .A2(_3736_),
    .B1(_3744_),
    .B2(_3745_),
    .X(net452));
 sky130_fd_sc_hd__nand2_1 _8490_ (.A(_3377_),
    .B(_0646_),
    .Y(_3746_));
 sky130_fd_sc_hd__nand2_1 _8491_ (.A(_3353_),
    .B(_0646_),
    .Y(_3747_));
 sky130_fd_sc_hd__mux2_1 _8492_ (.A0(_3746_),
    .A1(_3747_),
    .S(_0183_),
    .X(_3748_));
 sky130_fd_sc_hd__mux2_1 _8493_ (.A0(_3700_),
    .A1(_3748_),
    .S(_3565_),
    .X(_3749_));
 sky130_fd_sc_hd__inv_2 _8494_ (.A(_3749_),
    .Y(_3750_));
 sky130_fd_sc_hd__a22o_1 _8495_ (.A1(_3379_),
    .A2(_3536_),
    .B1(_3381_),
    .B2(_3537_),
    .X(_3751_));
 sky130_fd_sc_hd__mux2_1 _8496_ (.A0(_3751_),
    .A1(net731),
    .S(_3546_),
    .X(_3752_));
 sky130_fd_sc_hd__mux2_2 _8497_ (.A0(_3750_),
    .A1(_3752_),
    .S(_3542_),
    .X(_3753_));
 sky130_fd_sc_hd__buf_1 _8498_ (.A(_3753_),
    .X(net453));
 sky130_fd_sc_hd__nand2_1 _8499_ (.A(_3389_),
    .B(_0469_),
    .Y(_3754_));
 sky130_fd_sc_hd__mux2_1 _8500_ (.A0(_3754_),
    .A1(_3733_),
    .S(_0183_),
    .X(_3755_));
 sky130_fd_sc_hd__mux2_1 _8501_ (.A0(_3755_),
    .A1(_3711_),
    .S(_3564_),
    .X(_3756_));
 sky130_fd_sc_hd__inv_2 _8502_ (.A(_3756_),
    .Y(_3757_));
 sky130_fd_sc_hd__nand2_1 _8503_ (.A(_3391_),
    .B(_0427_),
    .Y(_3758_));
 sky130_fd_sc_hd__mux2_1 _8504_ (.A0(_3758_),
    .A1(_3740_),
    .S(_4153_),
    .X(_3759_));
 sky130_fd_sc_hd__mux2_1 _8505_ (.A0(_3759_),
    .A1(_3715_),
    .S(_3574_),
    .X(_3760_));
 sky130_fd_sc_hd__inv_2 _8506_ (.A(_3760_),
    .Y(_3761_));
 sky130_fd_sc_hd__a221o_1 _8507_ (.A1(_3393_),
    .A2(_3573_),
    .B1(_3761_),
    .B2(_3578_),
    .C1(_3547_),
    .X(_3762_));
 sky130_fd_sc_hd__o21a_1 _8508_ (.A1(_3539_),
    .A2(_3396_),
    .B1(_3542_),
    .X(_3763_));
 sky130_fd_sc_hd__a22o_2 _8509_ (.A1(_3595_),
    .A2(_3757_),
    .B1(_3762_),
    .B2(_3763_),
    .X(net454));
 sky130_fd_sc_hd__nand2_1 _8510_ (.A(_3403_),
    .B(_0427_),
    .Y(_3764_));
 sky130_fd_sc_hd__nand2_1 _8511_ (.A(_3379_),
    .B(_0427_),
    .Y(_3765_));
 sky130_fd_sc_hd__mux2_1 _8512_ (.A0(_3764_),
    .A1(_3765_),
    .S(_4153_),
    .X(_3766_));
 sky130_fd_sc_hd__nand2_1 _8513_ (.A(_3766_),
    .B(_3575_),
    .Y(_3767_));
 sky130_fd_sc_hd__a221o_1 _8514_ (.A1(_3405_),
    .A2(_3573_),
    .B1(_3767_),
    .B2(_3578_),
    .C1(_3546_),
    .X(_3768_));
 sky130_fd_sc_hd__nand2_1 _8515_ (.A(_3408_),
    .B(_0451_),
    .Y(_3769_));
 sky130_fd_sc_hd__nand2_1 _8516_ (.A(net731),
    .B(_0451_),
    .Y(_3770_));
 sky130_fd_sc_hd__mux2_1 _8517_ (.A0(_3769_),
    .A1(_3770_),
    .S(_0125_),
    .X(_3771_));
 sky130_fd_sc_hd__nand2_1 _8518_ (.A(_3771_),
    .B(_3547_),
    .Y(_3772_));
 sky130_fd_sc_hd__nand2_1 _8519_ (.A(_3401_),
    .B(_0469_),
    .Y(_3773_));
 sky130_fd_sc_hd__mux2_1 _8520_ (.A0(_3773_),
    .A1(_3746_),
    .S(_0183_),
    .X(_3774_));
 sky130_fd_sc_hd__a21oi_1 _8521_ (.A1(_3774_),
    .A2(_3565_),
    .B1(_3563_),
    .Y(_3775_));
 sky130_fd_sc_hd__a31o_2 _8522_ (.A1(_3768_),
    .A2(_3563_),
    .A3(_3772_),
    .B1(_3775_),
    .X(net455));
 sky130_fd_sc_hd__nand2_1 _8523_ (.A(_3413_),
    .B(_0469_),
    .Y(_3776_));
 sky130_fd_sc_hd__mux2_2 _8524_ (.A0(_3776_),
    .A1(_3754_),
    .S(_0183_),
    .X(_3777_));
 sky130_fd_sc_hd__inv_2 _8525_ (.A(_3777_),
    .Y(_3778_));
 sky130_fd_sc_hd__a221o_1 _8526_ (.A1(_3415_),
    .A2(_3578_),
    .B1(_3417_),
    .B2(_3573_),
    .C1(_3546_),
    .X(_3779_));
 sky130_fd_sc_hd__o21a_1 _8527_ (.A1(_3539_),
    .A2(_3420_),
    .B1(_3542_),
    .X(_3780_));
 sky130_fd_sc_hd__a22o_2 _8528_ (.A1(_3595_),
    .A2(_3778_),
    .B1(_3779_),
    .B2(_3780_),
    .X(net456));
 sky130_fd_sc_hd__a221o_1 _8529_ (.A1(_3431_),
    .A2(_3578_),
    .B1(_3434_),
    .B2(_3573_),
    .C1(_3546_),
    .X(_3781_));
 sky130_fd_sc_hd__a21oi_1 _8530_ (.A1(_3439_),
    .A2(_3547_),
    .B1(_3543_),
    .Y(_3782_));
 sky130_fd_sc_hd__a22o_1 _8531_ (.A1(_3423_),
    .A2(_3595_),
    .B1(_3781_),
    .B2(_3782_),
    .X(net458));
 sky130_fd_sc_hd__a221o_1 _8532_ (.A1(_3450_),
    .A2(_3578_),
    .B1(_3454_),
    .B2(_3573_),
    .C1(_3546_),
    .X(_3783_));
 sky130_fd_sc_hd__a21oi_1 _8533_ (.A1(_3460_),
    .A2(_3547_),
    .B1(_3543_),
    .Y(_3784_));
 sky130_fd_sc_hd__a22o_2 _8534_ (.A1(_3442_),
    .A2(_3595_),
    .B1(_3783_),
    .B2(_3784_),
    .X(net459));
 sky130_fd_sc_hd__nand2_1 _8535_ (.A(_3774_),
    .B(_3564_),
    .Y(_3785_));
 sky130_fd_sc_hd__o221a_1 _8536_ (.A1(_0473_),
    .A2(_3480_),
    .B1(_0480_),
    .B2(_3423_),
    .C1(_3785_),
    .X(_3786_));
 sky130_fd_sc_hd__a22o_1 _8537_ (.A1(_0126_),
    .A2(_3467_),
    .B1(_3439_),
    .B2(_0121_),
    .X(_3787_));
 sky130_fd_sc_hd__a21o_1 _8538_ (.A1(_3771_),
    .A2(_3548_),
    .B1(_3787_),
    .X(_3788_));
 sky130_fd_sc_hd__o21ai_1 _8539_ (.A1(_3568_),
    .A2(_3788_),
    .B1(_3563_),
    .Y(_3789_));
 sky130_fd_sc_hd__nand2_1 _8540_ (.A(_3766_),
    .B(_3574_),
    .Y(_3790_));
 sky130_fd_sc_hd__o221a_2 _8541_ (.A1(_0253_),
    .A2(_3431_),
    .B1(_0431_),
    .B2(_3471_),
    .C1(_3790_),
    .X(_3791_));
 sky130_fd_sc_hd__a22o_1 _8542_ (.A1(_3474_),
    .A2(_3537_),
    .B1(_3791_),
    .B2(_3536_),
    .X(_3792_));
 sky130_fd_sc_hd__and2_1 _8543_ (.A(_3792_),
    .B(_3568_),
    .X(_3793_));
 sky130_fd_sc_hd__o22a_1 _8544_ (.A1(_3563_),
    .A2(_3786_),
    .B1(_3789_),
    .B2(_3793_),
    .X(net460));
 sky130_fd_sc_hd__a21oi_1 _8545_ (.A1(_3420_),
    .A2(_0119_),
    .B1(_3630_),
    .Y(_3794_));
 sky130_fd_sc_hd__a221o_1 _8546_ (.A1(_0121_),
    .A2(_3460_),
    .B1(_3494_),
    .B2(_0126_),
    .C1(_3794_),
    .X(_3795_));
 sky130_fd_sc_hd__inv_2 _8547_ (.A(_3795_),
    .Y(_3796_));
 sky130_fd_sc_hd__a21o_1 _8548_ (.A1(_3417_),
    .A2(\arbiter.master_sel[1][0] ),
    .B1(_3584_),
    .X(_3797_));
 sky130_fd_sc_hd__o221a_1 _8549_ (.A1(_0414_),
    .A2(_3454_),
    .B1(_0410_),
    .B2(_3489_),
    .C1(_3797_),
    .X(_3798_));
 sky130_fd_sc_hd__nand2_1 _8550_ (.A(_3415_),
    .B(_0427_),
    .Y(_3799_));
 sky130_fd_sc_hd__nand2_1 _8551_ (.A(_3799_),
    .B(_3574_),
    .Y(_3800_));
 sky130_fd_sc_hd__o221a_1 _8552_ (.A1(_0253_),
    .A2(_3450_),
    .B1(_0431_),
    .B2(_3486_),
    .C1(_3800_),
    .X(_3801_));
 sky130_fd_sc_hd__a221o_1 _8553_ (.A1(_3798_),
    .A2(_3537_),
    .B1(_3801_),
    .B2(_3536_),
    .C1(_3545_),
    .X(_3802_));
 sky130_fd_sc_hd__o21a_1 _8554_ (.A1(_3539_),
    .A2(_3796_),
    .B1(_3802_),
    .X(_3803_));
 sky130_fd_sc_hd__nand2_1 _8555_ (.A(_3777_),
    .B(_3564_),
    .Y(_3804_));
 sky130_fd_sc_hd__o221a_1 _8556_ (.A1(_0480_),
    .A2(_3442_),
    .B1(_0473_),
    .B2(_3483_),
    .C1(_3804_),
    .X(_3805_));
 sky130_fd_sc_hd__mux2_1 _8557_ (.A0(_3803_),
    .A1(_3805_),
    .S(_3543_),
    .X(_3806_));
 sky130_fd_sc_hd__buf_1 _8558_ (.A(_3806_),
    .X(net461));
 sky130_fd_sc_hd__a221o_1 _8559_ (.A1(_3499_),
    .A2(_3578_),
    .B1(_3501_),
    .B2(_3573_),
    .C1(_3546_),
    .X(_3807_));
 sky130_fd_sc_hd__o21a_1 _8560_ (.A1(_3539_),
    .A2(_3504_),
    .B1(_3542_),
    .X(_3808_));
 sky130_fd_sc_hd__a22o_1 _8561_ (.A1(_3497_),
    .A2(_3595_),
    .B1(_3807_),
    .B2(_3808_),
    .X(net462));
 sky130_fd_sc_hd__o21ai_1 _8562_ (.A1(_3568_),
    .A2(_3516_),
    .B1(_3563_),
    .Y(_3809_));
 sky130_fd_sc_hd__a22o_1 _8563_ (.A1(_3511_),
    .A2(_3537_),
    .B1(_3513_),
    .B2(_3536_),
    .X(_3810_));
 sky130_fd_sc_hd__and2_1 _8564_ (.A(_3810_),
    .B(_3568_),
    .X(_3811_));
 sky130_fd_sc_hd__o22a_1 _8565_ (.A1(_3507_),
    .A2(_3563_),
    .B1(_3809_),
    .B2(_3811_),
    .X(net463));
 sky130_fd_sc_hd__a22o_1 _8566_ (.A1(_3519_),
    .A2(_3536_),
    .B1(_3520_),
    .B2(_3537_),
    .X(_3812_));
 sky130_fd_sc_hd__nand2_1 _8567_ (.A(_3812_),
    .B(_3539_),
    .Y(_3813_));
 sky130_fd_sc_hd__o211a_1 _8568_ (.A1(_3539_),
    .A2(_0118_),
    .B1(_3542_),
    .C1(_3813_),
    .X(_3814_));
 sky130_fd_sc_hd__a21oi_2 _8569_ (.A1(_0205_),
    .A2(_3595_),
    .B1(_3814_),
    .Y(net464));
 sky130_fd_sc_hd__a221o_1 _8570_ (.A1(_3526_),
    .A2(_3537_),
    .B1(_3528_),
    .B2(_3536_),
    .C1(_3545_),
    .X(_3815_));
 sky130_fd_sc_hd__o21a_1 _8571_ (.A1(_3531_),
    .A2(_3539_),
    .B1(_3815_),
    .X(_3816_));
 sky130_fd_sc_hd__mux2_1 _8572_ (.A0(_3816_),
    .A1(_3523_),
    .S(_3543_),
    .X(_3817_));
 sky130_fd_sc_hd__buf_1 _8573_ (.A(_3817_),
    .X(net465));
 sky130_fd_sc_hd__nand2_2 _8574_ (.A(_0188_),
    .B(_0209_),
    .Y(_3818_));
 sky130_fd_sc_hd__inv_2 _8575_ (.A(_3818_),
    .Y(_3819_));
 sky130_fd_sc_hd__clkbuf_8 _8576_ (.A(_3819_),
    .X(_3820_));
 sky130_fd_sc_hd__buf_4 _8577_ (.A(_3820_),
    .X(_3821_));
 sky130_fd_sc_hd__nand2_4 _8578_ (.A(_0319_),
    .B(_4233_),
    .Y(_3822_));
 sky130_fd_sc_hd__and3_1 _8579_ (.A(_3822_),
    .B(_0588_),
    .C(_0436_),
    .X(_3823_));
 sky130_fd_sc_hd__clkbuf_8 _8580_ (.A(_3823_),
    .X(_3824_));
 sky130_fd_sc_hd__buf_4 _8581_ (.A(_3824_),
    .X(_3825_));
 sky130_fd_sc_hd__inv_6 _8582_ (.A(_3822_),
    .Y(_3826_));
 sky130_fd_sc_hd__buf_4 _8583_ (.A(_3826_),
    .X(_3827_));
 sky130_fd_sc_hd__nand2_2 _8584_ (.A(_0121_),
    .B(_4239_),
    .Y(_3828_));
 sky130_fd_sc_hd__clkinv_4 _8585_ (.A(_3828_),
    .Y(_3829_));
 sky130_fd_sc_hd__clkbuf_8 _8586_ (.A(_3829_),
    .X(_3830_));
 sky130_fd_sc_hd__buf_4 _8587_ (.A(_3830_),
    .X(_3831_));
 sky130_fd_sc_hd__a221o_1 _8588_ (.A1(_3077_),
    .A2(_3825_),
    .B1(_3083_),
    .B2(_3827_),
    .C1(_3831_),
    .X(_3832_));
 sky130_fd_sc_hd__clkbuf_8 _8589_ (.A(_3828_),
    .X(_3833_));
 sky130_fd_sc_hd__clkbuf_8 _8590_ (.A(_3818_),
    .X(_3834_));
 sky130_fd_sc_hd__o21a_1 _8591_ (.A1(_3833_),
    .A2(_3092_),
    .B1(_3834_),
    .X(_3835_));
 sky130_fd_sc_hd__a22o_1 _8592_ (.A1(_3075_),
    .A2(_3821_),
    .B1(_3832_),
    .B2(_3835_),
    .X(net466));
 sky130_fd_sc_hd__a22o_1 _8593_ (.A1(_3097_),
    .A2(_3824_),
    .B1(_3099_),
    .B2(_3826_),
    .X(_3836_));
 sky130_fd_sc_hd__mux2_1 _8594_ (.A0(_3836_),
    .A1(_3102_),
    .S(_3830_),
    .X(_3837_));
 sky130_fd_sc_hd__mux2_1 _8595_ (.A0(_3837_),
    .A1(_3095_),
    .S(_3820_),
    .X(_3838_));
 sky130_fd_sc_hd__buf_1 _8596_ (.A(_3838_),
    .X(net467));
 sky130_fd_sc_hd__a221o_1 _8597_ (.A1(_3110_),
    .A2(_3827_),
    .B1(_3577_),
    .B2(_3825_),
    .C1(_3831_),
    .X(_3839_));
 sky130_fd_sc_hd__a21oi_1 _8598_ (.A1(_3571_),
    .A2(_3831_),
    .B1(_3820_),
    .Y(_3840_));
 sky130_fd_sc_hd__a22o_1 _8599_ (.A1(_3567_),
    .A2(_3821_),
    .B1(_3839_),
    .B2(_3840_),
    .X(net469));
 sky130_fd_sc_hd__a221o_1 _8600_ (.A1(_3582_),
    .A2(_3825_),
    .B1(_3586_),
    .B2(_3827_),
    .C1(_3831_),
    .X(_3841_));
 sky130_fd_sc_hd__o21a_1 _8601_ (.A1(_3833_),
    .A2(_3590_),
    .B1(_3834_),
    .X(_3842_));
 sky130_fd_sc_hd__a22o_1 _8602_ (.A1(_3593_),
    .A2(_3821_),
    .B1(_3841_),
    .B2(_3842_),
    .X(net470));
 sky130_fd_sc_hd__a221o_1 _8603_ (.A1(_3133_),
    .A2(_3827_),
    .B1(_3140_),
    .B2(_3825_),
    .C1(_3831_),
    .X(_3843_));
 sky130_fd_sc_hd__a21oi_1 _8604_ (.A1(_3145_),
    .A2(_3831_),
    .B1(_3820_),
    .Y(_3844_));
 sky130_fd_sc_hd__a22o_1 _8605_ (.A1(_3129_),
    .A2(_3821_),
    .B1(_3843_),
    .B2(_3844_),
    .X(net471));
 sky130_fd_sc_hd__a221o_1 _8606_ (.A1(_3158_),
    .A2(_3824_),
    .B1(_3163_),
    .B2(_3826_),
    .C1(_3829_),
    .X(_3845_));
 sky130_fd_sc_hd__o21a_1 _8607_ (.A1(_3588_),
    .A2(_3828_),
    .B1(_3845_),
    .X(_3846_));
 sky130_fd_sc_hd__mux2_1 _8608_ (.A0(_3846_),
    .A1(_3169_),
    .S(_3820_),
    .X(_3847_));
 sky130_fd_sc_hd__buf_1 _8609_ (.A(_3847_),
    .X(net472));
 sky130_fd_sc_hd__a221o_1 _8610_ (.A1(_3175_),
    .A2(_3825_),
    .B1(_3177_),
    .B2(_3827_),
    .C1(_3831_),
    .X(_3848_));
 sky130_fd_sc_hd__o21a_1 _8611_ (.A1(_3833_),
    .A2(_3184_),
    .B1(_3834_),
    .X(_3849_));
 sky130_fd_sc_hd__a22o_1 _8612_ (.A1(_3173_),
    .A2(_3821_),
    .B1(_3848_),
    .B2(_3849_),
    .X(net473));
 sky130_fd_sc_hd__a22o_1 _8613_ (.A1(_3193_),
    .A2(_3824_),
    .B1(_3195_),
    .B2(_3826_),
    .X(_3850_));
 sky130_fd_sc_hd__mux2_1 _8614_ (.A0(_3850_),
    .A1(_3602_),
    .S(_3830_),
    .X(_3851_));
 sky130_fd_sc_hd__mux2_1 _8615_ (.A0(_3851_),
    .A1(_3191_),
    .S(_3820_),
    .X(_3852_));
 sky130_fd_sc_hd__buf_1 _8616_ (.A(_3852_),
    .X(net474));
 sky130_fd_sc_hd__a221o_1 _8617_ (.A1(_3205_),
    .A2(_3825_),
    .B1(_3207_),
    .B2(_3827_),
    .C1(_3831_),
    .X(_3853_));
 sky130_fd_sc_hd__o21a_1 _8618_ (.A1(_3833_),
    .A2(_3210_),
    .B1(_3834_),
    .X(_3854_));
 sky130_fd_sc_hd__a22o_1 _8619_ (.A1(_3203_),
    .A2(_3821_),
    .B1(_3853_),
    .B2(_3854_),
    .X(net475));
 sky130_fd_sc_hd__a22o_1 _8620_ (.A1(_3217_),
    .A2(_3824_),
    .B1(_3219_),
    .B2(_3826_),
    .X(_3855_));
 sky130_fd_sc_hd__mux2_1 _8621_ (.A0(_3855_),
    .A1(_3222_),
    .S(_3830_),
    .X(_3856_));
 sky130_fd_sc_hd__mux2_1 _8622_ (.A0(_3856_),
    .A1(_3215_),
    .S(_3820_),
    .X(_3857_));
 sky130_fd_sc_hd__buf_1 _8623_ (.A(_3857_),
    .X(net476));
 sky130_fd_sc_hd__a221o_1 _8624_ (.A1(_3231_),
    .A2(_3827_),
    .B1(_3628_),
    .B2(_3825_),
    .C1(_3831_),
    .X(_3858_));
 sky130_fd_sc_hd__o21a_1 _8625_ (.A1(_3833_),
    .A2(_3632_),
    .B1(_3834_),
    .X(_3859_));
 sky130_fd_sc_hd__a22o_1 _8626_ (.A1(_3638_),
    .A2(_3821_),
    .B1(_3858_),
    .B2(_3859_),
    .X(net477));
 sky130_fd_sc_hd__a221o_1 _8627_ (.A1(_3649_),
    .A2(_3826_),
    .B1(_3651_),
    .B2(_3825_),
    .C1(_3831_),
    .X(_3860_));
 sky130_fd_sc_hd__a21oi_1 _8628_ (.A1(_3646_),
    .A2(_3831_),
    .B1(_3820_),
    .Y(_3861_));
 sky130_fd_sc_hd__a22o_1 _8629_ (.A1(_3644_),
    .A2(_3821_),
    .B1(_3860_),
    .B2(_3861_),
    .X(net478));
 sky130_fd_sc_hd__a221o_1 _8630_ (.A1(_3253_),
    .A2(_3825_),
    .B1(_3256_),
    .B2(_3827_),
    .C1(_3831_),
    .X(_3862_));
 sky130_fd_sc_hd__o21a_1 _8631_ (.A1(_3833_),
    .A2(_3259_),
    .B1(_3834_),
    .X(_3863_));
 sky130_fd_sc_hd__a22o_1 _8632_ (.A1(_3251_),
    .A2(_3821_),
    .B1(_3862_),
    .B2(_3863_),
    .X(net480));
 sky130_fd_sc_hd__a22o_1 _8633_ (.A1(_3266_),
    .A2(_3824_),
    .B1(_3268_),
    .B2(_3826_),
    .X(_3864_));
 sky130_fd_sc_hd__mux2_1 _8634_ (.A0(_3864_),
    .A1(_3271_),
    .S(_3829_),
    .X(_3865_));
 sky130_fd_sc_hd__mux2_1 _8635_ (.A0(_3865_),
    .A1(_3264_),
    .S(_3819_),
    .X(_3866_));
 sky130_fd_sc_hd__buf_1 _8636_ (.A(_3866_),
    .X(net481));
 sky130_fd_sc_hd__a221o_1 _8637_ (.A1(_3279_),
    .A2(_3825_),
    .B1(_3281_),
    .B2(_3827_),
    .C1(_3830_),
    .X(_3867_));
 sky130_fd_sc_hd__o21a_1 _8638_ (.A1(_3833_),
    .A2(_3284_),
    .B1(_3834_),
    .X(_3868_));
 sky130_fd_sc_hd__a22o_1 _8639_ (.A1(_3277_),
    .A2(_3821_),
    .B1(_3867_),
    .B2(_3868_),
    .X(net482));
 sky130_fd_sc_hd__a22o_1 _8640_ (.A1(_3291_),
    .A2(_3824_),
    .B1(_3687_),
    .B2(_3826_),
    .X(_3869_));
 sky130_fd_sc_hd__mux2_1 _8641_ (.A0(_3869_),
    .A1(_3296_),
    .S(_3829_),
    .X(_3870_));
 sky130_fd_sc_hd__mux2_1 _8642_ (.A0(_3870_),
    .A1(_3289_),
    .S(_3819_),
    .X(_3871_));
 sky130_fd_sc_hd__buf_1 _8643_ (.A(_3871_),
    .X(net483));
 sky130_fd_sc_hd__a221o_1 _8644_ (.A1(_3303_),
    .A2(_3825_),
    .B1(_3305_),
    .B2(_3827_),
    .C1(_3830_),
    .X(_3872_));
 sky130_fd_sc_hd__o21a_1 _8645_ (.A1(_3833_),
    .A2(_3308_),
    .B1(_3834_),
    .X(_3873_));
 sky130_fd_sc_hd__a22o_1 _8646_ (.A1(_3301_),
    .A2(_3821_),
    .B1(_3872_),
    .B2(_3873_),
    .X(net484));
 sky130_fd_sc_hd__a2bb2o_1 _8647_ (.A1_N(_3822_),
    .A2_N(_3718_),
    .B1(_3315_),
    .B2(_3824_),
    .X(_3874_));
 sky130_fd_sc_hd__mux2_1 _8648_ (.A0(_3874_),
    .A1(_3320_),
    .S(_3829_),
    .X(_3875_));
 sky130_fd_sc_hd__mux2_1 _8649_ (.A0(_3875_),
    .A1(_3313_),
    .S(_3819_),
    .X(_3876_));
 sky130_fd_sc_hd__buf_1 _8650_ (.A(_3876_),
    .X(net485));
 sky130_fd_sc_hd__a221o_1 _8651_ (.A1(_3330_),
    .A2(_3825_),
    .B1(_3729_),
    .B2(_3827_),
    .C1(_3830_),
    .X(_3877_));
 sky130_fd_sc_hd__o21a_1 _8652_ (.A1(_3833_),
    .A2(_3336_),
    .B1(_3834_),
    .X(_3878_));
 sky130_fd_sc_hd__a22o_1 _8653_ (.A1(_3327_),
    .A2(_3821_),
    .B1(_3877_),
    .B2(_3878_),
    .X(net486));
 sky130_fd_sc_hd__a2bb2o_1 _8654_ (.A1_N(_3822_),
    .A2_N(_3738_),
    .B1(_3343_),
    .B2(_3824_),
    .X(_3879_));
 sky130_fd_sc_hd__mux2_1 _8655_ (.A0(_3879_),
    .A1(_3348_),
    .S(_3829_),
    .X(_3880_));
 sky130_fd_sc_hd__mux2_1 _8656_ (.A0(_3880_),
    .A1(_3341_),
    .S(_3819_),
    .X(_3881_));
 sky130_fd_sc_hd__buf_1 _8657_ (.A(_3881_),
    .X(net487));
 sky130_fd_sc_hd__a221o_1 _8658_ (.A1(_3355_),
    .A2(_3825_),
    .B1(_3357_),
    .B2(_3827_),
    .C1(_3830_),
    .X(_3882_));
 sky130_fd_sc_hd__o21a_1 _8659_ (.A1(_3833_),
    .A2(_3360_),
    .B1(_3834_),
    .X(_3883_));
 sky130_fd_sc_hd__a22o_1 _8660_ (.A1(_3353_),
    .A2(_3821_),
    .B1(_3882_),
    .B2(_3883_),
    .X(net488));
 sky130_fd_sc_hd__a22o_1 _8661_ (.A1(_3367_),
    .A2(_3824_),
    .B1(_3369_),
    .B2(_3826_),
    .X(_3884_));
 sky130_fd_sc_hd__mux2_1 _8662_ (.A0(_3884_),
    .A1(_3372_),
    .S(_3829_),
    .X(_3885_));
 sky130_fd_sc_hd__mux2_1 _8663_ (.A0(_3885_),
    .A1(_3365_),
    .S(_3819_),
    .X(_3886_));
 sky130_fd_sc_hd__buf_1 _8664_ (.A(_3886_),
    .X(net489));
 sky130_fd_sc_hd__a221o_1 _8665_ (.A1(_3379_),
    .A2(_3825_),
    .B1(_3381_),
    .B2(_3827_),
    .C1(_3830_),
    .X(_3887_));
 sky130_fd_sc_hd__o21a_1 _8666_ (.A1(_3833_),
    .A2(net731),
    .B1(_3834_),
    .X(_3888_));
 sky130_fd_sc_hd__a22o_1 _8667_ (.A1(_3377_),
    .A2(_3821_),
    .B1(_3887_),
    .B2(_3888_),
    .X(net491));
 sky130_fd_sc_hd__a221o_1 _8668_ (.A1(_3391_),
    .A2(_3824_),
    .B1(_3393_),
    .B2(_3827_),
    .C1(_3830_),
    .X(_3889_));
 sky130_fd_sc_hd__o21a_1 _8669_ (.A1(_3833_),
    .A2(_3396_),
    .B1(_3834_),
    .X(_3890_));
 sky130_fd_sc_hd__a22o_1 _8670_ (.A1(_3389_),
    .A2(_3821_),
    .B1(_3889_),
    .B2(_3890_),
    .X(net492));
 sky130_fd_sc_hd__a221o_1 _8671_ (.A1(_3403_),
    .A2(_3824_),
    .B1(_3405_),
    .B2(_3827_),
    .C1(_3830_),
    .X(_3891_));
 sky130_fd_sc_hd__o21a_1 _8672_ (.A1(_3833_),
    .A2(_3408_),
    .B1(_3834_),
    .X(_3892_));
 sky130_fd_sc_hd__a22o_1 _8673_ (.A1(_3401_),
    .A2(_3820_),
    .B1(_3891_),
    .B2(_3892_),
    .X(net493));
 sky130_fd_sc_hd__a22o_1 _8674_ (.A1(_3415_),
    .A2(_3823_),
    .B1(_3417_),
    .B2(_3826_),
    .X(_3893_));
 sky130_fd_sc_hd__mux2_1 _8675_ (.A0(_3893_),
    .A1(_3420_),
    .S(_3829_),
    .X(_3894_));
 sky130_fd_sc_hd__mux2_1 _8676_ (.A0(_3894_),
    .A1(_3413_),
    .S(_3819_),
    .X(_3895_));
 sky130_fd_sc_hd__buf_1 _8677_ (.A(_3895_),
    .X(net494));
 sky130_fd_sc_hd__a221o_1 _8678_ (.A1(_3434_),
    .A2(_3826_),
    .B1(_3791_),
    .B2(_3825_),
    .C1(_3830_),
    .X(_3896_));
 sky130_fd_sc_hd__a21oi_1 _8679_ (.A1(_3788_),
    .A2(_3831_),
    .B1(_3820_),
    .Y(_3897_));
 sky130_fd_sc_hd__a22o_1 _8680_ (.A1(_3786_),
    .A2(_3820_),
    .B1(_3896_),
    .B2(_3897_),
    .X(net495));
 sky130_fd_sc_hd__a221o_1 _8681_ (.A1(_3801_),
    .A2(_3824_),
    .B1(_3798_),
    .B2(_3827_),
    .C1(_3830_),
    .X(_3898_));
 sky130_fd_sc_hd__a21oi_1 _8682_ (.A1(_3795_),
    .A2(_3831_),
    .B1(_3820_),
    .Y(_3899_));
 sky130_fd_sc_hd__a22o_1 _8683_ (.A1(_3805_),
    .A2(_3820_),
    .B1(_3898_),
    .B2(_3899_),
    .X(net496));
 sky130_fd_sc_hd__a221o_1 _8684_ (.A1(_3471_),
    .A2(_3824_),
    .B1(_3474_),
    .B2(_3826_),
    .C1(_3830_),
    .X(_3900_));
 sky130_fd_sc_hd__nand2_1 _8685_ (.A(_3467_),
    .B(_3831_),
    .Y(_3901_));
 sky130_fd_sc_hd__and2_1 _8686_ (.A(_3480_),
    .B(_3820_),
    .X(_3902_));
 sky130_fd_sc_hd__a31o_1 _8687_ (.A1(_3900_),
    .A2(_3834_),
    .A3(_3901_),
    .B1(_3902_),
    .X(net497));
 sky130_fd_sc_hd__a22o_1 _8688_ (.A1(_3486_),
    .A2(_3823_),
    .B1(_3489_),
    .B2(_3826_),
    .X(_3903_));
 sky130_fd_sc_hd__mux2_1 _8689_ (.A0(_3903_),
    .A1(_3493_),
    .S(_3829_),
    .X(_3904_));
 sky130_fd_sc_hd__mux2_1 _8690_ (.A0(_3904_),
    .A1(_3483_),
    .S(_3819_),
    .X(_3905_));
 sky130_fd_sc_hd__buf_1 _8691_ (.A(_3905_),
    .X(net498));
 sky130_fd_sc_hd__a22o_1 _8692_ (.A1(_3499_),
    .A2(_3824_),
    .B1(_3501_),
    .B2(_3826_),
    .X(_3906_));
 sky130_fd_sc_hd__a32o_1 _8693_ (.A1(_3533_),
    .A2(_4239_),
    .A3(\arbiter.master_sel[2][1] ),
    .B1(_3833_),
    .B2(_3906_),
    .X(_3907_));
 sky130_fd_sc_hd__a32o_2 _8694_ (.A1(_0209_),
    .A2(\arbiter.master_sel[3][1] ),
    .A3(_3541_),
    .B1(_3907_),
    .B2(_3834_),
    .X(net499));
 sky130_fd_sc_hd__o31a_1 _8695_ (.A1(_0083_),
    .A2(_0120_),
    .A3(_3550_),
    .B1(_3818_),
    .X(_3908_));
 sky130_fd_sc_hd__nor2_1 _8696_ (.A(_3822_),
    .B(_3510_),
    .Y(_3909_));
 sky130_fd_sc_hd__a41o_1 _8697_ (.A1(_3552_),
    .A2(_0589_),
    .A3(\arbiter.master_sel[0][1] ),
    .A4(_3822_),
    .B1(_3909_),
    .X(_3910_));
 sky130_fd_sc_hd__nand2_1 _8698_ (.A(_3910_),
    .B(_3833_),
    .Y(_3911_));
 sky130_fd_sc_hd__o2bb2a_2 _8699_ (.A1_N(_3908_),
    .A2_N(_3911_),
    .B1(_3507_),
    .B2(_3834_),
    .X(net500));
 sky130_fd_sc_hd__a21oi_1 _8700_ (.A1(_0118_),
    .A2(_3831_),
    .B1(_3820_),
    .Y(_3912_));
 sky130_fd_sc_hd__a221o_1 _8701_ (.A1(_3519_),
    .A2(_3824_),
    .B1(_3520_),
    .B2(_3826_),
    .C1(_3830_),
    .X(_3913_));
 sky130_fd_sc_hd__a22o_1 _8702_ (.A1(_3912_),
    .A2(_3913_),
    .B1(_0206_),
    .B2(_3821_),
    .X(net367));
 sky130_fd_sc_hd__a221o_1 _8703_ (.A1(_3526_),
    .A2(_3826_),
    .B1(_3528_),
    .B2(_3825_),
    .C1(_3830_),
    .X(_3914_));
 sky130_fd_sc_hd__o21a_1 _8704_ (.A1(_3833_),
    .A2(_3531_),
    .B1(_3818_),
    .X(_3915_));
 sky130_fd_sc_hd__a22o_1 _8705_ (.A1(_3523_),
    .A2(_3820_),
    .B1(_3914_),
    .B2(_3915_),
    .X(net368));
 sky130_fd_sc_hd__nor2_2 _8706_ (.A(_0138_),
    .B(_0476_),
    .Y(_3916_));
 sky130_fd_sc_hd__buf_6 _8707_ (.A(_3916_),
    .X(_3917_));
 sky130_fd_sc_hd__clkbuf_8 _8708_ (.A(_3917_),
    .X(_3918_));
 sky130_fd_sc_hd__nor2_2 _8709_ (.A(_4184_),
    .B(_0625_),
    .Y(_3919_));
 sky130_fd_sc_hd__buf_4 _8710_ (.A(_3919_),
    .X(_3920_));
 sky130_fd_sc_hd__buf_4 _8711_ (.A(_3920_),
    .X(_3921_));
 sky130_fd_sc_hd__inv_2 _8712_ (.A(_3919_),
    .Y(_3922_));
 sky130_fd_sc_hd__and3_1 _8713_ (.A(_3922_),
    .B(_0588_),
    .C(_0433_),
    .X(_3923_));
 sky130_fd_sc_hd__clkbuf_4 _8714_ (.A(_3923_),
    .X(_3924_));
 sky130_fd_sc_hd__clkbuf_8 _8715_ (.A(_3924_),
    .X(_3925_));
 sky130_fd_sc_hd__nor2_8 _8716_ (.A(_0083_),
    .B(_0455_),
    .Y(_3926_));
 sky130_fd_sc_hd__buf_4 _8717_ (.A(_3926_),
    .X(_3927_));
 sky130_fd_sc_hd__a221o_1 _8718_ (.A1(_3083_),
    .A2(_3921_),
    .B1(_3577_),
    .B2(_3925_),
    .C1(_3927_),
    .X(_3928_));
 sky130_fd_sc_hd__a21oi_1 _8719_ (.A1(_3571_),
    .A2(_3927_),
    .B1(_3917_),
    .Y(_3929_));
 sky130_fd_sc_hd__a22o_1 _8720_ (.A1(_3567_),
    .A2(_3918_),
    .B1(_3928_),
    .B2(_3929_),
    .X(net369));
 sky130_fd_sc_hd__a221o_1 _8721_ (.A1(_3582_),
    .A2(_3925_),
    .B1(_3586_),
    .B2(_3921_),
    .C1(_3927_),
    .X(_3930_));
 sky130_fd_sc_hd__inv_2 _8722_ (.A(_3926_),
    .Y(_3931_));
 sky130_fd_sc_hd__buf_4 _8723_ (.A(_3931_),
    .X(_3932_));
 sky130_fd_sc_hd__inv_2 _8724_ (.A(_3916_),
    .Y(_3933_));
 sky130_fd_sc_hd__buf_4 _8725_ (.A(_3933_),
    .X(_3934_));
 sky130_fd_sc_hd__o21a_1 _8726_ (.A1(_3932_),
    .A2(_3590_),
    .B1(_3934_),
    .X(_3935_));
 sky130_fd_sc_hd__a22o_1 _8727_ (.A1(_3593_),
    .A2(_3918_),
    .B1(_3930_),
    .B2(_3935_),
    .X(net370));
 sky130_fd_sc_hd__a221o_1 _8728_ (.A1(_3108_),
    .A2(_3925_),
    .B1(_3110_),
    .B2(_3921_),
    .C1(_3927_),
    .X(_3936_));
 sky130_fd_sc_hd__a21oi_1 _8729_ (.A1(_3113_),
    .A2(_3927_),
    .B1(_3917_),
    .Y(_3937_));
 sky130_fd_sc_hd__a22o_1 _8730_ (.A1(_3106_),
    .A2(_3918_),
    .B1(_3936_),
    .B2(_3937_),
    .X(net371));
 sky130_fd_sc_hd__o21ai_1 _8731_ (.A1(_3932_),
    .A2(_3123_),
    .B1(_3934_),
    .Y(_3938_));
 sky130_fd_sc_hd__a22o_1 _8732_ (.A1(_3118_),
    .A2(_3924_),
    .B1(_3120_),
    .B2(_3920_),
    .X(_3939_));
 sky130_fd_sc_hd__and2_1 _8733_ (.A(_3939_),
    .B(_3932_),
    .X(_3940_));
 sky130_fd_sc_hd__o22a_1 _8734_ (.A1(_3116_),
    .A2(_3934_),
    .B1(_3938_),
    .B2(_3940_),
    .X(net372));
 sky130_fd_sc_hd__a221o_1 _8735_ (.A1(_3133_),
    .A2(_3921_),
    .B1(_3140_),
    .B2(_3925_),
    .C1(_3927_),
    .X(_3941_));
 sky130_fd_sc_hd__a21oi_1 _8736_ (.A1(_3145_),
    .A2(_3927_),
    .B1(_3917_),
    .Y(_3942_));
 sky130_fd_sc_hd__a22o_1 _8737_ (.A1(_3129_),
    .A2(_3918_),
    .B1(_3941_),
    .B2(_3942_),
    .X(net373));
 sky130_fd_sc_hd__inv_2 _8738_ (.A(_3924_),
    .Y(_3943_));
 sky130_fd_sc_hd__o221a_1 _8739_ (.A1(_3922_),
    .A2(_3162_),
    .B1(_3157_),
    .B2(_3943_),
    .C1(_3931_),
    .X(_3944_));
 sky130_fd_sc_hd__a211o_1 _8740_ (.A1(_3152_),
    .A2(_3927_),
    .B1(_3917_),
    .C1(_3944_),
    .X(_3945_));
 sky130_fd_sc_hd__o21ai_2 _8741_ (.A1(_3168_),
    .A2(_3934_),
    .B1(_3945_),
    .Y(net374));
 sky130_fd_sc_hd__a221o_1 _8742_ (.A1(_3175_),
    .A2(_3925_),
    .B1(_3177_),
    .B2(_3921_),
    .C1(_3927_),
    .X(_3946_));
 sky130_fd_sc_hd__o21a_1 _8743_ (.A1(_3932_),
    .A2(_3184_),
    .B1(_3933_),
    .X(_3947_));
 sky130_fd_sc_hd__a22o_1 _8744_ (.A1(_3173_),
    .A2(_3918_),
    .B1(_3946_),
    .B2(_3947_),
    .X(net375));
 sky130_fd_sc_hd__a221o_1 _8745_ (.A1(_3193_),
    .A2(_3924_),
    .B1(_3195_),
    .B2(_3920_),
    .C1(_3926_),
    .X(_3948_));
 sky130_fd_sc_hd__o21a_1 _8746_ (.A1(_3602_),
    .A2(_3931_),
    .B1(_3948_),
    .X(_3949_));
 sky130_fd_sc_hd__mux2_1 _8747_ (.A0(_3949_),
    .A1(_3191_),
    .S(_3917_),
    .X(_3950_));
 sky130_fd_sc_hd__buf_1 _8748_ (.A(_3950_),
    .X(net376));
 sky130_fd_sc_hd__a221o_1 _8749_ (.A1(_3207_),
    .A2(_3921_),
    .B1(_3628_),
    .B2(_3925_),
    .C1(_3927_),
    .X(_3951_));
 sky130_fd_sc_hd__o21a_1 _8750_ (.A1(_3932_),
    .A2(_3632_),
    .B1(_3933_),
    .X(_3952_));
 sky130_fd_sc_hd__a22o_1 _8751_ (.A1(_3638_),
    .A2(_3918_),
    .B1(_3951_),
    .B2(_3952_),
    .X(net378));
 sky130_fd_sc_hd__a221o_1 _8752_ (.A1(_3649_),
    .A2(_3921_),
    .B1(_3651_),
    .B2(_3925_),
    .C1(_3927_),
    .X(_3953_));
 sky130_fd_sc_hd__a21oi_1 _8753_ (.A1(_3646_),
    .A2(_3927_),
    .B1(_3917_),
    .Y(_3954_));
 sky130_fd_sc_hd__a22o_1 _8754_ (.A1(_3644_),
    .A2(_3918_),
    .B1(_3953_),
    .B2(_3954_),
    .X(net379));
 sky130_fd_sc_hd__and3_2 _8755_ (.A(_3922_),
    .B(_3574_),
    .C(_0588_),
    .X(_3955_));
 sky130_fd_sc_hd__a221o_1 _8756_ (.A1(_3231_),
    .A2(_3920_),
    .B1(_3660_),
    .B2(_3955_),
    .C1(_3926_),
    .X(_3956_));
 sky130_fd_sc_hd__o211a_1 _8757_ (.A1(_3234_),
    .A2(_3932_),
    .B1(_3933_),
    .C1(_3956_),
    .X(_3957_));
 sky130_fd_sc_hd__a31o_1 _8758_ (.A1(_0470_),
    .A2(_3227_),
    .A3(_3917_),
    .B1(_3957_),
    .X(net380));
 sky130_fd_sc_hd__nor2_2 _8759_ (.A(_0138_),
    .B(_3565_),
    .Y(_3958_));
 sky130_fd_sc_hd__a22o_1 _8760_ (.A1(_3243_),
    .A2(_3920_),
    .B1(_3671_),
    .B2(_3955_),
    .X(_3959_));
 sky130_fd_sc_hd__clkbuf_8 _8761_ (.A(_3926_),
    .X(_3960_));
 sky130_fd_sc_hd__mux2_1 _8762_ (.A0(_3959_),
    .A1(_3246_),
    .S(_3960_),
    .X(_3961_));
 sky130_fd_sc_hd__a22o_1 _8763_ (.A1(_3665_),
    .A2(_3958_),
    .B1(_3961_),
    .B2(_3934_),
    .X(net381));
 sky130_fd_sc_hd__a221o_1 _8764_ (.A1(_3256_),
    .A2(_3920_),
    .B1(_3681_),
    .B2(_3955_),
    .C1(_3960_),
    .X(_3962_));
 sky130_fd_sc_hd__or2_1 _8765_ (.A(_3931_),
    .B(_3259_),
    .X(_3963_));
 sky130_fd_sc_hd__a32o_1 _8766_ (.A1(_3962_),
    .A2(_3934_),
    .A3(_3963_),
    .B1(_3677_),
    .B2(_3958_),
    .X(net382));
 sky130_fd_sc_hd__a32o_1 _8767_ (.A1(_3266_),
    .A2(_0427_),
    .A3(_3924_),
    .B1(_3268_),
    .B2(_3920_),
    .X(_3964_));
 sky130_fd_sc_hd__mux2_1 _8768_ (.A0(_3964_),
    .A1(_3271_),
    .S(_3960_),
    .X(_3965_));
 sky130_fd_sc_hd__a22o_1 _8769_ (.A1(_3697_),
    .A2(_3958_),
    .B1(_3965_),
    .B2(_3934_),
    .X(net383));
 sky130_fd_sc_hd__and2b_1 _8770_ (.A_N(_3707_),
    .B(_3955_),
    .X(_3966_));
 sky130_fd_sc_hd__a211o_1 _8771_ (.A1(_3281_),
    .A2(_3920_),
    .B1(_3960_),
    .C1(_3966_),
    .X(_3967_));
 sky130_fd_sc_hd__or2_1 _8772_ (.A(_3931_),
    .B(_3284_),
    .X(_3968_));
 sky130_fd_sc_hd__a32o_1 _8773_ (.A1(_3967_),
    .A2(_3934_),
    .A3(_3968_),
    .B1(_3702_),
    .B2(_3958_),
    .X(net384));
 sky130_fd_sc_hd__a221o_1 _8774_ (.A1(_3293_),
    .A2(_3921_),
    .B1(_3669_),
    .B2(_3925_),
    .C1(_3927_),
    .X(_3969_));
 sky130_fd_sc_hd__o21a_1 _8775_ (.A1(_3932_),
    .A2(_3296_),
    .B1(_3933_),
    .X(_3970_));
 sky130_fd_sc_hd__a22o_1 _8776_ (.A1(_3289_),
    .A2(_3918_),
    .B1(_3969_),
    .B2(_3970_),
    .X(net385));
 sky130_fd_sc_hd__a21o_1 _8777_ (.A1(_3305_),
    .A2(_3920_),
    .B1(_3926_),
    .X(_3971_));
 sky130_fd_sc_hd__a41o_1 _8778_ (.A1(_3680_),
    .A2(_0589_),
    .A3(_0433_),
    .A4(_3922_),
    .B1(_3971_),
    .X(_3972_));
 sky130_fd_sc_hd__o21a_1 _8779_ (.A1(_3932_),
    .A2(_3308_),
    .B1(_3933_),
    .X(_3973_));
 sky130_fd_sc_hd__a22o_1 _8780_ (.A1(_3301_),
    .A2(_3918_),
    .B1(_3972_),
    .B2(_3973_),
    .X(net386));
 sky130_fd_sc_hd__a221o_1 _8781_ (.A1(_3317_),
    .A2(_3920_),
    .B1(_3743_),
    .B2(_3955_),
    .C1(_3960_),
    .X(_3974_));
 sky130_fd_sc_hd__or2_1 _8782_ (.A(_3931_),
    .B(_3320_),
    .X(_3975_));
 sky130_fd_sc_hd__a32o_1 _8783_ (.A1(_3974_),
    .A2(_3934_),
    .A3(_3975_),
    .B1(_3736_),
    .B2(_3958_),
    .X(net387));
 sky130_fd_sc_hd__a22o_1 _8784_ (.A1(_3704_),
    .A2(_3924_),
    .B1(_3333_),
    .B2(_3920_),
    .X(_3976_));
 sky130_fd_sc_hd__mux2_1 _8785_ (.A0(_3976_),
    .A1(_3336_),
    .S(_3960_),
    .X(_3977_));
 sky130_fd_sc_hd__a22o_1 _8786_ (.A1(_3750_),
    .A2(_3958_),
    .B1(_3977_),
    .B2(_3934_),
    .X(net389));
 sky130_fd_sc_hd__a22o_1 _8787_ (.A1(_3345_),
    .A2(_3920_),
    .B1(_3761_),
    .B2(_3955_),
    .X(_3978_));
 sky130_fd_sc_hd__mux2_1 _8788_ (.A0(_3978_),
    .A1(_3348_),
    .S(_3960_),
    .X(_3979_));
 sky130_fd_sc_hd__a22o_1 _8789_ (.A1(_3757_),
    .A2(_3958_),
    .B1(_3979_),
    .B2(_3934_),
    .X(net390));
 sky130_fd_sc_hd__a221o_1 _8790_ (.A1(_3355_),
    .A2(_3925_),
    .B1(_3357_),
    .B2(_3921_),
    .C1(_3960_),
    .X(_3980_));
 sky130_fd_sc_hd__o21a_1 _8791_ (.A1(_3932_),
    .A2(_3360_),
    .B1(_3933_),
    .X(_3981_));
 sky130_fd_sc_hd__a22o_1 _8792_ (.A1(_3353_),
    .A2(_3918_),
    .B1(_3980_),
    .B2(_3981_),
    .X(net391));
 sky130_fd_sc_hd__a22o_1 _8793_ (.A1(_3367_),
    .A2(_3924_),
    .B1(_3369_),
    .B2(_3920_),
    .X(_3982_));
 sky130_fd_sc_hd__mux2_1 _8794_ (.A0(_3982_),
    .A1(_3372_),
    .S(_3926_),
    .X(_3983_));
 sky130_fd_sc_hd__mux2_1 _8795_ (.A0(_3983_),
    .A1(_3365_),
    .S(_3917_),
    .X(_3984_));
 sky130_fd_sc_hd__buf_1 _8796_ (.A(_3984_),
    .X(net392));
 sky130_fd_sc_hd__a221o_1 _8797_ (.A1(_3379_),
    .A2(_3925_),
    .B1(_3381_),
    .B2(_3921_),
    .C1(_3960_),
    .X(_3985_));
 sky130_fd_sc_hd__o21a_1 _8798_ (.A1(_3932_),
    .A2(net731),
    .B1(_3933_),
    .X(_3986_));
 sky130_fd_sc_hd__a22o_1 _8799_ (.A1(_3377_),
    .A2(_3918_),
    .B1(_3985_),
    .B2(_3986_),
    .X(net393));
 sky130_fd_sc_hd__a221o_1 _8800_ (.A1(_3391_),
    .A2(_3925_),
    .B1(_3393_),
    .B2(_3921_),
    .C1(_3960_),
    .X(_3987_));
 sky130_fd_sc_hd__o21a_1 _8801_ (.A1(_3932_),
    .A2(_3396_),
    .B1(_3933_),
    .X(_3988_));
 sky130_fd_sc_hd__a22o_1 _8802_ (.A1(_3389_),
    .A2(_3918_),
    .B1(_3987_),
    .B2(_3988_),
    .X(net394));
 sky130_fd_sc_hd__nand2_1 _8803_ (.A(_3791_),
    .B(_3925_),
    .Y(_3989_));
 sky130_fd_sc_hd__a21oi_1 _8804_ (.A1(_3405_),
    .A2(_3921_),
    .B1(_3960_),
    .Y(_3990_));
 sky130_fd_sc_hd__a22o_1 _8805_ (.A1(_3788_),
    .A2(_3960_),
    .B1(_3989_),
    .B2(_3990_),
    .X(_3991_));
 sky130_fd_sc_hd__nand2_1 _8806_ (.A(_3786_),
    .B(_3918_),
    .Y(_3992_));
 sky130_fd_sc_hd__o21ai_4 _8807_ (.A1(_3917_),
    .A2(_3991_),
    .B1(_3992_),
    .Y(net395));
 sky130_fd_sc_hd__a2bb2o_1 _8808_ (.A1_N(_3799_),
    .A2_N(_3943_),
    .B1(_3919_),
    .B2(_3798_),
    .X(_3993_));
 sky130_fd_sc_hd__mux2_1 _8809_ (.A0(_3993_),
    .A1(_3796_),
    .S(_3926_),
    .X(_3994_));
 sky130_fd_sc_hd__mux2_2 _8810_ (.A0(_3994_),
    .A1(_3778_),
    .S(_3917_),
    .X(_3995_));
 sky130_fd_sc_hd__buf_1 _8811_ (.A(_3995_),
    .X(net396));
 sky130_fd_sc_hd__a221o_1 _8812_ (.A1(_3431_),
    .A2(_3925_),
    .B1(_3434_),
    .B2(_3921_),
    .C1(_3960_),
    .X(_3996_));
 sky130_fd_sc_hd__a21oi_1 _8813_ (.A1(_3439_),
    .A2(_3927_),
    .B1(_3917_),
    .Y(_3997_));
 sky130_fd_sc_hd__a22o_1 _8814_ (.A1(_3423_),
    .A2(_3918_),
    .B1(_3996_),
    .B2(_3997_),
    .X(net397));
 sky130_fd_sc_hd__o21ai_1 _8815_ (.A1(_3932_),
    .A2(_3460_),
    .B1(_3934_),
    .Y(_3998_));
 sky130_fd_sc_hd__a22o_1 _8816_ (.A1(_3450_),
    .A2(_3924_),
    .B1(_3454_),
    .B2(_3920_),
    .X(_3999_));
 sky130_fd_sc_hd__and2_1 _8817_ (.A(_3999_),
    .B(_3932_),
    .X(_4000_));
 sky130_fd_sc_hd__o22a_2 _8818_ (.A1(_3442_),
    .A2(_3934_),
    .B1(_3998_),
    .B2(_4000_),
    .X(net398));
 sky130_fd_sc_hd__a221o_1 _8819_ (.A1(_3471_),
    .A2(_3925_),
    .B1(_3474_),
    .B2(_3921_),
    .C1(_3960_),
    .X(_4001_));
 sky130_fd_sc_hd__nand2_1 _8820_ (.A(_3467_),
    .B(_3927_),
    .Y(_4002_));
 sky130_fd_sc_hd__and2_1 _8821_ (.A(_3480_),
    .B(_3917_),
    .X(_4003_));
 sky130_fd_sc_hd__a31o_1 _8822_ (.A1(_4001_),
    .A2(_3934_),
    .A3(_4002_),
    .B1(_4003_),
    .X(net400));
 sky130_fd_sc_hd__a22o_1 _8823_ (.A1(_3486_),
    .A2(_3924_),
    .B1(_3489_),
    .B2(_3919_),
    .X(_4004_));
 sky130_fd_sc_hd__mux2_1 _8824_ (.A0(_4004_),
    .A1(_3493_),
    .S(_3926_),
    .X(_4005_));
 sky130_fd_sc_hd__mux2_1 _8825_ (.A0(_4005_),
    .A1(_3483_),
    .S(_3917_),
    .X(_4006_));
 sky130_fd_sc_hd__clkbuf_2 _8826_ (.A(_4006_),
    .X(net401));
 sky130_fd_sc_hd__a221o_1 _8827_ (.A1(_3499_),
    .A2(_3924_),
    .B1(_3501_),
    .B2(_3920_),
    .C1(_3926_),
    .X(_4007_));
 sky130_fd_sc_hd__o21a_1 _8828_ (.A1(_3504_),
    .A2(_3931_),
    .B1(_4007_),
    .X(_4008_));
 sky130_fd_sc_hd__mux2_1 _8829_ (.A0(_4008_),
    .A1(_3497_),
    .S(_3917_),
    .X(_4009_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _8830_ (.A(_4009_),
    .X(net402));
 sky130_fd_sc_hd__o21ai_1 _8831_ (.A1(_3932_),
    .A2(_3516_),
    .B1(_3934_),
    .Y(_4010_));
 sky130_fd_sc_hd__a22o_1 _8832_ (.A1(_3511_),
    .A2(_3920_),
    .B1(_3513_),
    .B2(_3924_),
    .X(_4011_));
 sky130_fd_sc_hd__and2_1 _8833_ (.A(_4011_),
    .B(_3932_),
    .X(_4012_));
 sky130_fd_sc_hd__o22a_2 _8834_ (.A1(_3507_),
    .A2(_3934_),
    .B1(_4010_),
    .B2(_4012_),
    .X(net403));
 sky130_fd_sc_hd__a21oi_1 _8835_ (.A1(_0118_),
    .A2(_3927_),
    .B1(_3917_),
    .Y(_4013_));
 sky130_fd_sc_hd__a221o_1 _8836_ (.A1(_3519_),
    .A2(_3925_),
    .B1(_3520_),
    .B2(_3921_),
    .C1(_3960_),
    .X(_4014_));
 sky130_fd_sc_hd__a22o_2 _8837_ (.A1(_4013_),
    .A2(_4014_),
    .B1(_0206_),
    .B2(_3918_),
    .X(net404));
 sky130_fd_sc_hd__a221o_1 _8838_ (.A1(_3526_),
    .A2(_3921_),
    .B1(_3528_),
    .B2(_3925_),
    .C1(_3960_),
    .X(_4015_));
 sky130_fd_sc_hd__o21a_1 _8839_ (.A1(_3932_),
    .A2(_3531_),
    .B1(_3933_),
    .X(_4016_));
 sky130_fd_sc_hd__a22o_1 _8840_ (.A1(_3523_),
    .A2(_3918_),
    .B1(_4015_),
    .B2(_4016_),
    .X(net405));
 sky130_fd_sc_hd__a21oi_1 _8841_ (.A1(_0139_),
    .A2(_0373_),
    .B1(_0165_),
    .Y(_4017_));
 sky130_fd_sc_hd__nand2_1 _8842_ (.A(_0137_),
    .B(_0855_),
    .Y(_4018_));
 sky130_fd_sc_hd__a21bo_1 _8843_ (.A1(_4018_),
    .A2(_0164_),
    .B1_N(_0147_),
    .X(_4019_));
 sky130_fd_sc_hd__nand2_1 _8844_ (.A(_4019_),
    .B(_0157_),
    .Y(_4020_));
 sky130_fd_sc_hd__nand3_1 _8845_ (.A(_0137_),
    .B(_0164_),
    .C(_0199_),
    .Y(_4021_));
 sky130_fd_sc_hd__nand2_1 _8846_ (.A(_0147_),
    .B(_0157_),
    .Y(_4022_));
 sky130_fd_sc_hd__inv_2 _8847_ (.A(_4022_),
    .Y(_4023_));
 sky130_fd_sc_hd__nand2_1 _8848_ (.A(_4021_),
    .B(_4023_),
    .Y(_4024_));
 sky130_fd_sc_hd__inv_2 _8849_ (.A(_4024_),
    .Y(_4025_));
 sky130_fd_sc_hd__nor2_1 _8850_ (.A(_0174_),
    .B(_4025_),
    .Y(_4026_));
 sky130_fd_sc_hd__nand2_1 _8851_ (.A(_4020_),
    .B(_4026_),
    .Y(_4027_));
 sky130_fd_sc_hd__o21a_1 _8852_ (.A1(_4017_),
    .A2(_4027_),
    .B1(_0156_),
    .X(_4028_));
 sky130_fd_sc_hd__a211o_1 _8853_ (.A1(_0208_),
    .A2(_2439_),
    .B1(_1757_),
    .C1(_0156_),
    .X(_4029_));
 sky130_fd_sc_hd__o21ai_1 _8854_ (.A1(_0483_),
    .A2(_4028_),
    .B1(_4029_),
    .Y(_0032_));
 sky130_fd_sc_hd__nor2_1 _8855_ (.A(_4017_),
    .B(_4020_),
    .Y(_4030_));
 sky130_fd_sc_hd__nand2_1 _8856_ (.A(_4030_),
    .B(_4026_),
    .Y(_4031_));
 sky130_fd_sc_hd__nand2_1 _8857_ (.A(_0208_),
    .B(_0652_),
    .Y(_4032_));
 sky130_fd_sc_hd__a31o_1 _8858_ (.A1(_0142_),
    .A2(_0145_),
    .A3(_4032_),
    .B1(_1757_),
    .X(_4033_));
 sky130_fd_sc_hd__a21boi_1 _8859_ (.A1(_4031_),
    .A2(_0146_),
    .B1_N(_4033_),
    .Y(_0033_));
 sky130_fd_sc_hd__nor2_1 _8860_ (.A(_0174_),
    .B(_4024_),
    .Y(_4034_));
 sky130_fd_sc_hd__nand2_1 _8861_ (.A(_4020_),
    .B(_4034_),
    .Y(_4035_));
 sky130_fd_sc_hd__o21ai_1 _8862_ (.A1(_4017_),
    .A2(_4035_),
    .B1(_0163_),
    .Y(_4036_));
 sky130_fd_sc_hd__a211o_1 _8863_ (.A1(_0208_),
    .A2(_0767_),
    .B1(_1757_),
    .C1(_0163_),
    .X(_4037_));
 sky130_fd_sc_hd__a21bo_1 _8864_ (.A1(_4036_),
    .A2(_1757_),
    .B1_N(_4037_),
    .X(_0034_));
 sky130_fd_sc_hd__nand2_1 _8865_ (.A(_4030_),
    .B(_4034_),
    .Y(_4038_));
 sky130_fd_sc_hd__a21o_1 _8866_ (.A1(_4038_),
    .A2(_0136_),
    .B1(_0483_),
    .X(_4039_));
 sky130_fd_sc_hd__a211o_1 _8867_ (.A1(_0194_),
    .A2(_0208_),
    .B1(_1757_),
    .C1(_0136_),
    .X(_4040_));
 sky130_fd_sc_hd__nand2_1 _8868_ (.A(_4039_),
    .B(_4040_),
    .Y(_0035_));
 sky130_fd_sc_hd__or2_1 _8869_ (.A(net763),
    .B(_0356_),
    .X(_4041_));
 sky130_fd_sc_hd__nand2_1 _8870_ (.A(_0363_),
    .B(_0368_),
    .Y(_4042_));
 sky130_fd_sc_hd__inv_2 _8871_ (.A(_4042_),
    .Y(_4043_));
 sky130_fd_sc_hd__nand2_1 _8872_ (.A(_4041_),
    .B(_4043_),
    .Y(_4044_));
 sky130_fd_sc_hd__inv_2 _8873_ (.A(_4044_),
    .Y(_4045_));
 sky130_fd_sc_hd__nor2_1 _8874_ (.A(_0174_),
    .B(_4045_),
    .Y(_4046_));
 sky130_fd_sc_hd__nand2_1 _8875_ (.A(_0345_),
    .B(_0183_),
    .Y(_4047_));
 sky130_fd_sc_hd__a21bo_1 _8876_ (.A1(_4047_),
    .A2(_0355_),
    .B1_N(_0368_),
    .X(_4048_));
 sky130_fd_sc_hd__nand2_1 _8877_ (.A(_4048_),
    .B(_0363_),
    .Y(_4049_));
 sky130_fd_sc_hd__a211o_1 _8878_ (.A1(net751),
    .A2(_0138_),
    .B1(_4042_),
    .C1(_0356_),
    .X(_4050_));
 sky130_fd_sc_hd__nand3_1 _8879_ (.A(_4046_),
    .B(_4049_),
    .C(_4050_),
    .Y(_4051_));
 sky130_fd_sc_hd__inv_2 _8880_ (.A(_0210_),
    .Y(_4052_));
 sky130_fd_sc_hd__a21o_1 _8881_ (.A1(_4051_),
    .A2(_0362_),
    .B1(_4052_),
    .X(_4053_));
 sky130_fd_sc_hd__o31ai_1 _8882_ (.A1(_4150_),
    .A2(_0470_),
    .A3(_0206_),
    .B1(_0209_),
    .Y(_4054_));
 sky130_fd_sc_hd__a21o_1 _8883_ (.A1(_0166_),
    .A2(_4054_),
    .B1(_0362_),
    .X(_4055_));
 sky130_fd_sc_hd__nand2_1 _8884_ (.A(_4053_),
    .B(_4055_),
    .Y(_0028_));
 sky130_fd_sc_hd__inv_2 _8885_ (.A(_4049_),
    .Y(_4056_));
 sky130_fd_sc_hd__nand3_1 _8886_ (.A(_4046_),
    .B(_4056_),
    .C(_4050_),
    .Y(_4057_));
 sky130_fd_sc_hd__nand2_1 _8887_ (.A(_0364_),
    .B(_0367_),
    .Y(_4058_));
 sky130_fd_sc_hd__inv_2 _8888_ (.A(_4058_),
    .Y(_4059_));
 sky130_fd_sc_hd__a21o_1 _8889_ (.A1(_4057_),
    .A2(_4059_),
    .B1(_4052_),
    .X(_4060_));
 sky130_fd_sc_hd__a31o_1 _8890_ (.A1(_0205_),
    .A2(_0124_),
    .A3(_0184_),
    .B1(_0138_),
    .X(_4061_));
 sky130_fd_sc_hd__a21o_1 _8891_ (.A1(_0166_),
    .A2(_4061_),
    .B1(_4059_),
    .X(_4062_));
 sky130_fd_sc_hd__nand2_1 _8892_ (.A(_4060_),
    .B(_4062_),
    .Y(_0029_));
 sky130_fd_sc_hd__nor2_1 _8893_ (.A(_0174_),
    .B(_4044_),
    .Y(_4063_));
 sky130_fd_sc_hd__nand3_1 _8894_ (.A(_4050_),
    .B(_4063_),
    .C(_4049_),
    .Y(_4064_));
 sky130_fd_sc_hd__a21o_1 _8895_ (.A1(_4064_),
    .A2(_0354_),
    .B1(_4052_),
    .X(_4065_));
 sky130_fd_sc_hd__o31ai_1 _8896_ (.A1(net74),
    .A2(_0480_),
    .A3(_0206_),
    .B1(_0209_),
    .Y(_4066_));
 sky130_fd_sc_hd__a21o_1 _8897_ (.A1(_0166_),
    .A2(_4066_),
    .B1(_0354_),
    .X(_4067_));
 sky130_fd_sc_hd__nand2_1 _8898_ (.A(_4065_),
    .B(_4067_),
    .Y(_0030_));
 sky130_fd_sc_hd__nand3_1 _8899_ (.A(_4056_),
    .B(_4050_),
    .C(_4063_),
    .Y(_4068_));
 sky130_fd_sc_hd__a21o_1 _8900_ (.A1(_4068_),
    .A2(_0344_),
    .B1(_4052_),
    .X(_4069_));
 sky130_fd_sc_hd__o31ai_1 _8901_ (.A1(net138),
    .A2(_0476_),
    .A3(_0206_),
    .B1(_0209_),
    .Y(_4070_));
 sky130_fd_sc_hd__a21o_1 _8902_ (.A1(_0166_),
    .A2(_4070_),
    .B1(_0344_),
    .X(_4071_));
 sky130_fd_sc_hd__nand2_1 _8903_ (.A(_4069_),
    .B(_4071_),
    .Y(_0031_));
 sky130_fd_sc_hd__nor2_1 _8904_ (.A(_0125_),
    .B(_0380_),
    .Y(_4072_));
 sky130_fd_sc_hd__a31o_1 _8905_ (.A1(_0328_),
    .A2(_0291_),
    .A3(_0380_),
    .B1(_4072_),
    .X(_0002_));
 sky130_fd_sc_hd__o2bb2a_1 _8906_ (.A1_N(_0341_),
    .A2_N(_0357_),
    .B1(net754),
    .B2(_0380_),
    .X(_0003_));
 sky130_fd_sc_hd__mux2_1 _8907_ (.A0(_4056_),
    .A1(net764),
    .S(_0211_),
    .X(_4073_));
 sky130_fd_sc_hd__clkbuf_1 _8908_ (.A(_4073_),
    .X(_0004_));
 sky130_fd_sc_hd__mux2_1 _8909_ (.A0(_4045_),
    .A1(net763),
    .S(_0211_),
    .X(_4074_));
 sky130_fd_sc_hd__clkbuf_1 _8910_ (.A(_4074_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _8911_ (.A0(_0060_),
    .A1(_0558_),
    .S(_4236_),
    .X(_4075_));
 sky130_fd_sc_hd__clkbuf_1 _8912_ (.A(_4075_),
    .X(_0006_));
 sky130_fd_sc_hd__nand2_1 _8913_ (.A(_4236_),
    .B(net756),
    .Y(_4076_));
 sky130_fd_sc_hd__o21ai_1 _8914_ (.A1(_4236_),
    .A2(_4247_),
    .B1(net757),
    .Y(_0007_));
 sky130_fd_sc_hd__mux2_1 _8915_ (.A0(_4216_),
    .A1(_0523_),
    .S(_4181_),
    .X(_4077_));
 sky130_fd_sc_hd__clkbuf_1 _8916_ (.A(_4077_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _8917_ (.A0(_4207_),
    .A1(_4118_),
    .S(_4181_),
    .X(_4078_));
 sky130_fd_sc_hd__clkbuf_1 _8918_ (.A(net771),
    .X(_0009_));
 sky130_fd_sc_hd__nand2_1 _8919_ (.A(_0287_),
    .B(net743),
    .Y(_4079_));
 sky130_fd_sc_hd__mux2_1 _8920_ (.A0(_0294_),
    .A1(net769),
    .S(_4079_),
    .X(_4080_));
 sky130_fd_sc_hd__clkbuf_1 _8921_ (.A(_4080_),
    .X(_0010_));
 sky130_fd_sc_hd__nand2_1 _8922_ (.A(_4079_),
    .B(net748),
    .Y(_4081_));
 sky130_fd_sc_hd__o21ai_1 _8923_ (.A1(_4079_),
    .A2(_0304_),
    .B1(net749),
    .Y(_0011_));
 sky130_fd_sc_hd__nand2_1 _8924_ (.A(_0169_),
    .B(_0769_),
    .Y(_4082_));
 sky130_fd_sc_hd__o21ai_1 _8925_ (.A1(_0169_),
    .A2(_4020_),
    .B1(_4082_),
    .Y(_0012_));
 sky130_fd_sc_hd__mux2_1 _8926_ (.A0(_4025_),
    .A1(net777),
    .S(_0169_),
    .X(_4083_));
 sky130_fd_sc_hd__clkbuf_1 _8927_ (.A(_4083_),
    .X(_0013_));
 sky130_fd_sc_hd__o21ai_1 _8928_ (.A1(_0180_),
    .A2(_0388_),
    .B1(net740),
    .Y(_4084_));
 sky130_fd_sc_hd__nor2_1 _8929_ (.A(_0398_),
    .B(_0393_),
    .Y(_4085_));
 sky130_fd_sc_hd__nand3_1 _8930_ (.A(_0390_),
    .B(_0391_),
    .C(_4085_),
    .Y(_4086_));
 sky130_fd_sc_hd__nand2_1 _8931_ (.A(net741),
    .B(_4086_),
    .Y(_0014_));
 sky130_fd_sc_hd__o21ai_1 _8932_ (.A1(_0180_),
    .A2(_0388_),
    .B1(net743),
    .Y(_4087_));
 sky130_fd_sc_hd__and2_1 _8933_ (.A(_0396_),
    .B(_0401_),
    .X(_4088_));
 sky130_fd_sc_hd__nand3_1 _8934_ (.A(_0390_),
    .B(_0391_),
    .C(_4088_),
    .Y(_4089_));
 sky130_fd_sc_hd__nand2_1 _8935_ (.A(net744),
    .B(_4089_),
    .Y(_0015_));
 sky130_fd_sc_hd__nand2_1 _8936_ (.A(_4165_),
    .B(net759),
    .Y(_4090_));
 sky130_fd_sc_hd__o21ai_1 _8937_ (.A1(_4165_),
    .A2(_0238_),
    .B1(net760),
    .Y(_0016_));
 sky130_fd_sc_hd__mux2_1 _8938_ (.A0(net774),
    .A1(_0223_),
    .S(_4164_),
    .X(_4091_));
 sky130_fd_sc_hd__clkbuf_1 _8939_ (.A(net775),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _8940_ (.A0(_0093_),
    .A1(_0771_),
    .S(_4242_),
    .X(_4092_));
 sky130_fd_sc_hd__clkbuf_1 _8941_ (.A(_4092_),
    .X(_0018_));
 sky130_fd_sc_hd__nand2_1 _8942_ (.A(_4242_),
    .B(net745),
    .Y(_4093_));
 sky130_fd_sc_hd__o21ai_1 _8943_ (.A1(_4242_),
    .A2(_0098_),
    .B1(net746),
    .Y(_0019_));
 sky130_fd_sc_hd__dfrtp_1 _8944_ (.CLK(clknet_2_0__leaf_clk_i),
    .D(_0024_),
    .RESET_B(net732),
    .Q(\arbiter.state[2][0] ));
 sky130_fd_sc_hd__dfrtp_1 _8945_ (.CLK(clknet_2_0__leaf_clk_i),
    .D(_0025_),
    .RESET_B(net732),
    .Q(\arbiter.state[2][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8946_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(_0002_),
    .RESET_B(net733),
    .Q(\arbiter.master_sel[2][0] ));
 sky130_fd_sc_hd__dfrtp_4 _8947_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(net755),
    .RESET_B(net733),
    .Q(\arbiter.master_sel[2][1] ));
 sky130_fd_sc_hd__dfrtp_4 _8948_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(_0004_),
    .RESET_B(net732),
    .Q(\arbiter.master_sel[3][0] ));
 sky130_fd_sc_hd__dfrtp_4 _8949_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(_0005_),
    .RESET_B(net732),
    .Q(\arbiter.master_sel[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8950_ (.CLK(clknet_2_3__leaf_clk_i),
    .D(_0006_),
    .RESET_B(net733),
    .Q(\arbiter.slave_sel[1][0] ));
 sky130_fd_sc_hd__dfrtp_4 _8951_ (.CLK(clknet_2_3__leaf_clk_i),
    .D(net758),
    .RESET_B(net733),
    .Q(\arbiter.slave_sel[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8952_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(_0022_),
    .RESET_B(net732),
    .Q(\arbiter.state[3][0] ));
 sky130_fd_sc_hd__dfrtp_4 _8953_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(_0023_),
    .RESET_B(net732),
    .Q(\arbiter.state[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8954_ (.CLK(clknet_2_3__leaf_clk_i),
    .D(_0008_),
    .RESET_B(net733),
    .Q(\arbiter.slave_sel[0][0] ));
 sky130_fd_sc_hd__dfrtp_1 _8955_ (.CLK(clknet_2_3__leaf_clk_i),
    .D(_0009_),
    .RESET_B(net733),
    .Q(\arbiter.slave_sel[0][1] ));
 sky130_fd_sc_hd__dfrtp_4 _8956_ (.CLK(clknet_2_2__leaf_clk_i),
    .D(_0010_),
    .RESET_B(net733),
    .Q(\arbiter.master_sel[1][0] ));
 sky130_fd_sc_hd__dfrtp_4 _8957_ (.CLK(clknet_2_2__leaf_clk_i),
    .D(net750),
    .RESET_B(net733),
    .Q(\arbiter.master_sel[1][1] ));
 sky130_fd_sc_hd__dfrtp_4 _8958_ (.CLK(clknet_2_0__leaf_clk_i),
    .D(_0012_),
    .RESET_B(net732),
    .Q(\arbiter.slave_sel[3][0] ));
 sky130_fd_sc_hd__dfrtp_4 _8959_ (.CLK(clknet_2_0__leaf_clk_i),
    .D(_0013_),
    .RESET_B(net732),
    .Q(\arbiter.slave_sel[3][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8960_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(net742),
    .RESET_B(net732),
    .Q(\arbiter.crossbar[3] ));
 sky130_fd_sc_hd__dfrtp_4 _8961_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(_0015_),
    .RESET_B(net732),
    .Q(\arbiter.crossbar[2] ));
 sky130_fd_sc_hd__dfstp_1 _8962_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(net739),
    .SET_B(net732),
    .Q(\arbiter.crossbar[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8963_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(net736),
    .RESET_B(net732),
    .Q(\arbiter.crossbar[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8964_ (.CLK(clknet_2_3__leaf_clk_i),
    .D(net761),
    .RESET_B(net733),
    .Q(\arbiter.master_sel[0][0] ));
 sky130_fd_sc_hd__dfrtp_4 _8965_ (.CLK(clknet_2_3__leaf_clk_i),
    .D(_0017_),
    .RESET_B(net733),
    .Q(\arbiter.master_sel[0][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8966_ (.CLK(clknet_2_3__leaf_clk_i),
    .D(_0020_),
    .RESET_B(net733),
    .Q(\arbiter.state[0][0] ));
 sky130_fd_sc_hd__dfrtp_4 _8967_ (.CLK(clknet_2_3__leaf_clk_i),
    .D(_0021_),
    .RESET_B(net229),
    .Q(\arbiter.state[0][1] ));
 sky130_fd_sc_hd__dfrtp_4 _8968_ (.CLK(clknet_2_0__leaf_clk_i),
    .D(_0032_),
    .RESET_B(net229),
    .Q(\arbiter.slave_handled[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8969_ (.CLK(clknet_2_0__leaf_clk_i),
    .D(_0033_),
    .RESET_B(net732),
    .Q(\arbiter.slave_handled[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8970_ (.CLK(clknet_2_0__leaf_clk_i),
    .D(_0034_),
    .RESET_B(net732),
    .Q(\arbiter.slave_handled[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8971_ (.CLK(clknet_2_0__leaf_clk_i),
    .D(_0035_),
    .RESET_B(net732),
    .Q(\arbiter.slave_handled[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8972_ (.CLK(clknet_2_2__leaf_clk_i),
    .D(_0028_),
    .RESET_B(net733),
    .Q(\arbiter.master_handled[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8973_ (.CLK(clknet_2_2__leaf_clk_i),
    .D(_0029_),
    .RESET_B(net733),
    .Q(\arbiter.master_handled[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8974_ (.CLK(clknet_2_2__leaf_clk_i),
    .D(_0030_),
    .RESET_B(net733),
    .Q(\arbiter.master_handled[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8975_ (.CLK(clknet_2_2__leaf_clk_i),
    .D(_0031_),
    .RESET_B(net733),
    .Q(\arbiter.master_handled[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8976_ (.CLK(clknet_2_2__leaf_clk_i),
    .D(_0026_),
    .RESET_B(net733),
    .Q(\arbiter.state[1][0] ));
 sky130_fd_sc_hd__dfrtp_4 _8977_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(_0027_),
    .RESET_B(net229),
    .Q(\arbiter.state[1][1] ));
 sky130_fd_sc_hd__dfrtp_1 _8978_ (.CLK(clknet_2_0__leaf_clk_i),
    .D(_0018_),
    .RESET_B(net732),
    .Q(\arbiter.slave_sel[2][0] ));
 sky130_fd_sc_hd__dfrtp_4 _8979_ (.CLK(clknet_2_1__leaf_clk_i),
    .D(net747),
    .RESET_B(net229),
    .Q(\arbiter.slave_sel[2][1] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk_i (.A(clk_i),
    .X(clknet_0_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_0__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_1__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_2__leaf_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk_i (.A(clknet_0_clk_i),
    .X(clknet_2_3__leaf_clk_i));
 sky130_fd_sc_hd__buf_6 fanout732 (.A(net229),
    .X(net732));
 sky130_fd_sc_hd__buf_6 fanout733 (.A(net229),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_2 hold1 (.A(\arbiter.crossbar[1] ),
    .X(net734));
 sky130_fd_sc_hd__clkbuf_4 hold10 (.A(\arbiter.crossbar[2] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(_4087_),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_4 hold12 (.A(\arbiter.slave_sel[2][1] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(_4093_),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(_0019_),
    .X(net747));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold15 (.A(\arbiter.master_sel[1][1] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(_4081_),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(_0011_),
    .X(net750));
 sky130_fd_sc_hd__buf_2 hold18 (.A(\arbiter.state[3][0] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(_0375_),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(_0404_),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_4 hold20 (.A(\arbiter.state[3][1] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\arbiter.master_sel[2][1] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(_0003_),
    .X(net755));
 sky130_fd_sc_hd__buf_2 hold23 (.A(\arbiter.slave_sel[1][1] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_4076_),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(_0007_),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\arbiter.master_sel[0][0] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_4090_),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(_0016_),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_2 hold29 (.A(\arbiter.state[2][0] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_0001_),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\arbiter.master_sel[3][1] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\arbiter.master_sel[3][0] ),
    .X(net764));
 sky130_fd_sc_hd__buf_2 hold32 (.A(\arbiter.state[1][0] ),
    .X(net765));
 sky130_fd_sc_hd__buf_1 hold33 (.A(\arbiter.master_handled[0] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\arbiter.master_handled[3] ),
    .X(net767));
 sky130_fd_sc_hd__clkdlybuf4s25_1 hold35 (.A(\arbiter.master_handled[2] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\arbiter.master_sel[1][0] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\arbiter.slave_sel[0][1] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(_4078_),
    .X(net771));
 sky130_fd_sc_hd__clkbuf_2 hold39 (.A(\arbiter.state[0][1] ),
    .X(net772));
 sky130_fd_sc_hd__buf_2 hold4 (.A(\arbiter.crossbar[0] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(_4112_),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\arbiter.master_sel[0][1] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_4091_),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\arbiter.master_sel[2][0] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\arbiter.slave_sel[3][1] ),
    .X(net777));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold45 (.A(\arbiter.state[0][0] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(_4159_),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(_0389_),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_0000_),
    .X(net739));
 sky130_fd_sc_hd__buf_2 hold7 (.A(\arbiter.crossbar[3] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(_4084_),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_0014_),
    .X(net742));
 sky130_fd_sc_hd__buf_2 input1 (.A(mports_i[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input10 (.A(mports_i[108]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input100 (.A(mports_i[18]),
    .X(net100));
 sky130_fd_sc_hd__buf_2 input101 (.A(mports_i[190]),
    .X(net101));
 sky130_fd_sc_hd__buf_2 input102 (.A(mports_i[191]),
    .X(net102));
 sky130_fd_sc_hd__buf_2 input103 (.A(mports_i[192]),
    .X(net103));
 sky130_fd_sc_hd__buf_2 input104 (.A(mports_i[193]),
    .X(net104));
 sky130_fd_sc_hd__buf_2 input105 (.A(mports_i[194]),
    .X(net105));
 sky130_fd_sc_hd__buf_2 input106 (.A(mports_i[195]),
    .X(net106));
 sky130_fd_sc_hd__clkbuf_2 input107 (.A(mports_i[196]),
    .X(net107));
 sky130_fd_sc_hd__buf_2 input108 (.A(mports_i[197]),
    .X(net108));
 sky130_fd_sc_hd__buf_2 input109 (.A(mports_i[198]),
    .X(net109));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(mports_i[109]),
    .X(net11));
 sky130_fd_sc_hd__buf_2 input110 (.A(mports_i[199]),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_4 input111 (.A(mports_i[19]),
    .X(net111));
 sky130_fd_sc_hd__buf_2 input112 (.A(mports_i[1]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 input113 (.A(mports_i[200]),
    .X(net113));
 sky130_fd_sc_hd__buf_2 input114 (.A(mports_i[201]),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_2 input115 (.A(mports_i[202]),
    .X(net115));
 sky130_fd_sc_hd__buf_2 input116 (.A(mports_i[203]),
    .X(net116));
 sky130_fd_sc_hd__buf_2 input117 (.A(mports_i[204]),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_2 input118 (.A(mports_i[205]),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 input119 (.A(mports_i[206]),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_4 input12 (.A(mports_i[10]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input120 (.A(mports_i[207]),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 input121 (.A(mports_i[208]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_2 input122 (.A(mports_i[209]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_4 input123 (.A(mports_i[20]),
    .X(net123));
 sky130_fd_sc_hd__buf_2 input124 (.A(mports_i[210]),
    .X(net124));
 sky130_fd_sc_hd__buf_2 input125 (.A(mports_i[211]),
    .X(net125));
 sky130_fd_sc_hd__buf_2 input126 (.A(mports_i[212]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_4 input127 (.A(mports_i[213]),
    .X(net127));
 sky130_fd_sc_hd__buf_2 input128 (.A(mports_i[214]),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_4 input129 (.A(mports_i[215]),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(mports_i[110]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input130 (.A(mports_i[216]),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_4 input131 (.A(mports_i[217]),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 input132 (.A(mports_i[218]),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 input133 (.A(mports_i[219]),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_4 input134 (.A(mports_i[21]),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_4 input135 (.A(mports_i[220]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_4 input136 (.A(mports_i[221]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_4 input137 (.A(mports_i[222]),
    .X(net137));
 sky130_fd_sc_hd__buf_6 input138 (.A(mports_i[223]),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_4 input139 (.A(mports_i[224]),
    .X(net139));
 sky130_fd_sc_hd__buf_2 input14 (.A(mports_i[111]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input140 (.A(mports_i[225]),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_4 input141 (.A(mports_i[226]),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_4 input142 (.A(mports_i[227]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_4 input143 (.A(mports_i[22]),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_4 input144 (.A(mports_i[23]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_4 input145 (.A(mports_i[24]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_4 input146 (.A(mports_i[25]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_4 input147 (.A(mports_i[26]),
    .X(net147));
 sky130_fd_sc_hd__buf_4 input148 (.A(mports_i[27]),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_4 input149 (.A(mports_i[28]),
    .X(net149));
 sky130_fd_sc_hd__buf_2 input15 (.A(mports_i[112]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input150 (.A(mports_i[29]),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_4 input151 (.A(mports_i[2]),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 input152 (.A(mports_i[30]),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 input153 (.A(mports_i[31]),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 input154 (.A(mports_i[32]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 input155 (.A(mports_i[33]),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_4 input156 (.A(mports_i[34]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 input157 (.A(mports_i[35]),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 input158 (.A(mports_i[36]),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_4 input159 (.A(mports_i[37]),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(mports_i[113]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 input160 (.A(mports_i[38]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_4 input161 (.A(mports_i[39]),
    .X(net161));
 sky130_fd_sc_hd__buf_2 input162 (.A(mports_i[3]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_4 input163 (.A(mports_i[40]),
    .X(net163));
 sky130_fd_sc_hd__buf_2 input164 (.A(mports_i[41]),
    .X(net164));
 sky130_fd_sc_hd__buf_2 input165 (.A(mports_i[42]),
    .X(net165));
 sky130_fd_sc_hd__buf_2 input166 (.A(mports_i[43]),
    .X(net166));
 sky130_fd_sc_hd__buf_2 input167 (.A(mports_i[44]),
    .X(net167));
 sky130_fd_sc_hd__buf_2 input168 (.A(mports_i[45]),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_2 input169 (.A(mports_i[46]),
    .X(net169));
 sky130_fd_sc_hd__buf_2 input17 (.A(mports_i[114]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input170 (.A(mports_i[47]),
    .X(net170));
 sky130_fd_sc_hd__dlymetal6s2s_1 input171 (.A(mports_i[48]),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_4 input172 (.A(mports_i[49]),
    .X(net172));
 sky130_fd_sc_hd__buf_2 input173 (.A(mports_i[4]),
    .X(net173));
 sky130_fd_sc_hd__buf_2 input174 (.A(mports_i[50]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_2 input175 (.A(mports_i[51]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(mports_i[52]),
    .X(net176));
 sky130_fd_sc_hd__dlymetal6s2s_1 input177 (.A(mports_i[53]),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_2 input178 (.A(mports_i[54]),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_2 input179 (.A(mports_i[55]),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(mports_i[115]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input180 (.A(mports_i[56]),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 input181 (.A(mports_i[57]),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_2 input182 (.A(mports_i[58]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 input183 (.A(mports_i[59]),
    .X(net183));
 sky130_fd_sc_hd__buf_2 input184 (.A(mports_i[5]),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 input185 (.A(mports_i[60]),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_2 input186 (.A(mports_i[61]),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_2 input187 (.A(mports_i[62]),
    .X(net187));
 sky130_fd_sc_hd__buf_2 input188 (.A(mports_i[63]),
    .X(net188));
 sky130_fd_sc_hd__buf_2 input189 (.A(mports_i[64]),
    .X(net189));
 sky130_fd_sc_hd__buf_2 input19 (.A(mports_i[116]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input190 (.A(mports_i[65]),
    .X(net190));
 sky130_fd_sc_hd__buf_2 input191 (.A(mports_i[66]),
    .X(net191));
 sky130_fd_sc_hd__buf_2 input192 (.A(mports_i[67]),
    .X(net192));
 sky130_fd_sc_hd__buf_2 input193 (.A(mports_i[68]),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 input194 (.A(mports_i[69]),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 input195 (.A(mports_i[6]),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 input196 (.A(mports_i[70]),
    .X(net196));
 sky130_fd_sc_hd__buf_2 input197 (.A(mports_i[71]),
    .X(net197));
 sky130_fd_sc_hd__buf_2 input198 (.A(mports_i[72]),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_4 input199 (.A(mports_i[73]),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(mports_i[100]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(mports_i[117]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input200 (.A(mports_i[74]),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 input201 (.A(mports_i[75]),
    .X(net201));
 sky130_fd_sc_hd__buf_2 input202 (.A(mports_i[76]),
    .X(net202));
 sky130_fd_sc_hd__buf_2 input203 (.A(mports_i[77]),
    .X(net203));
 sky130_fd_sc_hd__buf_2 input204 (.A(mports_i[78]),
    .X(net204));
 sky130_fd_sc_hd__buf_2 input205 (.A(mports_i[79]),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_4 input206 (.A(mports_i[7]),
    .X(net206));
 sky130_fd_sc_hd__buf_2 input207 (.A(mports_i[80]),
    .X(net207));
 sky130_fd_sc_hd__buf_2 input208 (.A(mports_i[81]),
    .X(net208));
 sky130_fd_sc_hd__buf_2 input209 (.A(mports_i[82]),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(mports_i[118]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input210 (.A(mports_i[83]),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 input211 (.A(mports_i[84]),
    .X(net211));
 sky130_fd_sc_hd__buf_2 input212 (.A(mports_i[85]),
    .X(net212));
 sky130_fd_sc_hd__buf_2 input213 (.A(mports_i[86]),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_4 input214 (.A(mports_i[87]),
    .X(net214));
 sky130_fd_sc_hd__clkbuf_4 input215 (.A(mports_i[88]),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_4 input216 (.A(mports_i[89]),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_4 input217 (.A(mports_i[8]),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_4 input218 (.A(mports_i[90]),
    .X(net218));
 sky130_fd_sc_hd__buf_2 input219 (.A(mports_i[91]),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(mports_i[119]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input220 (.A(mports_i[92]),
    .X(net220));
 sky130_fd_sc_hd__buf_2 input221 (.A(mports_i[93]),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 input222 (.A(mports_i[94]),
    .X(net222));
 sky130_fd_sc_hd__buf_2 input223 (.A(mports_i[95]),
    .X(net223));
 sky130_fd_sc_hd__buf_2 input224 (.A(mports_i[96]),
    .X(net224));
 sky130_fd_sc_hd__buf_2 input225 (.A(mports_i[97]),
    .X(net225));
 sky130_fd_sc_hd__buf_2 input226 (.A(mports_i[98]),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 input227 (.A(mports_i[99]),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_4 input228 (.A(mports_i[9]),
    .X(net228));
 sky130_fd_sc_hd__buf_8 input229 (.A(nrst_i),
    .X(net229));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(mports_i[11]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input230 (.A(sports_i[0]),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_8 input231 (.A(sports_i[100]),
    .X(net231));
 sky130_fd_sc_hd__clkbuf_4 input232 (.A(sports_i[101]),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_4 input233 (.A(sports_i[102]),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_4 input234 (.A(sports_i[103]),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_4 input235 (.A(sports_i[104]),
    .X(net235));
 sky130_fd_sc_hd__buf_4 input236 (.A(sports_i[105]),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_4 input237 (.A(sports_i[106]),
    .X(net237));
 sky130_fd_sc_hd__buf_1 input238 (.A(sports_i[107]),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_4 input239 (.A(sports_i[108]),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 input24 (.A(mports_i[120]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 input240 (.A(sports_i[109]),
    .X(net240));
 sky130_fd_sc_hd__dlymetal6s2s_1 input241 (.A(sports_i[10]),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_4 input242 (.A(sports_i[110]),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_4 input243 (.A(sports_i[111]),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_4 input244 (.A(sports_i[112]),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_4 input245 (.A(sports_i[113]),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_4 input246 (.A(sports_i[114]),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_4 input247 (.A(sports_i[115]),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_4 input248 (.A(sports_i[116]),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_4 input249 (.A(sports_i[117]),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_2 input25 (.A(mports_i[121]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_4 input250 (.A(sports_i[118]),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_4 input251 (.A(sports_i[119]),
    .X(net251));
 sky130_fd_sc_hd__buf_1 input252 (.A(sports_i[11]),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 input253 (.A(sports_i[120]),
    .X(net253));
 sky130_fd_sc_hd__clkbuf_4 input254 (.A(sports_i[121]),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_4 input255 (.A(sports_i[122]),
    .X(net255));
 sky130_fd_sc_hd__clkbuf_4 input256 (.A(sports_i[123]),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_4 input257 (.A(sports_i[124]),
    .X(net257));
 sky130_fd_sc_hd__buf_4 input258 (.A(sports_i[125]),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_4 input259 (.A(sports_i[126]),
    .X(net259));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(mports_i[122]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input260 (.A(sports_i[127]),
    .X(net260));
 sky130_fd_sc_hd__clkbuf_4 input261 (.A(sports_i[128]),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_4 input262 (.A(sports_i[129]),
    .X(net262));
 sky130_fd_sc_hd__dlymetal6s2s_1 input263 (.A(sports_i[12]),
    .X(net263));
 sky130_fd_sc_hd__clkbuf_4 input264 (.A(sports_i[130]),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_4 input265 (.A(sports_i[131]),
    .X(net265));
 sky130_fd_sc_hd__clkbuf_4 input266 (.A(sports_i[132]),
    .X(net266));
 sky130_fd_sc_hd__buf_4 input267 (.A(sports_i[133]),
    .X(net267));
 sky130_fd_sc_hd__clkbuf_2 input268 (.A(sports_i[134]),
    .X(net268));
 sky130_fd_sc_hd__clkbuf_4 input269 (.A(sports_i[135]),
    .X(net269));
 sky130_fd_sc_hd__buf_2 input27 (.A(mports_i[123]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input270 (.A(sports_i[13]),
    .X(net270));
 sky130_fd_sc_hd__buf_1 input271 (.A(sports_i[14]),
    .X(net271));
 sky130_fd_sc_hd__buf_1 input272 (.A(sports_i[15]),
    .X(net272));
 sky130_fd_sc_hd__buf_1 input273 (.A(sports_i[16]),
    .X(net273));
 sky130_fd_sc_hd__buf_1 input274 (.A(sports_i[17]),
    .X(net274));
 sky130_fd_sc_hd__buf_1 input275 (.A(sports_i[18]),
    .X(net275));
 sky130_fd_sc_hd__buf_1 input276 (.A(sports_i[19]),
    .X(net276));
 sky130_fd_sc_hd__buf_2 input277 (.A(sports_i[1]),
    .X(net277));
 sky130_fd_sc_hd__buf_1 input278 (.A(sports_i[20]),
    .X(net278));
 sky130_fd_sc_hd__buf_1 input279 (.A(sports_i[21]),
    .X(net279));
 sky130_fd_sc_hd__buf_2 input28 (.A(mports_i[124]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input280 (.A(sports_i[22]),
    .X(net280));
 sky130_fd_sc_hd__buf_1 input281 (.A(sports_i[23]),
    .X(net281));
 sky130_fd_sc_hd__buf_1 input282 (.A(sports_i[24]),
    .X(net282));
 sky130_fd_sc_hd__buf_1 input283 (.A(sports_i[25]),
    .X(net283));
 sky130_fd_sc_hd__buf_2 input284 (.A(sports_i[26]),
    .X(net284));
 sky130_fd_sc_hd__clkbuf_4 input285 (.A(sports_i[27]),
    .X(net285));
 sky130_fd_sc_hd__clkbuf_4 input286 (.A(sports_i[28]),
    .X(net286));
 sky130_fd_sc_hd__buf_2 input287 (.A(sports_i[29]),
    .X(net287));
 sky130_fd_sc_hd__buf_2 input288 (.A(sports_i[2]),
    .X(net288));
 sky130_fd_sc_hd__clkbuf_2 input289 (.A(sports_i[30]),
    .X(net289));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(mports_i[125]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 input290 (.A(sports_i[31]),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_8 input291 (.A(sports_i[32]),
    .X(net291));
 sky130_fd_sc_hd__buf_2 input292 (.A(sports_i[33]),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_4 input293 (.A(sports_i[34]),
    .X(net293));
 sky130_fd_sc_hd__buf_2 input294 (.A(sports_i[35]),
    .X(net294));
 sky130_fd_sc_hd__clkbuf_4 input295 (.A(sports_i[36]),
    .X(net295));
 sky130_fd_sc_hd__clkbuf_2 input296 (.A(sports_i[37]),
    .X(net296));
 sky130_fd_sc_hd__clkbuf_2 input297 (.A(sports_i[38]),
    .X(net297));
 sky130_fd_sc_hd__clkbuf_2 input298 (.A(sports_i[39]),
    .X(net298));
 sky130_fd_sc_hd__buf_2 input299 (.A(sports_i[3]),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(mports_i[101]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(mports_i[126]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input300 (.A(sports_i[40]),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_1 input301 (.A(sports_i[41]),
    .X(net301));
 sky130_fd_sc_hd__buf_1 input302 (.A(sports_i[42]),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_1 input303 (.A(sports_i[43]),
    .X(net303));
 sky130_fd_sc_hd__buf_1 input304 (.A(sports_i[44]),
    .X(net304));
 sky130_fd_sc_hd__buf_1 input305 (.A(sports_i[45]),
    .X(net305));
 sky130_fd_sc_hd__clkbuf_1 input306 (.A(sports_i[46]),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_1 input307 (.A(sports_i[47]),
    .X(net307));
 sky130_fd_sc_hd__buf_1 input308 (.A(sports_i[48]),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_1 input309 (.A(sports_i[49]),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(mports_i[127]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input310 (.A(sports_i[4]),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_1 input311 (.A(sports_i[50]),
    .X(net311));
 sky130_fd_sc_hd__clkbuf_1 input312 (.A(sports_i[51]),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_1 input313 (.A(sports_i[52]),
    .X(net313));
 sky130_fd_sc_hd__clkbuf_1 input314 (.A(sports_i[53]),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_1 input315 (.A(sports_i[54]),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_1 input316 (.A(sports_i[55]),
    .X(net316));
 sky130_fd_sc_hd__buf_1 input317 (.A(sports_i[56]),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_1 input318 (.A(sports_i[57]),
    .X(net318));
 sky130_fd_sc_hd__buf_1 input319 (.A(sports_i[58]),
    .X(net319));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(mports_i[128]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input320 (.A(sports_i[59]),
    .X(net320));
 sky130_fd_sc_hd__buf_2 input321 (.A(sports_i[5]),
    .X(net321));
 sky130_fd_sc_hd__buf_2 input322 (.A(sports_i[60]),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_2 input323 (.A(sports_i[61]),
    .X(net323));
 sky130_fd_sc_hd__buf_2 input324 (.A(sports_i[62]),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 input325 (.A(sports_i[63]),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_4 input326 (.A(sports_i[64]),
    .X(net326));
 sky130_fd_sc_hd__clkbuf_2 input327 (.A(sports_i[65]),
    .X(net327));
 sky130_fd_sc_hd__buf_4 input328 (.A(sports_i[66]),
    .X(net328));
 sky130_fd_sc_hd__buf_2 input329 (.A(sports_i[67]),
    .X(net329));
 sky130_fd_sc_hd__buf_2 input33 (.A(mports_i[129]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input330 (.A(sports_i[68]),
    .X(net330));
 sky130_fd_sc_hd__buf_2 input331 (.A(sports_i[69]),
    .X(net331));
 sky130_fd_sc_hd__buf_1 input332 (.A(sports_i[6]),
    .X(net332));
 sky130_fd_sc_hd__buf_4 input333 (.A(sports_i[70]),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_4 input334 (.A(sports_i[71]),
    .X(net334));
 sky130_fd_sc_hd__buf_2 input335 (.A(sports_i[72]),
    .X(net335));
 sky130_fd_sc_hd__buf_1 input336 (.A(sports_i[73]),
    .X(net336));
 sky130_fd_sc_hd__clkbuf_4 input337 (.A(sports_i[74]),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_1 input338 (.A(sports_i[75]),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_4 input339 (.A(sports_i[76]),
    .X(net339));
 sky130_fd_sc_hd__buf_2 input34 (.A(mports_i[12]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input340 (.A(sports_i[77]),
    .X(net340));
 sky130_fd_sc_hd__clkbuf_4 input341 (.A(sports_i[78]),
    .X(net341));
 sky130_fd_sc_hd__buf_2 input342 (.A(sports_i[79]),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 input343 (.A(sports_i[7]),
    .X(net343));
 sky130_fd_sc_hd__buf_2 input344 (.A(sports_i[80]),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_4 input345 (.A(sports_i[81]),
    .X(net345));
 sky130_fd_sc_hd__buf_2 input346 (.A(sports_i[82]),
    .X(net346));
 sky130_fd_sc_hd__clkbuf_4 input347 (.A(sports_i[83]),
    .X(net347));
 sky130_fd_sc_hd__buf_2 input348 (.A(sports_i[84]),
    .X(net348));
 sky130_fd_sc_hd__buf_2 input349 (.A(sports_i[85]),
    .X(net349));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(mports_i[130]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input350 (.A(sports_i[86]),
    .X(net350));
 sky130_fd_sc_hd__buf_2 input351 (.A(sports_i[87]),
    .X(net351));
 sky130_fd_sc_hd__clkbuf_4 input352 (.A(sports_i[88]),
    .X(net352));
 sky130_fd_sc_hd__buf_2 input353 (.A(sports_i[89]),
    .X(net353));
 sky130_fd_sc_hd__buf_1 input354 (.A(sports_i[8]),
    .X(net354));
 sky130_fd_sc_hd__buf_2 input355 (.A(sports_i[90]),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_4 input356 (.A(sports_i[91]),
    .X(net356));
 sky130_fd_sc_hd__clkbuf_4 input357 (.A(sports_i[92]),
    .X(net357));
 sky130_fd_sc_hd__buf_2 input358 (.A(sports_i[93]),
    .X(net358));
 sky130_fd_sc_hd__buf_2 input359 (.A(sports_i[94]),
    .X(net359));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(mports_i[131]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input360 (.A(sports_i[95]),
    .X(net360));
 sky130_fd_sc_hd__buf_2 input361 (.A(sports_i[96]),
    .X(net361));
 sky130_fd_sc_hd__buf_2 input362 (.A(sports_i[97]),
    .X(net362));
 sky130_fd_sc_hd__clkbuf_4 input363 (.A(sports_i[98]),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_4 input364 (.A(sports_i[99]),
    .X(net364));
 sky130_fd_sc_hd__buf_1 input365 (.A(sports_i[9]),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(mports_i[132]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(mports_i[133]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(mports_i[134]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(mports_i[102]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(mports_i[135]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(mports_i[136]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(mports_i[137]),
    .X(net42));
 sky130_fd_sc_hd__dlymetal6s2s_1 input43 (.A(mports_i[138]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(mports_i[139]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 input45 (.A(mports_i[13]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(mports_i[140]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(mports_i[141]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(mports_i[142]),
    .X(net48));
 sky130_fd_sc_hd__dlymetal6s2s_1 input49 (.A(mports_i[143]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(mports_i[103]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input50 (.A(mports_i[144]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_2 input51 (.A(mports_i[145]),
    .X(net51));
 sky130_fd_sc_hd__dlymetal6s2s_1 input52 (.A(mports_i[146]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(mports_i[147]),
    .X(net53));
 sky130_fd_sc_hd__dlymetal6s2s_1 input54 (.A(mports_i[148]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(mports_i[149]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 input56 (.A(mports_i[14]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(mports_i[150]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(mports_i[151]),
    .X(net58));
 sky130_fd_sc_hd__dlymetal6s2s_1 input59 (.A(mports_i[152]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(mports_i[104]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(mports_i[153]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 input61 (.A(mports_i[154]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(mports_i[155]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 input63 (.A(mports_i[156]),
    .X(net63));
 sky130_fd_sc_hd__buf_2 input64 (.A(mports_i[157]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 input65 (.A(mports_i[158]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 input66 (.A(mports_i[159]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_4 input67 (.A(mports_i[15]),
    .X(net67));
 sky130_fd_sc_hd__buf_2 input68 (.A(mports_i[160]),
    .X(net68));
 sky130_fd_sc_hd__buf_2 input69 (.A(mports_i[161]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(mports_i[105]),
    .X(net7));
 sky130_fd_sc_hd__buf_2 input70 (.A(mports_i[162]),
    .X(net70));
 sky130_fd_sc_hd__buf_2 input71 (.A(mports_i[163]),
    .X(net71));
 sky130_fd_sc_hd__buf_2 input72 (.A(mports_i[164]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 input73 (.A(mports_i[165]),
    .X(net73));
 sky130_fd_sc_hd__buf_6 input74 (.A(mports_i[166]),
    .X(net74));
 sky130_fd_sc_hd__buf_2 input75 (.A(mports_i[167]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_4 input76 (.A(mports_i[168]),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_4 input77 (.A(mports_i[169]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_4 input78 (.A(mports_i[16]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 input79 (.A(mports_i[170]),
    .X(net79));
 sky130_fd_sc_hd__buf_2 input8 (.A(mports_i[106]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_4 input80 (.A(mports_i[171]),
    .X(net80));
 sky130_fd_sc_hd__buf_2 input81 (.A(mports_i[172]),
    .X(net81));
 sky130_fd_sc_hd__buf_2 input82 (.A(mports_i[173]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_4 input83 (.A(mports_i[174]),
    .X(net83));
 sky130_fd_sc_hd__buf_2 input84 (.A(mports_i[175]),
    .X(net84));
 sky130_fd_sc_hd__buf_2 input85 (.A(mports_i[176]),
    .X(net85));
 sky130_fd_sc_hd__buf_2 input86 (.A(mports_i[177]),
    .X(net86));
 sky130_fd_sc_hd__buf_2 input87 (.A(mports_i[178]),
    .X(net87));
 sky130_fd_sc_hd__buf_2 input88 (.A(mports_i[179]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_4 input89 (.A(mports_i[17]),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(mports_i[107]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_4 input90 (.A(mports_i[180]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_4 input91 (.A(mports_i[181]),
    .X(net91));
 sky130_fd_sc_hd__buf_2 input92 (.A(mports_i[182]),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_4 input93 (.A(mports_i[183]),
    .X(net93));
 sky130_fd_sc_hd__buf_2 input94 (.A(mports_i[184]),
    .X(net94));
 sky130_fd_sc_hd__buf_2 input95 (.A(mports_i[185]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_4 input96 (.A(mports_i[186]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_2 input97 (.A(mports_i[187]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_2 input98 (.A(mports_i[188]),
    .X(net98));
 sky130_fd_sc_hd__buf_2 input99 (.A(mports_i[189]),
    .X(net99));
 sky130_fd_sc_hd__buf_12 output366 (.A(net366),
    .X(mports_o[0]));
 sky130_fd_sc_hd__buf_12 output367 (.A(net367),
    .X(mports_o[100]));
 sky130_fd_sc_hd__buf_12 output368 (.A(net368),
    .X(mports_o[101]));
 sky130_fd_sc_hd__buf_12 output369 (.A(net369),
    .X(mports_o[102]));
 sky130_fd_sc_hd__buf_12 output370 (.A(net370),
    .X(mports_o[103]));
 sky130_fd_sc_hd__buf_12 output371 (.A(net371),
    .X(mports_o[104]));
 sky130_fd_sc_hd__buf_12 output372 (.A(net372),
    .X(mports_o[105]));
 sky130_fd_sc_hd__buf_12 output373 (.A(net373),
    .X(mports_o[106]));
 sky130_fd_sc_hd__buf_12 output374 (.A(net374),
    .X(mports_o[107]));
 sky130_fd_sc_hd__buf_12 output375 (.A(net375),
    .X(mports_o[108]));
 sky130_fd_sc_hd__buf_12 output376 (.A(net376),
    .X(mports_o[109]));
 sky130_fd_sc_hd__buf_12 output377 (.A(net377),
    .X(mports_o[10]));
 sky130_fd_sc_hd__buf_12 output378 (.A(net378),
    .X(mports_o[110]));
 sky130_fd_sc_hd__buf_12 output379 (.A(net379),
    .X(mports_o[111]));
 sky130_fd_sc_hd__buf_12 output380 (.A(net380),
    .X(mports_o[112]));
 sky130_fd_sc_hd__buf_12 output381 (.A(net381),
    .X(mports_o[113]));
 sky130_fd_sc_hd__buf_12 output382 (.A(net382),
    .X(mports_o[114]));
 sky130_fd_sc_hd__buf_12 output383 (.A(net383),
    .X(mports_o[115]));
 sky130_fd_sc_hd__buf_12 output384 (.A(net384),
    .X(mports_o[116]));
 sky130_fd_sc_hd__buf_12 output385 (.A(net385),
    .X(mports_o[117]));
 sky130_fd_sc_hd__buf_12 output386 (.A(net386),
    .X(mports_o[118]));
 sky130_fd_sc_hd__buf_12 output387 (.A(net387),
    .X(mports_o[119]));
 sky130_fd_sc_hd__buf_12 output388 (.A(net388),
    .X(mports_o[11]));
 sky130_fd_sc_hd__buf_12 output389 (.A(net389),
    .X(mports_o[120]));
 sky130_fd_sc_hd__buf_12 output390 (.A(net390),
    .X(mports_o[121]));
 sky130_fd_sc_hd__buf_12 output391 (.A(net391),
    .X(mports_o[122]));
 sky130_fd_sc_hd__buf_12 output392 (.A(net392),
    .X(mports_o[123]));
 sky130_fd_sc_hd__buf_12 output393 (.A(net393),
    .X(mports_o[124]));
 sky130_fd_sc_hd__buf_12 output394 (.A(net394),
    .X(mports_o[125]));
 sky130_fd_sc_hd__buf_12 output395 (.A(net395),
    .X(mports_o[126]));
 sky130_fd_sc_hd__buf_12 output396 (.A(net396),
    .X(mports_o[127]));
 sky130_fd_sc_hd__buf_12 output397 (.A(net397),
    .X(mports_o[128]));
 sky130_fd_sc_hd__buf_12 output398 (.A(net398),
    .X(mports_o[129]));
 sky130_fd_sc_hd__buf_12 output399 (.A(net399),
    .X(mports_o[12]));
 sky130_fd_sc_hd__buf_12 output400 (.A(net400),
    .X(mports_o[130]));
 sky130_fd_sc_hd__buf_12 output401 (.A(net401),
    .X(mports_o[131]));
 sky130_fd_sc_hd__buf_12 output402 (.A(net402),
    .X(mports_o[132]));
 sky130_fd_sc_hd__buf_12 output403 (.A(net403),
    .X(mports_o[133]));
 sky130_fd_sc_hd__buf_12 output404 (.A(net404),
    .X(mports_o[134]));
 sky130_fd_sc_hd__buf_12 output405 (.A(net405),
    .X(mports_o[135]));
 sky130_fd_sc_hd__buf_12 output406 (.A(net406),
    .X(mports_o[13]));
 sky130_fd_sc_hd__buf_12 output407 (.A(net407),
    .X(mports_o[14]));
 sky130_fd_sc_hd__buf_12 output408 (.A(net408),
    .X(mports_o[15]));
 sky130_fd_sc_hd__buf_12 output409 (.A(net409),
    .X(mports_o[16]));
 sky130_fd_sc_hd__buf_12 output410 (.A(net410),
    .X(mports_o[17]));
 sky130_fd_sc_hd__buf_12 output411 (.A(net411),
    .X(mports_o[18]));
 sky130_fd_sc_hd__buf_12 output412 (.A(net412),
    .X(mports_o[19]));
 sky130_fd_sc_hd__buf_12 output413 (.A(net413),
    .X(mports_o[1]));
 sky130_fd_sc_hd__buf_12 output414 (.A(net414),
    .X(mports_o[20]));
 sky130_fd_sc_hd__buf_12 output415 (.A(net415),
    .X(mports_o[21]));
 sky130_fd_sc_hd__buf_12 output416 (.A(net416),
    .X(mports_o[22]));
 sky130_fd_sc_hd__buf_12 output417 (.A(net417),
    .X(mports_o[23]));
 sky130_fd_sc_hd__buf_12 output418 (.A(net418),
    .X(mports_o[24]));
 sky130_fd_sc_hd__buf_12 output419 (.A(net419),
    .X(mports_o[25]));
 sky130_fd_sc_hd__buf_12 output420 (.A(net420),
    .X(mports_o[26]));
 sky130_fd_sc_hd__buf_12 output421 (.A(net421),
    .X(mports_o[27]));
 sky130_fd_sc_hd__buf_12 output422 (.A(net422),
    .X(mports_o[28]));
 sky130_fd_sc_hd__buf_12 output423 (.A(net423),
    .X(mports_o[29]));
 sky130_fd_sc_hd__buf_12 output424 (.A(net424),
    .X(mports_o[2]));
 sky130_fd_sc_hd__buf_12 output425 (.A(net425),
    .X(mports_o[30]));
 sky130_fd_sc_hd__buf_12 output426 (.A(net426),
    .X(mports_o[31]));
 sky130_fd_sc_hd__buf_12 output427 (.A(net427),
    .X(mports_o[32]));
 sky130_fd_sc_hd__buf_12 output428 (.A(net428),
    .X(mports_o[33]));
 sky130_fd_sc_hd__buf_12 output429 (.A(net429),
    .X(mports_o[34]));
 sky130_fd_sc_hd__buf_12 output430 (.A(net430),
    .X(mports_o[35]));
 sky130_fd_sc_hd__buf_12 output431 (.A(net431),
    .X(mports_o[36]));
 sky130_fd_sc_hd__buf_12 output432 (.A(net432),
    .X(mports_o[37]));
 sky130_fd_sc_hd__buf_12 output433 (.A(net433),
    .X(mports_o[38]));
 sky130_fd_sc_hd__buf_12 output434 (.A(net434),
    .X(mports_o[39]));
 sky130_fd_sc_hd__buf_12 output435 (.A(net435),
    .X(mports_o[3]));
 sky130_fd_sc_hd__buf_12 output436 (.A(net436),
    .X(mports_o[40]));
 sky130_fd_sc_hd__buf_12 output437 (.A(net437),
    .X(mports_o[41]));
 sky130_fd_sc_hd__buf_12 output438 (.A(net438),
    .X(mports_o[42]));
 sky130_fd_sc_hd__buf_12 output439 (.A(net439),
    .X(mports_o[43]));
 sky130_fd_sc_hd__buf_12 output440 (.A(net440),
    .X(mports_o[44]));
 sky130_fd_sc_hd__buf_12 output441 (.A(net441),
    .X(mports_o[45]));
 sky130_fd_sc_hd__buf_12 output442 (.A(net442),
    .X(mports_o[46]));
 sky130_fd_sc_hd__buf_12 output443 (.A(net443),
    .X(mports_o[47]));
 sky130_fd_sc_hd__buf_12 output444 (.A(net444),
    .X(mports_o[48]));
 sky130_fd_sc_hd__buf_12 output445 (.A(net445),
    .X(mports_o[49]));
 sky130_fd_sc_hd__buf_12 output446 (.A(net446),
    .X(mports_o[4]));
 sky130_fd_sc_hd__buf_12 output447 (.A(net447),
    .X(mports_o[50]));
 sky130_fd_sc_hd__buf_12 output448 (.A(net448),
    .X(mports_o[51]));
 sky130_fd_sc_hd__buf_12 output449 (.A(net449),
    .X(mports_o[52]));
 sky130_fd_sc_hd__buf_12 output450 (.A(net450),
    .X(mports_o[53]));
 sky130_fd_sc_hd__buf_12 output451 (.A(net451),
    .X(mports_o[54]));
 sky130_fd_sc_hd__buf_12 output452 (.A(net452),
    .X(mports_o[55]));
 sky130_fd_sc_hd__buf_12 output453 (.A(net453),
    .X(mports_o[56]));
 sky130_fd_sc_hd__buf_12 output454 (.A(net454),
    .X(mports_o[57]));
 sky130_fd_sc_hd__buf_12 output455 (.A(net455),
    .X(mports_o[58]));
 sky130_fd_sc_hd__buf_12 output456 (.A(net456),
    .X(mports_o[59]));
 sky130_fd_sc_hd__buf_12 output457 (.A(net457),
    .X(mports_o[5]));
 sky130_fd_sc_hd__buf_12 output458 (.A(net458),
    .X(mports_o[60]));
 sky130_fd_sc_hd__buf_12 output459 (.A(net459),
    .X(mports_o[61]));
 sky130_fd_sc_hd__buf_12 output460 (.A(net460),
    .X(mports_o[62]));
 sky130_fd_sc_hd__buf_12 output461 (.A(net461),
    .X(mports_o[63]));
 sky130_fd_sc_hd__buf_12 output462 (.A(net462),
    .X(mports_o[64]));
 sky130_fd_sc_hd__buf_12 output463 (.A(net463),
    .X(mports_o[65]));
 sky130_fd_sc_hd__buf_12 output464 (.A(net464),
    .X(mports_o[66]));
 sky130_fd_sc_hd__buf_12 output465 (.A(net465),
    .X(mports_o[67]));
 sky130_fd_sc_hd__buf_12 output466 (.A(net466),
    .X(mports_o[68]));
 sky130_fd_sc_hd__buf_12 output467 (.A(net467),
    .X(mports_o[69]));
 sky130_fd_sc_hd__buf_12 output468 (.A(net468),
    .X(mports_o[6]));
 sky130_fd_sc_hd__buf_12 output469 (.A(net469),
    .X(mports_o[70]));
 sky130_fd_sc_hd__buf_12 output470 (.A(net470),
    .X(mports_o[71]));
 sky130_fd_sc_hd__buf_12 output471 (.A(net471),
    .X(mports_o[72]));
 sky130_fd_sc_hd__buf_12 output472 (.A(net472),
    .X(mports_o[73]));
 sky130_fd_sc_hd__buf_12 output473 (.A(net473),
    .X(mports_o[74]));
 sky130_fd_sc_hd__buf_12 output474 (.A(net474),
    .X(mports_o[75]));
 sky130_fd_sc_hd__buf_12 output475 (.A(net475),
    .X(mports_o[76]));
 sky130_fd_sc_hd__buf_12 output476 (.A(net476),
    .X(mports_o[77]));
 sky130_fd_sc_hd__buf_12 output477 (.A(net477),
    .X(mports_o[78]));
 sky130_fd_sc_hd__buf_12 output478 (.A(net478),
    .X(mports_o[79]));
 sky130_fd_sc_hd__buf_12 output479 (.A(net479),
    .X(mports_o[7]));
 sky130_fd_sc_hd__buf_12 output480 (.A(net480),
    .X(mports_o[80]));
 sky130_fd_sc_hd__buf_12 output481 (.A(net481),
    .X(mports_o[81]));
 sky130_fd_sc_hd__buf_12 output482 (.A(net482),
    .X(mports_o[82]));
 sky130_fd_sc_hd__buf_12 output483 (.A(net483),
    .X(mports_o[83]));
 sky130_fd_sc_hd__buf_12 output484 (.A(net484),
    .X(mports_o[84]));
 sky130_fd_sc_hd__buf_12 output485 (.A(net485),
    .X(mports_o[85]));
 sky130_fd_sc_hd__buf_12 output486 (.A(net486),
    .X(mports_o[86]));
 sky130_fd_sc_hd__buf_12 output487 (.A(net487),
    .X(mports_o[87]));
 sky130_fd_sc_hd__buf_12 output488 (.A(net488),
    .X(mports_o[88]));
 sky130_fd_sc_hd__buf_12 output489 (.A(net489),
    .X(mports_o[89]));
 sky130_fd_sc_hd__buf_12 output490 (.A(net490),
    .X(mports_o[8]));
 sky130_fd_sc_hd__buf_12 output491 (.A(net491),
    .X(mports_o[90]));
 sky130_fd_sc_hd__buf_12 output492 (.A(net492),
    .X(mports_o[91]));
 sky130_fd_sc_hd__buf_12 output493 (.A(net493),
    .X(mports_o[92]));
 sky130_fd_sc_hd__buf_12 output494 (.A(net494),
    .X(mports_o[93]));
 sky130_fd_sc_hd__buf_12 output495 (.A(net495),
    .X(mports_o[94]));
 sky130_fd_sc_hd__buf_12 output496 (.A(net496),
    .X(mports_o[95]));
 sky130_fd_sc_hd__buf_12 output497 (.A(net497),
    .X(mports_o[96]));
 sky130_fd_sc_hd__buf_12 output498 (.A(net498),
    .X(mports_o[97]));
 sky130_fd_sc_hd__buf_12 output499 (.A(net499),
    .X(mports_o[98]));
 sky130_fd_sc_hd__buf_12 output500 (.A(net500),
    .X(mports_o[99]));
 sky130_fd_sc_hd__buf_12 output501 (.A(net501),
    .X(mports_o[9]));
 sky130_fd_sc_hd__buf_12 output502 (.A(net502),
    .X(sports_o[0]));
 sky130_fd_sc_hd__buf_12 output503 (.A(net503),
    .X(sports_o[100]));
 sky130_fd_sc_hd__buf_12 output504 (.A(net504),
    .X(sports_o[101]));
 sky130_fd_sc_hd__buf_12 output505 (.A(net505),
    .X(sports_o[102]));
 sky130_fd_sc_hd__buf_12 output506 (.A(net506),
    .X(sports_o[103]));
 sky130_fd_sc_hd__buf_12 output507 (.A(net507),
    .X(sports_o[104]));
 sky130_fd_sc_hd__buf_12 output508 (.A(net508),
    .X(sports_o[105]));
 sky130_fd_sc_hd__buf_12 output509 (.A(net509),
    .X(sports_o[106]));
 sky130_fd_sc_hd__buf_12 output510 (.A(net510),
    .X(sports_o[107]));
 sky130_fd_sc_hd__buf_12 output511 (.A(net511),
    .X(sports_o[108]));
 sky130_fd_sc_hd__buf_12 output512 (.A(net512),
    .X(sports_o[109]));
 sky130_fd_sc_hd__buf_12 output513 (.A(net513),
    .X(sports_o[10]));
 sky130_fd_sc_hd__buf_12 output514 (.A(net514),
    .X(sports_o[110]));
 sky130_fd_sc_hd__buf_12 output515 (.A(net515),
    .X(sports_o[111]));
 sky130_fd_sc_hd__buf_12 output516 (.A(net516),
    .X(sports_o[112]));
 sky130_fd_sc_hd__buf_12 output517 (.A(net517),
    .X(sports_o[113]));
 sky130_fd_sc_hd__buf_12 output518 (.A(net518),
    .X(sports_o[114]));
 sky130_fd_sc_hd__buf_12 output519 (.A(net519),
    .X(sports_o[115]));
 sky130_fd_sc_hd__buf_12 output520 (.A(net520),
    .X(sports_o[116]));
 sky130_fd_sc_hd__buf_12 output521 (.A(net521),
    .X(sports_o[117]));
 sky130_fd_sc_hd__buf_12 output522 (.A(net522),
    .X(sports_o[118]));
 sky130_fd_sc_hd__buf_12 output523 (.A(net523),
    .X(sports_o[119]));
 sky130_fd_sc_hd__buf_12 output524 (.A(net524),
    .X(sports_o[11]));
 sky130_fd_sc_hd__buf_12 output525 (.A(net525),
    .X(sports_o[120]));
 sky130_fd_sc_hd__buf_12 output526 (.A(net526),
    .X(sports_o[121]));
 sky130_fd_sc_hd__buf_12 output527 (.A(net527),
    .X(sports_o[122]));
 sky130_fd_sc_hd__buf_12 output528 (.A(net528),
    .X(sports_o[123]));
 sky130_fd_sc_hd__buf_12 output529 (.A(net529),
    .X(sports_o[124]));
 sky130_fd_sc_hd__buf_12 output530 (.A(net530),
    .X(sports_o[125]));
 sky130_fd_sc_hd__buf_12 output531 (.A(net531),
    .X(sports_o[126]));
 sky130_fd_sc_hd__buf_12 output532 (.A(net532),
    .X(sports_o[127]));
 sky130_fd_sc_hd__buf_12 output533 (.A(net533),
    .X(sports_o[128]));
 sky130_fd_sc_hd__buf_12 output534 (.A(net534),
    .X(sports_o[129]));
 sky130_fd_sc_hd__buf_12 output535 (.A(net535),
    .X(sports_o[12]));
 sky130_fd_sc_hd__buf_12 output536 (.A(net536),
    .X(sports_o[130]));
 sky130_fd_sc_hd__buf_12 output537 (.A(net537),
    .X(sports_o[131]));
 sky130_fd_sc_hd__buf_12 output538 (.A(net538),
    .X(sports_o[132]));
 sky130_fd_sc_hd__buf_12 output539 (.A(net539),
    .X(sports_o[133]));
 sky130_fd_sc_hd__buf_12 output540 (.A(net540),
    .X(sports_o[134]));
 sky130_fd_sc_hd__buf_12 output541 (.A(net541),
    .X(sports_o[135]));
 sky130_fd_sc_hd__buf_12 output542 (.A(net542),
    .X(sports_o[136]));
 sky130_fd_sc_hd__buf_12 output543 (.A(net543),
    .X(sports_o[137]));
 sky130_fd_sc_hd__buf_12 output544 (.A(net544),
    .X(sports_o[138]));
 sky130_fd_sc_hd__buf_12 output545 (.A(net545),
    .X(sports_o[139]));
 sky130_fd_sc_hd__buf_12 output546 (.A(net546),
    .X(sports_o[13]));
 sky130_fd_sc_hd__buf_12 output547 (.A(net547),
    .X(sports_o[140]));
 sky130_fd_sc_hd__buf_12 output548 (.A(net548),
    .X(sports_o[141]));
 sky130_fd_sc_hd__buf_12 output549 (.A(net549),
    .X(sports_o[142]));
 sky130_fd_sc_hd__buf_12 output550 (.A(net550),
    .X(sports_o[143]));
 sky130_fd_sc_hd__buf_12 output551 (.A(net551),
    .X(sports_o[144]));
 sky130_fd_sc_hd__buf_12 output552 (.A(net552),
    .X(sports_o[145]));
 sky130_fd_sc_hd__buf_12 output553 (.A(net553),
    .X(sports_o[146]));
 sky130_fd_sc_hd__buf_12 output554 (.A(net554),
    .X(sports_o[147]));
 sky130_fd_sc_hd__buf_12 output555 (.A(net555),
    .X(sports_o[148]));
 sky130_fd_sc_hd__buf_12 output556 (.A(net556),
    .X(sports_o[149]));
 sky130_fd_sc_hd__buf_12 output557 (.A(net557),
    .X(sports_o[14]));
 sky130_fd_sc_hd__buf_12 output558 (.A(net558),
    .X(sports_o[150]));
 sky130_fd_sc_hd__buf_12 output559 (.A(net559),
    .X(sports_o[151]));
 sky130_fd_sc_hd__buf_12 output560 (.A(net560),
    .X(sports_o[152]));
 sky130_fd_sc_hd__buf_12 output561 (.A(net561),
    .X(sports_o[153]));
 sky130_fd_sc_hd__buf_12 output562 (.A(net562),
    .X(sports_o[154]));
 sky130_fd_sc_hd__buf_12 output563 (.A(net563),
    .X(sports_o[155]));
 sky130_fd_sc_hd__buf_12 output564 (.A(net564),
    .X(sports_o[156]));
 sky130_fd_sc_hd__buf_12 output565 (.A(net565),
    .X(sports_o[157]));
 sky130_fd_sc_hd__buf_12 output566 (.A(net566),
    .X(sports_o[158]));
 sky130_fd_sc_hd__buf_12 output567 (.A(net567),
    .X(sports_o[159]));
 sky130_fd_sc_hd__buf_12 output568 (.A(net568),
    .X(sports_o[15]));
 sky130_fd_sc_hd__buf_12 output569 (.A(net569),
    .X(sports_o[160]));
 sky130_fd_sc_hd__buf_12 output570 (.A(net570),
    .X(sports_o[161]));
 sky130_fd_sc_hd__buf_12 output571 (.A(net571),
    .X(sports_o[162]));
 sky130_fd_sc_hd__buf_12 output572 (.A(net572),
    .X(sports_o[163]));
 sky130_fd_sc_hd__buf_12 output573 (.A(net573),
    .X(sports_o[164]));
 sky130_fd_sc_hd__buf_12 output574 (.A(net574),
    .X(sports_o[165]));
 sky130_fd_sc_hd__buf_12 output575 (.A(net575),
    .X(sports_o[166]));
 sky130_fd_sc_hd__buf_12 output576 (.A(net576),
    .X(sports_o[167]));
 sky130_fd_sc_hd__buf_12 output577 (.A(net577),
    .X(sports_o[168]));
 sky130_fd_sc_hd__buf_12 output578 (.A(net578),
    .X(sports_o[169]));
 sky130_fd_sc_hd__buf_12 output579 (.A(net579),
    .X(sports_o[16]));
 sky130_fd_sc_hd__buf_12 output580 (.A(net580),
    .X(sports_o[170]));
 sky130_fd_sc_hd__buf_12 output581 (.A(net581),
    .X(sports_o[171]));
 sky130_fd_sc_hd__buf_12 output582 (.A(net582),
    .X(sports_o[172]));
 sky130_fd_sc_hd__buf_12 output583 (.A(net583),
    .X(sports_o[173]));
 sky130_fd_sc_hd__buf_12 output584 (.A(net584),
    .X(sports_o[174]));
 sky130_fd_sc_hd__buf_12 output585 (.A(net585),
    .X(sports_o[175]));
 sky130_fd_sc_hd__buf_12 output586 (.A(net586),
    .X(sports_o[176]));
 sky130_fd_sc_hd__buf_12 output587 (.A(net587),
    .X(sports_o[177]));
 sky130_fd_sc_hd__buf_12 output588 (.A(net588),
    .X(sports_o[178]));
 sky130_fd_sc_hd__buf_12 output589 (.A(net589),
    .X(sports_o[179]));
 sky130_fd_sc_hd__buf_12 output590 (.A(net590),
    .X(sports_o[17]));
 sky130_fd_sc_hd__buf_12 output591 (.A(net591),
    .X(sports_o[180]));
 sky130_fd_sc_hd__buf_12 output592 (.A(net592),
    .X(sports_o[181]));
 sky130_fd_sc_hd__buf_12 output593 (.A(net593),
    .X(sports_o[182]));
 sky130_fd_sc_hd__buf_12 output594 (.A(net594),
    .X(sports_o[183]));
 sky130_fd_sc_hd__buf_12 output595 (.A(net595),
    .X(sports_o[184]));
 sky130_fd_sc_hd__buf_12 output596 (.A(net596),
    .X(sports_o[185]));
 sky130_fd_sc_hd__buf_12 output597 (.A(net597),
    .X(sports_o[186]));
 sky130_fd_sc_hd__buf_12 output598 (.A(net598),
    .X(sports_o[187]));
 sky130_fd_sc_hd__buf_12 output599 (.A(net599),
    .X(sports_o[188]));
 sky130_fd_sc_hd__buf_12 output600 (.A(net600),
    .X(sports_o[189]));
 sky130_fd_sc_hd__buf_12 output601 (.A(net601),
    .X(sports_o[18]));
 sky130_fd_sc_hd__buf_12 output602 (.A(net602),
    .X(sports_o[190]));
 sky130_fd_sc_hd__buf_12 output603 (.A(net603),
    .X(sports_o[191]));
 sky130_fd_sc_hd__buf_12 output604 (.A(net604),
    .X(sports_o[192]));
 sky130_fd_sc_hd__buf_12 output605 (.A(net605),
    .X(sports_o[193]));
 sky130_fd_sc_hd__buf_12 output606 (.A(net606),
    .X(sports_o[194]));
 sky130_fd_sc_hd__buf_12 output607 (.A(net607),
    .X(sports_o[195]));
 sky130_fd_sc_hd__buf_12 output608 (.A(net608),
    .X(sports_o[196]));
 sky130_fd_sc_hd__buf_12 output609 (.A(net609),
    .X(sports_o[197]));
 sky130_fd_sc_hd__buf_12 output610 (.A(net610),
    .X(sports_o[198]));
 sky130_fd_sc_hd__buf_12 output611 (.A(net611),
    .X(sports_o[199]));
 sky130_fd_sc_hd__buf_12 output612 (.A(net612),
    .X(sports_o[19]));
 sky130_fd_sc_hd__buf_12 output613 (.A(net613),
    .X(sports_o[1]));
 sky130_fd_sc_hd__buf_12 output614 (.A(net614),
    .X(sports_o[200]));
 sky130_fd_sc_hd__buf_12 output615 (.A(net615),
    .X(sports_o[201]));
 sky130_fd_sc_hd__buf_12 output616 (.A(net616),
    .X(sports_o[202]));
 sky130_fd_sc_hd__buf_12 output617 (.A(net617),
    .X(sports_o[203]));
 sky130_fd_sc_hd__buf_12 output618 (.A(net618),
    .X(sports_o[204]));
 sky130_fd_sc_hd__buf_12 output619 (.A(net619),
    .X(sports_o[205]));
 sky130_fd_sc_hd__buf_12 output620 (.A(net620),
    .X(sports_o[206]));
 sky130_fd_sc_hd__buf_12 output621 (.A(net621),
    .X(sports_o[207]));
 sky130_fd_sc_hd__buf_12 output622 (.A(net622),
    .X(sports_o[208]));
 sky130_fd_sc_hd__buf_12 output623 (.A(net623),
    .X(sports_o[209]));
 sky130_fd_sc_hd__buf_12 output624 (.A(net624),
    .X(sports_o[20]));
 sky130_fd_sc_hd__buf_12 output625 (.A(net625),
    .X(sports_o[210]));
 sky130_fd_sc_hd__buf_12 output626 (.A(net626),
    .X(sports_o[211]));
 sky130_fd_sc_hd__buf_12 output627 (.A(net627),
    .X(sports_o[212]));
 sky130_fd_sc_hd__buf_12 output628 (.A(net628),
    .X(sports_o[213]));
 sky130_fd_sc_hd__buf_12 output629 (.A(net629),
    .X(sports_o[214]));
 sky130_fd_sc_hd__buf_12 output630 (.A(net630),
    .X(sports_o[215]));
 sky130_fd_sc_hd__buf_12 output631 (.A(net631),
    .X(sports_o[216]));
 sky130_fd_sc_hd__buf_12 output632 (.A(net632),
    .X(sports_o[217]));
 sky130_fd_sc_hd__buf_12 output633 (.A(net633),
    .X(sports_o[218]));
 sky130_fd_sc_hd__buf_12 output634 (.A(net634),
    .X(sports_o[219]));
 sky130_fd_sc_hd__buf_12 output635 (.A(net635),
    .X(sports_o[21]));
 sky130_fd_sc_hd__buf_12 output636 (.A(net636),
    .X(sports_o[220]));
 sky130_fd_sc_hd__buf_12 output637 (.A(net637),
    .X(sports_o[221]));
 sky130_fd_sc_hd__buf_12 output638 (.A(net638),
    .X(sports_o[222]));
 sky130_fd_sc_hd__buf_12 output639 (.A(net639),
    .X(sports_o[223]));
 sky130_fd_sc_hd__buf_12 output640 (.A(net640),
    .X(sports_o[224]));
 sky130_fd_sc_hd__buf_12 output641 (.A(net641),
    .X(sports_o[225]));
 sky130_fd_sc_hd__buf_12 output642 (.A(net642),
    .X(sports_o[226]));
 sky130_fd_sc_hd__buf_12 output643 (.A(net643),
    .X(sports_o[227]));
 sky130_fd_sc_hd__buf_12 output644 (.A(net644),
    .X(sports_o[22]));
 sky130_fd_sc_hd__buf_12 output645 (.A(net645),
    .X(sports_o[23]));
 sky130_fd_sc_hd__buf_12 output646 (.A(net646),
    .X(sports_o[24]));
 sky130_fd_sc_hd__buf_12 output647 (.A(net647),
    .X(sports_o[25]));
 sky130_fd_sc_hd__buf_12 output648 (.A(net648),
    .X(sports_o[26]));
 sky130_fd_sc_hd__buf_12 output649 (.A(net649),
    .X(sports_o[27]));
 sky130_fd_sc_hd__buf_12 output650 (.A(net650),
    .X(sports_o[28]));
 sky130_fd_sc_hd__buf_12 output651 (.A(net651),
    .X(sports_o[29]));
 sky130_fd_sc_hd__buf_12 output652 (.A(net652),
    .X(sports_o[2]));
 sky130_fd_sc_hd__buf_12 output653 (.A(net653),
    .X(sports_o[30]));
 sky130_fd_sc_hd__buf_12 output654 (.A(net654),
    .X(sports_o[31]));
 sky130_fd_sc_hd__buf_12 output655 (.A(net655),
    .X(sports_o[32]));
 sky130_fd_sc_hd__buf_12 output656 (.A(net656),
    .X(sports_o[33]));
 sky130_fd_sc_hd__buf_12 output657 (.A(net657),
    .X(sports_o[34]));
 sky130_fd_sc_hd__buf_12 output658 (.A(net658),
    .X(sports_o[35]));
 sky130_fd_sc_hd__buf_12 output659 (.A(net659),
    .X(sports_o[36]));
 sky130_fd_sc_hd__buf_12 output660 (.A(net660),
    .X(sports_o[37]));
 sky130_fd_sc_hd__buf_12 output661 (.A(net661),
    .X(sports_o[38]));
 sky130_fd_sc_hd__buf_12 output662 (.A(net662),
    .X(sports_o[39]));
 sky130_fd_sc_hd__buf_12 output663 (.A(net663),
    .X(sports_o[3]));
 sky130_fd_sc_hd__buf_12 output664 (.A(net664),
    .X(sports_o[40]));
 sky130_fd_sc_hd__buf_12 output665 (.A(net665),
    .X(sports_o[41]));
 sky130_fd_sc_hd__buf_12 output666 (.A(net666),
    .X(sports_o[42]));
 sky130_fd_sc_hd__buf_12 output667 (.A(net667),
    .X(sports_o[43]));
 sky130_fd_sc_hd__buf_12 output668 (.A(net668),
    .X(sports_o[44]));
 sky130_fd_sc_hd__buf_12 output669 (.A(net669),
    .X(sports_o[45]));
 sky130_fd_sc_hd__buf_12 output670 (.A(net670),
    .X(sports_o[46]));
 sky130_fd_sc_hd__buf_12 output671 (.A(net671),
    .X(sports_o[47]));
 sky130_fd_sc_hd__buf_12 output672 (.A(net672),
    .X(sports_o[48]));
 sky130_fd_sc_hd__buf_12 output673 (.A(net673),
    .X(sports_o[49]));
 sky130_fd_sc_hd__buf_12 output674 (.A(net674),
    .X(sports_o[4]));
 sky130_fd_sc_hd__buf_12 output675 (.A(net675),
    .X(sports_o[50]));
 sky130_fd_sc_hd__buf_12 output676 (.A(net676),
    .X(sports_o[51]));
 sky130_fd_sc_hd__buf_12 output677 (.A(net677),
    .X(sports_o[52]));
 sky130_fd_sc_hd__buf_12 output678 (.A(net678),
    .X(sports_o[53]));
 sky130_fd_sc_hd__buf_12 output679 (.A(net679),
    .X(sports_o[54]));
 sky130_fd_sc_hd__buf_12 output680 (.A(net680),
    .X(sports_o[55]));
 sky130_fd_sc_hd__buf_12 output681 (.A(net681),
    .X(sports_o[56]));
 sky130_fd_sc_hd__buf_12 output682 (.A(net682),
    .X(sports_o[57]));
 sky130_fd_sc_hd__buf_12 output683 (.A(net683),
    .X(sports_o[58]));
 sky130_fd_sc_hd__buf_12 output684 (.A(net684),
    .X(sports_o[59]));
 sky130_fd_sc_hd__buf_12 output685 (.A(net685),
    .X(sports_o[5]));
 sky130_fd_sc_hd__buf_12 output686 (.A(net686),
    .X(sports_o[60]));
 sky130_fd_sc_hd__buf_12 output687 (.A(net687),
    .X(sports_o[61]));
 sky130_fd_sc_hd__buf_12 output688 (.A(net688),
    .X(sports_o[62]));
 sky130_fd_sc_hd__buf_12 output689 (.A(net689),
    .X(sports_o[63]));
 sky130_fd_sc_hd__buf_12 output690 (.A(net690),
    .X(sports_o[64]));
 sky130_fd_sc_hd__buf_12 output691 (.A(net691),
    .X(sports_o[65]));
 sky130_fd_sc_hd__buf_12 output692 (.A(net692),
    .X(sports_o[66]));
 sky130_fd_sc_hd__buf_12 output693 (.A(net693),
    .X(sports_o[67]));
 sky130_fd_sc_hd__buf_12 output694 (.A(net694),
    .X(sports_o[68]));
 sky130_fd_sc_hd__buf_12 output695 (.A(net695),
    .X(sports_o[69]));
 sky130_fd_sc_hd__buf_12 output696 (.A(net696),
    .X(sports_o[6]));
 sky130_fd_sc_hd__buf_12 output697 (.A(net697),
    .X(sports_o[70]));
 sky130_fd_sc_hd__buf_12 output698 (.A(net698),
    .X(sports_o[71]));
 sky130_fd_sc_hd__buf_12 output699 (.A(net699),
    .X(sports_o[72]));
 sky130_fd_sc_hd__buf_12 output700 (.A(net700),
    .X(sports_o[73]));
 sky130_fd_sc_hd__buf_12 output701 (.A(net701),
    .X(sports_o[74]));
 sky130_fd_sc_hd__buf_12 output702 (.A(net702),
    .X(sports_o[75]));
 sky130_fd_sc_hd__buf_12 output703 (.A(net703),
    .X(sports_o[76]));
 sky130_fd_sc_hd__buf_12 output704 (.A(net704),
    .X(sports_o[77]));
 sky130_fd_sc_hd__buf_12 output705 (.A(net705),
    .X(sports_o[78]));
 sky130_fd_sc_hd__buf_12 output706 (.A(net706),
    .X(sports_o[79]));
 sky130_fd_sc_hd__buf_12 output707 (.A(net707),
    .X(sports_o[7]));
 sky130_fd_sc_hd__buf_12 output708 (.A(net708),
    .X(sports_o[80]));
 sky130_fd_sc_hd__buf_12 output709 (.A(net709),
    .X(sports_o[81]));
 sky130_fd_sc_hd__buf_12 output710 (.A(net710),
    .X(sports_o[82]));
 sky130_fd_sc_hd__buf_12 output711 (.A(net711),
    .X(sports_o[83]));
 sky130_fd_sc_hd__buf_12 output712 (.A(net712),
    .X(sports_o[84]));
 sky130_fd_sc_hd__buf_12 output713 (.A(net713),
    .X(sports_o[85]));
 sky130_fd_sc_hd__buf_12 output714 (.A(net714),
    .X(sports_o[86]));
 sky130_fd_sc_hd__buf_12 output715 (.A(net715),
    .X(sports_o[87]));
 sky130_fd_sc_hd__buf_12 output716 (.A(net716),
    .X(sports_o[88]));
 sky130_fd_sc_hd__buf_12 output717 (.A(net717),
    .X(sports_o[89]));
 sky130_fd_sc_hd__buf_12 output718 (.A(net718),
    .X(sports_o[8]));
 sky130_fd_sc_hd__buf_12 output719 (.A(net719),
    .X(sports_o[90]));
 sky130_fd_sc_hd__buf_12 output720 (.A(net720),
    .X(sports_o[91]));
 sky130_fd_sc_hd__buf_12 output721 (.A(net721),
    .X(sports_o[92]));
 sky130_fd_sc_hd__buf_12 output722 (.A(net722),
    .X(sports_o[93]));
 sky130_fd_sc_hd__buf_12 output723 (.A(net723),
    .X(sports_o[94]));
 sky130_fd_sc_hd__buf_12 output724 (.A(net724),
    .X(sports_o[95]));
 sky130_fd_sc_hd__buf_12 output725 (.A(net725),
    .X(sports_o[96]));
 sky130_fd_sc_hd__buf_12 output726 (.A(net726),
    .X(sports_o[97]));
 sky130_fd_sc_hd__buf_12 output727 (.A(net727),
    .X(sports_o[98]));
 sky130_fd_sc_hd__buf_12 output728 (.A(net728),
    .X(sports_o[99]));
 sky130_fd_sc_hd__buf_12 output729 (.A(net729),
    .X(sports_o[9]));
 sky130_fd_sc_hd__clkbuf_4 wire730 (.A(_0666_),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_4 wire731 (.A(_3384_),
    .X(net731));
endmodule

