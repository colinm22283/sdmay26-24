// This is the unpowered netlist.
module wishbone_register_m (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    access_read_mask_i,
    access_write_mask_i,
    reg_o,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [31:0] access_read_mask_i;
 input [31:0] access_write_mask_i;
 output [31:0] reg_o;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire net165;
 wire net166;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA__095__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__096__D (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA__098__A0 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__100__A0 (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__102__A0 (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__104__A0 (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__106__A0 (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__108__A0 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__110__A0 (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__112__A0 (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__114__A0 (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__114__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__116__A0 (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__116__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__118__A0 (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__118__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__120__A0 (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__A0 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__128__A0 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__A0 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__132__A0 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__136__A0 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__138__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__A0 (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__140__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__142__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__A0 (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__144__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__146__A0 (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__146__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__148__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__150__A0 (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__150__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__152__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__154__A0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__154__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__156__A0 (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__156__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__158__S (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__161__A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA__162__A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__164__A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA__166__A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA__167__A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA__169__A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA__171__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__173__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__174__A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__175__A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__176__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__179__A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA__180__A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA__181__A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__182__A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA__183__A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA__184__A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA__185__A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__186__A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA__187__A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA__188__A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA__189__A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA__190__A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__191__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__192__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__193__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__194__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__195__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__196__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__197__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__198__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__199__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__200__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__217__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__218__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__219__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__220__A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold94_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_A (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_A (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net160));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_68 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_101 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_99 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__inv_2 _095_ (.A(net164),
    .Y(_001_));
 sky130_fd_sc_hd__and4_1 _096_ (.A(net96),
    .B(net97),
    .C(net64),
    .D(net129),
    .X(_063_));
 sky130_fd_sc_hd__and2_1 _097_ (.A(net55),
    .B(net210),
    .X(_064_));
 sky130_fd_sc_hd__mux2_1 _098_ (.A0(net121),
    .A1(_064_),
    .S(net161),
    .X(_062_));
 sky130_fd_sc_hd__and2_1 _099_ (.A(net53),
    .B(net237),
    .X(_065_));
 sky130_fd_sc_hd__mux2_1 _100_ (.A0(net119),
    .A1(_065_),
    .S(net161),
    .X(_061_));
 sky130_fd_sc_hd__and2_1 _101_ (.A(net52),
    .B(net219),
    .X(_066_));
 sky130_fd_sc_hd__mux2_1 _102_ (.A0(net118),
    .A1(_066_),
    .S(net161),
    .X(_060_));
 sky130_fd_sc_hd__and2_1 _103_ (.A(net51),
    .B(net252),
    .X(_067_));
 sky130_fd_sc_hd__mux2_1 _104_ (.A0(net117),
    .A1(_067_),
    .S(net161),
    .X(_059_));
 sky130_fd_sc_hd__and2_1 _105_ (.A(net50),
    .B(net207),
    .X(_068_));
 sky130_fd_sc_hd__mux2_1 _106_ (.A0(net116),
    .A1(_068_),
    .S(net161),
    .X(_058_));
 sky130_fd_sc_hd__and2_1 _107_ (.A(net49),
    .B(net243),
    .X(_069_));
 sky130_fd_sc_hd__mux2_1 _108_ (.A0(net115),
    .A1(_069_),
    .S(net161),
    .X(_057_));
 sky130_fd_sc_hd__and2_1 _109_ (.A(net48),
    .B(net246),
    .X(_070_));
 sky130_fd_sc_hd__mux2_1 _110_ (.A0(net114),
    .A1(_070_),
    .S(net161),
    .X(_056_));
 sky130_fd_sc_hd__and2_1 _111_ (.A(net47),
    .B(net258),
    .X(_071_));
 sky130_fd_sc_hd__mux2_1 _112_ (.A0(net113),
    .A1(_071_),
    .S(net161),
    .X(_055_));
 sky130_fd_sc_hd__and2_1 _113_ (.A(net46),
    .B(net249),
    .X(_072_));
 sky130_fd_sc_hd__mux2_1 _114_ (.A0(net112),
    .A1(_072_),
    .S(net162),
    .X(_054_));
 sky130_fd_sc_hd__and2_1 _115_ (.A(net45),
    .B(net240),
    .X(_073_));
 sky130_fd_sc_hd__mux2_1 _116_ (.A0(net111),
    .A1(_073_),
    .S(net162),
    .X(_053_));
 sky130_fd_sc_hd__and2_1 _117_ (.A(net44),
    .B(net213),
    .X(_074_));
 sky130_fd_sc_hd__mux2_1 _118_ (.A0(net110),
    .A1(_074_),
    .S(net162),
    .X(_052_));
 sky130_fd_sc_hd__and2_1 _119_ (.A(net42),
    .B(net255),
    .X(_075_));
 sky130_fd_sc_hd__mux2_1 _120_ (.A0(net108),
    .A1(_075_),
    .S(net161),
    .X(_051_));
 sky130_fd_sc_hd__and2_1 _121_ (.A(net41),
    .B(net216),
    .X(_076_));
 sky130_fd_sc_hd__mux2_1 _122_ (.A0(net107),
    .A1(_076_),
    .S(net162),
    .X(_050_));
 sky130_fd_sc_hd__and2_1 _123_ (.A(net40),
    .B(net222),
    .X(_077_));
 sky130_fd_sc_hd__mux2_1 _124_ (.A0(net106),
    .A1(_077_),
    .S(net161),
    .X(_049_));
 sky130_fd_sc_hd__and2_1 _125_ (.A(net39),
    .B(net234),
    .X(_078_));
 sky130_fd_sc_hd__mux2_1 _126_ (.A0(net105),
    .A1(_078_),
    .S(net161),
    .X(_048_));
 sky130_fd_sc_hd__and2_1 _127_ (.A(net38),
    .B(net195),
    .X(_079_));
 sky130_fd_sc_hd__mux2_1 _128_ (.A0(net104),
    .A1(_079_),
    .S(net161),
    .X(_047_));
 sky130_fd_sc_hd__and2_1 _129_ (.A(net37),
    .B(net231),
    .X(_080_));
 sky130_fd_sc_hd__mux2_1 _130_ (.A0(net103),
    .A1(_080_),
    .S(net161),
    .X(_046_));
 sky130_fd_sc_hd__and2_1 _131_ (.A(net36),
    .B(net228),
    .X(_081_));
 sky130_fd_sc_hd__mux2_1 _132_ (.A0(net102),
    .A1(_081_),
    .S(net161),
    .X(_045_));
 sky130_fd_sc_hd__and2_1 _133_ (.A(net35),
    .B(net225),
    .X(_082_));
 sky130_fd_sc_hd__mux2_1 _134_ (.A0(net101),
    .A1(_082_),
    .S(net161),
    .X(_044_));
 sky130_fd_sc_hd__and2_1 _135_ (.A(net34),
    .B(net189),
    .X(_083_));
 sky130_fd_sc_hd__mux2_1 _136_ (.A0(net100),
    .A1(_083_),
    .S(net161),
    .X(_043_));
 sky130_fd_sc_hd__and2_1 _137_ (.A(net33),
    .B(net201),
    .X(_084_));
 sky130_fd_sc_hd__mux2_1 _138_ (.A0(net99),
    .A1(_084_),
    .S(net162),
    .X(_042_));
 sky130_fd_sc_hd__and2_1 _139_ (.A(net62),
    .B(net183),
    .X(_085_));
 sky130_fd_sc_hd__mux2_1 _140_ (.A0(net128),
    .A1(_085_),
    .S(net162),
    .X(_041_));
 sky130_fd_sc_hd__and2_1 _141_ (.A(net61),
    .B(net204),
    .X(_086_));
 sky130_fd_sc_hd__mux2_1 _142_ (.A0(net127),
    .A1(_086_),
    .S(net162),
    .X(_040_));
 sky130_fd_sc_hd__and2_1 _143_ (.A(net60),
    .B(net186),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _144_ (.A0(net126),
    .A1(_087_),
    .S(net162),
    .X(_039_));
 sky130_fd_sc_hd__and2_1 _145_ (.A(net59),
    .B(net180),
    .X(_088_));
 sky130_fd_sc_hd__mux2_1 _146_ (.A0(net125),
    .A1(_088_),
    .S(net162),
    .X(_038_));
 sky130_fd_sc_hd__and2_1 _147_ (.A(net58),
    .B(net198),
    .X(_089_));
 sky130_fd_sc_hd__mux2_1 _148_ (.A0(net124),
    .A1(_089_),
    .S(net162),
    .X(_037_));
 sky130_fd_sc_hd__and2_1 _149_ (.A(net57),
    .B(net174),
    .X(_090_));
 sky130_fd_sc_hd__mux2_1 _150_ (.A0(net123),
    .A1(_090_),
    .S(net162),
    .X(_036_));
 sky130_fd_sc_hd__and2_1 _151_ (.A(net56),
    .B(net192),
    .X(_091_));
 sky130_fd_sc_hd__mux2_1 _152_ (.A0(net122),
    .A1(_091_),
    .S(net162),
    .X(_035_));
 sky130_fd_sc_hd__and2_1 _153_ (.A(net54),
    .B(net177),
    .X(_092_));
 sky130_fd_sc_hd__mux2_1 _154_ (.A0(net120),
    .A1(_092_),
    .S(net162),
    .X(_034_));
 sky130_fd_sc_hd__and2_1 _155_ (.A(net43),
    .B(net171),
    .X(_093_));
 sky130_fd_sc_hd__mux2_1 _156_ (.A0(net109),
    .A1(_093_),
    .S(net162),
    .X(_033_));
 sky130_fd_sc_hd__and2_1 _157_ (.A(net32),
    .B(net168),
    .X(_094_));
 sky130_fd_sc_hd__mux2_1 _158_ (.A0(net98),
    .A1(_094_),
    .S(net162),
    .X(_032_));
 sky130_fd_sc_hd__and3b_1 _159_ (.A_N(net260),
    .B(net64),
    .C(net96),
    .X(_000_));
 sky130_fd_sc_hd__and2_1 _160_ (.A(net98),
    .B(net1),
    .X(net130));
 sky130_fd_sc_hd__and2_1 _161_ (.A(net109),
    .B(net12),
    .X(net141));
 sky130_fd_sc_hd__and2_1 _162_ (.A(net120),
    .B(net23),
    .X(net152));
 sky130_fd_sc_hd__and2_1 _163_ (.A(net122),
    .B(net25),
    .X(net154));
 sky130_fd_sc_hd__and2_2 _164_ (.A(net123),
    .B(net26),
    .X(net155));
 sky130_fd_sc_hd__and2_1 _165_ (.A(net124),
    .B(net27),
    .X(net156));
 sky130_fd_sc_hd__and2_2 _166_ (.A(net125),
    .B(net28),
    .X(net157));
 sky130_fd_sc_hd__and2_1 _167_ (.A(net126),
    .B(net29),
    .X(net158));
 sky130_fd_sc_hd__and2_1 _168_ (.A(net127),
    .B(net30),
    .X(net159));
 sky130_fd_sc_hd__and2_2 _169_ (.A(net128),
    .B(net31),
    .X(net160));
 sky130_fd_sc_hd__and2_1 _170_ (.A(net99),
    .B(net2),
    .X(net131));
 sky130_fd_sc_hd__and2_2 _171_ (.A(net100),
    .B(net3),
    .X(net132));
 sky130_fd_sc_hd__and2_1 _172_ (.A(net101),
    .B(net4),
    .X(net133));
 sky130_fd_sc_hd__and2_2 _173_ (.A(net102),
    .B(net5),
    .X(net134));
 sky130_fd_sc_hd__and2_2 _174_ (.A(net103),
    .B(net6),
    .X(net135));
 sky130_fd_sc_hd__and2_1 _175_ (.A(net104),
    .B(net7),
    .X(net136));
 sky130_fd_sc_hd__and2_2 _176_ (.A(net105),
    .B(net8),
    .X(net137));
 sky130_fd_sc_hd__and2_1 _177_ (.A(net106),
    .B(net9),
    .X(net138));
 sky130_fd_sc_hd__and2_1 _178_ (.A(net107),
    .B(net10),
    .X(net139));
 sky130_fd_sc_hd__and2_2 _179_ (.A(net108),
    .B(net11),
    .X(net140));
 sky130_fd_sc_hd__and2_1 _180_ (.A(net110),
    .B(net13),
    .X(net142));
 sky130_fd_sc_hd__and2_2 _181_ (.A(net111),
    .B(net14),
    .X(net143));
 sky130_fd_sc_hd__and2_1 _182_ (.A(net112),
    .B(net15),
    .X(net144));
 sky130_fd_sc_hd__and2_1 _183_ (.A(net113),
    .B(net16),
    .X(net145));
 sky130_fd_sc_hd__and2_1 _184_ (.A(net114),
    .B(net17),
    .X(net146));
 sky130_fd_sc_hd__and2_1 _185_ (.A(net115),
    .B(net18),
    .X(net147));
 sky130_fd_sc_hd__and2_1 _186_ (.A(net116),
    .B(net19),
    .X(net148));
 sky130_fd_sc_hd__and2_1 _187_ (.A(net117),
    .B(net20),
    .X(net149));
 sky130_fd_sc_hd__and2_1 _188_ (.A(net118),
    .B(net21),
    .X(net150));
 sky130_fd_sc_hd__and2_1 _189_ (.A(net119),
    .B(net22),
    .X(net151));
 sky130_fd_sc_hd__and2_1 _190_ (.A(net121),
    .B(net24),
    .X(net153));
 sky130_fd_sc_hd__inv_2 _191_ (.A(net164),
    .Y(_002_));
 sky130_fd_sc_hd__inv_2 _192_ (.A(net164),
    .Y(_003_));
 sky130_fd_sc_hd__inv_2 _193_ (.A(net164),
    .Y(_004_));
 sky130_fd_sc_hd__inv_2 _194_ (.A(net164),
    .Y(_005_));
 sky130_fd_sc_hd__inv_2 _195_ (.A(net164),
    .Y(_006_));
 sky130_fd_sc_hd__inv_2 _196_ (.A(net164),
    .Y(_007_));
 sky130_fd_sc_hd__inv_2 _197_ (.A(net164),
    .Y(_008_));
 sky130_fd_sc_hd__inv_2 _198_ (.A(net164),
    .Y(_009_));
 sky130_fd_sc_hd__inv_2 _199_ (.A(net164),
    .Y(_010_));
 sky130_fd_sc_hd__inv_2 _200_ (.A(net164),
    .Y(_011_));
 sky130_fd_sc_hd__inv_2 _201_ (.A(net163),
    .Y(_012_));
 sky130_fd_sc_hd__inv_2 _202_ (.A(net163),
    .Y(_013_));
 sky130_fd_sc_hd__inv_2 _203_ (.A(net163),
    .Y(_014_));
 sky130_fd_sc_hd__inv_2 _204_ (.A(net163),
    .Y(_015_));
 sky130_fd_sc_hd__inv_2 _205_ (.A(net163),
    .Y(_016_));
 sky130_fd_sc_hd__inv_2 _206_ (.A(net163),
    .Y(_017_));
 sky130_fd_sc_hd__inv_2 _207_ (.A(net163),
    .Y(_018_));
 sky130_fd_sc_hd__inv_2 _208_ (.A(net163),
    .Y(_019_));
 sky130_fd_sc_hd__inv_2 _209_ (.A(net163),
    .Y(_020_));
 sky130_fd_sc_hd__inv_2 _210_ (.A(net163),
    .Y(_021_));
 sky130_fd_sc_hd__inv_2 _211_ (.A(net163),
    .Y(_022_));
 sky130_fd_sc_hd__inv_2 _212_ (.A(net163),
    .Y(_023_));
 sky130_fd_sc_hd__inv_2 _213_ (.A(net163),
    .Y(_024_));
 sky130_fd_sc_hd__inv_2 _214_ (.A(net163),
    .Y(_025_));
 sky130_fd_sc_hd__inv_2 _215_ (.A(net163),
    .Y(_026_));
 sky130_fd_sc_hd__inv_2 _216_ (.A(net163),
    .Y(_027_));
 sky130_fd_sc_hd__inv_2 _217_ (.A(net164),
    .Y(_028_));
 sky130_fd_sc_hd__inv_2 _218_ (.A(net164),
    .Y(_029_));
 sky130_fd_sc_hd__inv_2 _219_ (.A(net164),
    .Y(_030_));
 sky130_fd_sc_hd__inv_2 _220_ (.A(net164),
    .Y(_031_));
 sky130_fd_sc_hd__dfrtp_2 _221_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(net169),
    .RESET_B(_001_),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_4 _222_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(net172),
    .RESET_B(_002_),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_4 _223_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(net178),
    .RESET_B(_003_),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_4 _224_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(net193),
    .RESET_B(_004_),
    .Q(net122));
 sky130_fd_sc_hd__dfrtp_4 _225_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(net175),
    .RESET_B(_005_),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_4 _226_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(net199),
    .RESET_B(_006_),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_4 _227_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(net181),
    .RESET_B(_007_),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_4 _228_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(net187),
    .RESET_B(_008_),
    .Q(net126));
 sky130_fd_sc_hd__dfrtp_2 _229_ (.CLK(clknet_2_1__leaf_wb_clk_i),
    .D(net205),
    .RESET_B(_009_),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_4 _230_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(net184),
    .RESET_B(_010_),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_2 _231_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net202),
    .RESET_B(_011_),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_4 _232_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(net190),
    .RESET_B(_012_),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_4 _233_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net226),
    .RESET_B(_013_),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_4 _234_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(net229),
    .RESET_B(_014_),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_4 _235_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(net232),
    .RESET_B(_015_),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_4 _236_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(net196),
    .RESET_B(_016_),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_4 _237_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(net235),
    .RESET_B(_017_),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_4 _238_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net223),
    .RESET_B(_018_),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_4 _239_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net217),
    .RESET_B(_019_),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_4 _240_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(net256),
    .RESET_B(_020_),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_4 _241_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(net214),
    .RESET_B(_021_),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_4 _242_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(net241),
    .RESET_B(_022_),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_4 _243_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(net250),
    .RESET_B(_023_),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_4 _244_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net259),
    .RESET_B(_024_),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_4 _245_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net247),
    .RESET_B(_025_),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_4 _246_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net244),
    .RESET_B(_026_),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_4 _247_ (.CLK(clknet_2_2__leaf_wb_clk_i),
    .D(net208),
    .RESET_B(_027_),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_4 _248_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net253),
    .RESET_B(_028_),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_4 _249_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net220),
    .RESET_B(_029_),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_4 _250_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net238),
    .RESET_B(_030_),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_4 _251_ (.CLK(clknet_2_3__leaf_wb_clk_i),
    .D(net211),
    .RESET_B(_031_),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_2 _252_ (.CLK(clknet_2_0__leaf_wb_clk_i),
    .D(net261),
    .Q(net129));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_2__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_2_3__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_8 fanout161 (.A(net162),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_8 fanout162 (.A(_063_),
    .X(net162));
 sky130_fd_sc_hd__buf_8 fanout163 (.A(net164),
    .X(net163));
 sky130_fd_sc_hd__buf_8 fanout164 (.A(net63),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(wbs_dat_i[0]),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(wbs_dat_i[2]),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net87),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(_034_),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(wbs_dat_i[6]),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net92),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(_038_),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(wbs_dat_i[9]),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net95),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(_041_),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(wbs_dat_i[7]),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net65),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net93),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(_039_),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(wbs_dat_i[11]),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net67),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(_043_),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(wbs_dat_i[3]),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net89),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(_035_),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(wbs_dat_i[15]),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net71),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_032_),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(_047_),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(wbs_dat_i[5]),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(net91),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_037_),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(wbs_dat_i[10]),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net66),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(_042_),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(wbs_dat_i[8]),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net94),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(_040_),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(wbs_dat_i[1]),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(wbs_dat_i[26]),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net83),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(_058_),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(wbs_dat_i[30]),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net88),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(_062_),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(wbs_dat_i[20]),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net77),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(_052_),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(wbs_dat_i[18]),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net76),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net74),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(_050_),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(wbs_dat_i[28]),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net85),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(_060_),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(wbs_dat_i[17]),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net73),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(_049_),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(wbs_dat_i[12]),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net68),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(_033_),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(_044_),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(wbs_dat_i[13]),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net69),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(_045_),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(wbs_dat_i[14]),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net70),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(_046_),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(wbs_dat_i[16]),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net72),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(_048_),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(wbs_dat_i[4]),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(wbs_dat_i[29]),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net86),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(_061_),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(wbs_dat_i[21]),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net78),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(_053_),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(wbs_dat_i[25]),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net82),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_057_),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(wbs_dat_i[24]),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net90),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net81),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(_056_),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(wbs_dat_i[22]),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net79),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(_054_),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(wbs_dat_i[27]),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(net84),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(_059_),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(wbs_dat_i[19]),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(net75),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(_036_),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(_051_),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(wbs_dat_i[23]),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net80),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(_055_),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net129),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(_000_),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(access_read_mask_i[0]),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input10 (.A(access_read_mask_i[18]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(access_read_mask_i[19]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(access_read_mask_i[1]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(access_read_mask_i[20]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(access_read_mask_i[21]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(access_read_mask_i[22]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(access_read_mask_i[23]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(access_read_mask_i[24]),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(access_read_mask_i[25]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(access_read_mask_i[26]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(access_read_mask_i[10]),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(access_read_mask_i[27]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(access_read_mask_i[28]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(access_read_mask_i[29]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(access_read_mask_i[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(access_read_mask_i[30]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(access_read_mask_i[3]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(access_read_mask_i[4]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(access_read_mask_i[5]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_1 input28 (.A(access_read_mask_i[6]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(access_read_mask_i[7]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(access_read_mask_i[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(access_read_mask_i[8]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(access_read_mask_i[9]),
    .X(net31));
 sky130_fd_sc_hd__buf_1 input32 (.A(access_write_mask_i[0]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(access_write_mask_i[10]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_1 input34 (.A(access_write_mask_i[11]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(access_write_mask_i[12]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(access_write_mask_i[13]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(access_write_mask_i[14]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(access_write_mask_i[15]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 input39 (.A(access_write_mask_i[16]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input4 (.A(access_read_mask_i[12]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input40 (.A(access_write_mask_i[17]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(access_write_mask_i[18]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(access_write_mask_i[19]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(access_write_mask_i[1]),
    .X(net43));
 sky130_fd_sc_hd__buf_1 input44 (.A(access_write_mask_i[20]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(access_write_mask_i[21]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(access_write_mask_i[22]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(access_write_mask_i[23]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(access_write_mask_i[24]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(access_write_mask_i[25]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input5 (.A(access_read_mask_i[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input50 (.A(access_write_mask_i[26]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(access_write_mask_i[27]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(access_write_mask_i[28]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(access_write_mask_i[29]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(access_write_mask_i[2]),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(access_write_mask_i[30]),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(access_write_mask_i[3]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(access_write_mask_i[4]),
    .X(net57));
 sky130_fd_sc_hd__buf_1 input58 (.A(access_write_mask_i[5]),
    .X(net58));
 sky130_fd_sc_hd__buf_1 input59 (.A(access_write_mask_i[6]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(access_read_mask_i[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_1 input60 (.A(access_write_mask_i[7]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(access_write_mask_i[8]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 input62 (.A(access_write_mask_i[9]),
    .X(net62));
 sky130_fd_sc_hd__buf_1 input63 (.A(wb_rst_i),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(wbs_cyc_i),
    .X(net64));
 sky130_fd_sc_hd__buf_1 input65 (.A(net167),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(net200),
    .X(net66));
 sky130_fd_sc_hd__buf_1 input67 (.A(net188),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(net224),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(net227),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input7 (.A(access_read_mask_i[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(net230),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(net194),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(net233),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(net221),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 input74 (.A(net215),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 input75 (.A(net254),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(net170),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 input77 (.A(net212),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 input78 (.A(net239),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(net248),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(access_read_mask_i[16]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input80 (.A(net257),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(net245),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(net242),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(net206),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(net251),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(net218),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(net236),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(net176),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 input88 (.A(net209),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(net191),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input9 (.A(access_read_mask_i[17]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(net173),
    .X(net90));
 sky130_fd_sc_hd__buf_1 input91 (.A(net197),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(net179),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 input93 (.A(net185),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(net203),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 input95 (.A(net182),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(wbs_stb_i),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(wbs_we_i),
    .X(net97));
 sky130_fd_sc_hd__buf_12 output100 (.A(net100),
    .X(reg_o[11]));
 sky130_fd_sc_hd__buf_12 output101 (.A(net101),
    .X(reg_o[12]));
 sky130_fd_sc_hd__buf_12 output102 (.A(net102),
    .X(reg_o[13]));
 sky130_fd_sc_hd__buf_12 output103 (.A(net103),
    .X(reg_o[14]));
 sky130_fd_sc_hd__buf_12 output104 (.A(net104),
    .X(reg_o[15]));
 sky130_fd_sc_hd__buf_12 output105 (.A(net105),
    .X(reg_o[16]));
 sky130_fd_sc_hd__buf_12 output106 (.A(net106),
    .X(reg_o[17]));
 sky130_fd_sc_hd__buf_12 output107 (.A(net107),
    .X(reg_o[18]));
 sky130_fd_sc_hd__buf_12 output108 (.A(net108),
    .X(reg_o[19]));
 sky130_fd_sc_hd__buf_12 output109 (.A(net109),
    .X(reg_o[1]));
 sky130_fd_sc_hd__buf_12 output110 (.A(net110),
    .X(reg_o[20]));
 sky130_fd_sc_hd__buf_12 output111 (.A(net111),
    .X(reg_o[21]));
 sky130_fd_sc_hd__buf_12 output112 (.A(net112),
    .X(reg_o[22]));
 sky130_fd_sc_hd__buf_12 output113 (.A(net113),
    .X(reg_o[23]));
 sky130_fd_sc_hd__buf_12 output114 (.A(net114),
    .X(reg_o[24]));
 sky130_fd_sc_hd__buf_12 output115 (.A(net115),
    .X(reg_o[25]));
 sky130_fd_sc_hd__buf_12 output116 (.A(net116),
    .X(reg_o[26]));
 sky130_fd_sc_hd__buf_12 output117 (.A(net117),
    .X(reg_o[27]));
 sky130_fd_sc_hd__buf_12 output118 (.A(net118),
    .X(reg_o[28]));
 sky130_fd_sc_hd__buf_12 output119 (.A(net119),
    .X(reg_o[29]));
 sky130_fd_sc_hd__buf_12 output120 (.A(net120),
    .X(reg_o[2]));
 sky130_fd_sc_hd__buf_12 output121 (.A(net121),
    .X(reg_o[30]));
 sky130_fd_sc_hd__buf_12 output122 (.A(net122),
    .X(reg_o[3]));
 sky130_fd_sc_hd__buf_12 output123 (.A(net123),
    .X(reg_o[4]));
 sky130_fd_sc_hd__buf_12 output124 (.A(net124),
    .X(reg_o[5]));
 sky130_fd_sc_hd__buf_12 output125 (.A(net125),
    .X(reg_o[6]));
 sky130_fd_sc_hd__buf_12 output126 (.A(net126),
    .X(reg_o[7]));
 sky130_fd_sc_hd__buf_12 output127 (.A(net127),
    .X(reg_o[8]));
 sky130_fd_sc_hd__buf_12 output128 (.A(net128),
    .X(reg_o[9]));
 sky130_fd_sc_hd__buf_12 output129 (.A(net129),
    .X(wbs_ack_o));
 sky130_fd_sc_hd__buf_12 output130 (.A(net130),
    .X(wbs_dat_o[0]));
 sky130_fd_sc_hd__buf_12 output131 (.A(net131),
    .X(wbs_dat_o[10]));
 sky130_fd_sc_hd__buf_12 output132 (.A(net132),
    .X(wbs_dat_o[11]));
 sky130_fd_sc_hd__buf_12 output133 (.A(net133),
    .X(wbs_dat_o[12]));
 sky130_fd_sc_hd__buf_12 output134 (.A(net134),
    .X(wbs_dat_o[13]));
 sky130_fd_sc_hd__buf_12 output135 (.A(net135),
    .X(wbs_dat_o[14]));
 sky130_fd_sc_hd__buf_12 output136 (.A(net136),
    .X(wbs_dat_o[15]));
 sky130_fd_sc_hd__buf_12 output137 (.A(net137),
    .X(wbs_dat_o[16]));
 sky130_fd_sc_hd__buf_12 output138 (.A(net138),
    .X(wbs_dat_o[17]));
 sky130_fd_sc_hd__buf_12 output139 (.A(net139),
    .X(wbs_dat_o[18]));
 sky130_fd_sc_hd__buf_12 output140 (.A(net140),
    .X(wbs_dat_o[19]));
 sky130_fd_sc_hd__buf_12 output141 (.A(net141),
    .X(wbs_dat_o[1]));
 sky130_fd_sc_hd__buf_12 output142 (.A(net142),
    .X(wbs_dat_o[20]));
 sky130_fd_sc_hd__buf_12 output143 (.A(net143),
    .X(wbs_dat_o[21]));
 sky130_fd_sc_hd__buf_12 output144 (.A(net144),
    .X(wbs_dat_o[22]));
 sky130_fd_sc_hd__buf_12 output145 (.A(net145),
    .X(wbs_dat_o[23]));
 sky130_fd_sc_hd__buf_12 output146 (.A(net146),
    .X(wbs_dat_o[24]));
 sky130_fd_sc_hd__buf_12 output147 (.A(net147),
    .X(wbs_dat_o[25]));
 sky130_fd_sc_hd__buf_12 output148 (.A(net148),
    .X(wbs_dat_o[26]));
 sky130_fd_sc_hd__buf_12 output149 (.A(net149),
    .X(wbs_dat_o[27]));
 sky130_fd_sc_hd__buf_12 output150 (.A(net150),
    .X(wbs_dat_o[28]));
 sky130_fd_sc_hd__buf_12 output151 (.A(net151),
    .X(wbs_dat_o[29]));
 sky130_fd_sc_hd__buf_12 output152 (.A(net152),
    .X(wbs_dat_o[2]));
 sky130_fd_sc_hd__buf_12 output153 (.A(net153),
    .X(wbs_dat_o[30]));
 sky130_fd_sc_hd__buf_12 output154 (.A(net154),
    .X(wbs_dat_o[3]));
 sky130_fd_sc_hd__buf_12 output155 (.A(net155),
    .X(wbs_dat_o[4]));
 sky130_fd_sc_hd__buf_12 output156 (.A(net156),
    .X(wbs_dat_o[5]));
 sky130_fd_sc_hd__buf_12 output157 (.A(net157),
    .X(wbs_dat_o[6]));
 sky130_fd_sc_hd__buf_12 output158 (.A(net158),
    .X(wbs_dat_o[7]));
 sky130_fd_sc_hd__buf_12 output159 (.A(net159),
    .X(wbs_dat_o[8]));
 sky130_fd_sc_hd__buf_12 output160 (.A(net160),
    .X(wbs_dat_o[9]));
 sky130_fd_sc_hd__buf_12 output98 (.A(net98),
    .X(reg_o[0]));
 sky130_fd_sc_hd__buf_12 output99 (.A(net99),
    .X(reg_o[10]));
 sky130_fd_sc_hd__conb_1 wishbone_register_m_165 (.LO(net165));
 sky130_fd_sc_hd__conb_1 wishbone_register_m_166 (.LO(net166));
 assign reg_o[31] = net165;
 assign wbs_dat_o[31] = net166;
endmodule

